magic
tech sky130A
magscale 1 2
timestamp 1624074425
<< locali >>
rect 51199 56294 51233 56408
rect 39679 44750 39713 45012
rect 7903 21144 7937 21184
rect 8191 21144 8225 21184
rect 7903 21110 8225 21144
rect 7903 19812 7937 19852
rect 8191 19812 8225 19852
rect 7903 19778 8225 19812
rect 9343 18480 9377 18520
rect 8321 18446 8479 18480
rect 8993 18446 9377 18480
rect 8767 17188 9089 17222
rect 8767 17148 8801 17188
rect 8671 17114 8801 17148
rect 8671 16926 8705 17114
rect 9055 17074 9089 17188
rect 56863 11672 56897 11786
rect 37951 10858 37985 11046
rect 8191 9156 8225 9196
rect 8095 9122 8225 9156
rect 8095 8860 8129 9122
rect 9343 8268 9377 8456
rect 25087 8194 25121 8308
rect 37951 8194 37985 8382
rect 46015 8342 46049 8456
rect 47743 8416 47777 8530
rect 46015 8308 46241 8342
rect 46207 8120 46241 8308
rect 8479 7824 8513 7864
rect 8383 7790 8513 7824
rect 8383 7528 8417 7790
rect 19327 7602 19361 7716
rect 28927 7528 28961 7790
rect 34015 7528 34049 7716
rect 37087 7528 37121 7864
rect 45823 7602 45857 7716
rect 46687 7602 46721 7790
rect 10015 6862 10049 6976
rect 18175 6270 18209 6458
rect 27775 6344 27809 6458
rect 28447 6270 28481 6458
rect 29599 6122 29633 6236
rect 32767 6122 32801 6310
rect 36031 6270 36065 6384
rect 36223 6270 36257 6458
rect 7711 5160 7745 5200
rect 7903 5200 8225 5234
rect 7903 5160 7937 5200
rect 7711 5126 7937 5160
rect 8191 5160 8225 5200
rect 8191 5126 8383 5160
rect 10687 3606 10721 3794
rect 24223 3606 24257 3794
rect 12703 3088 12737 3202
rect 48511 2792 48545 3202
<< viali >>
rect 56767 57148 56801 57182
rect 9919 57000 9953 57034
rect 13951 57000 13985 57034
rect 32575 57000 32609 57034
rect 1951 56926 1985 56960
rect 2815 56926 2849 56960
rect 5311 56926 5345 56960
rect 5791 56926 5825 56960
rect 7423 56926 7457 56960
rect 8095 56926 8129 56960
rect 11455 56926 11489 56960
rect 13183 56926 13217 56960
rect 15103 56926 15137 56960
rect 16351 56926 16385 56960
rect 18175 56926 18209 56960
rect 19519 56926 19553 56960
rect 21055 56926 21089 56960
rect 22015 56926 22049 56960
rect 24223 56926 24257 56960
rect 25951 56926 25985 56960
rect 27391 56926 27425 56960
rect 28639 56926 28673 56960
rect 30271 56926 30305 56960
rect 31711 56926 31745 56960
rect 34303 56926 34337 56960
rect 34879 56926 34913 56960
rect 38047 56926 38081 56960
rect 41983 56926 42017 56960
rect 47551 56926 47585 56960
rect 52735 56926 52769 56960
rect 1759 56852 1793 56886
rect 2623 56852 2657 56886
rect 5119 56852 5153 56886
rect 7231 56852 7265 56886
rect 11263 56852 11297 56886
rect 12991 56852 13025 56886
rect 14047 56852 14081 56886
rect 16159 56852 16193 56886
rect 17983 56852 18017 56886
rect 19327 56852 19361 56886
rect 20863 56852 20897 56886
rect 24031 56852 24065 56886
rect 27199 56852 27233 56886
rect 30079 56852 30113 56886
rect 32671 56852 32705 56886
rect 34111 56852 34145 56886
rect 36991 56852 37025 56886
rect 40063 56852 40097 56886
rect 40735 56852 40769 56886
rect 43231 56852 43265 56886
rect 45055 56852 45089 56886
rect 46303 56852 46337 56886
rect 48991 56852 49025 56886
rect 51103 56852 51137 56886
rect 54271 56852 54305 56886
rect 55807 56852 55841 56886
rect 57055 56852 57089 56886
rect 40543 56778 40577 56812
rect 9823 56704 9857 56738
rect 36703 56704 36737 56738
rect 39775 56704 39809 56738
rect 40831 56704 40865 56738
rect 42943 56704 42977 56738
rect 44767 56704 44801 56738
rect 46015 56704 46049 56738
rect 48703 56704 48737 56738
rect 50815 56704 50849 56738
rect 53983 56704 54017 56738
rect 55519 56704 55553 56738
rect 1663 56482 1697 56516
rect 2431 56482 2465 56516
rect 3199 56482 3233 56516
rect 4447 56482 4481 56516
rect 5503 56482 5537 56516
rect 6271 56482 6305 56516
rect 7135 56482 7169 56516
rect 8479 56482 8513 56516
rect 10303 56482 10337 56516
rect 11071 56482 11105 56516
rect 11839 56482 11873 56516
rect 12607 56482 12641 56516
rect 13471 56482 13505 56516
rect 15103 56482 15137 56516
rect 17215 56482 17249 56516
rect 18175 56482 18209 56516
rect 18943 56482 18977 56516
rect 20287 56482 20321 56516
rect 21439 56482 21473 56516
rect 22111 56482 22145 56516
rect 22975 56482 23009 56516
rect 24415 56482 24449 56516
rect 26047 56482 26081 56516
rect 26911 56482 26945 56516
rect 27775 56482 27809 56516
rect 28447 56482 28481 56516
rect 29695 56482 29729 56516
rect 30847 56482 30881 56516
rect 31615 56482 31649 56516
rect 32383 56482 32417 56516
rect 33919 56482 33953 56516
rect 34783 56482 34817 56516
rect 36127 56482 36161 56516
rect 36991 56482 37025 56516
rect 37759 56482 37793 56516
rect 38719 56482 38753 56516
rect 40159 56482 40193 56516
rect 41887 56482 41921 56516
rect 42751 56482 42785 56516
rect 43423 56482 43457 56516
rect 44191 56482 44225 56516
rect 45055 56482 45089 56516
rect 46687 56482 46721 56516
rect 48127 56482 48161 56516
rect 49759 56482 49793 56516
rect 50527 56482 50561 56516
rect 51967 56482 52001 56516
rect 53023 56482 53057 56516
rect 53791 56482 53825 56516
rect 54463 56482 54497 56516
rect 55231 56482 55265 56516
rect 56095 56482 56129 56516
rect 50335 56408 50369 56442
rect 51199 56408 51233 56442
rect 22207 56334 22241 56368
rect 31423 56334 31457 56368
rect 31711 56334 31745 56368
rect 41983 56334 42017 56368
rect 43519 56334 43553 56368
rect 26143 56260 26177 56294
rect 34015 56260 34049 56294
rect 45151 56260 45185 56294
rect 50623 56260 50657 56294
rect 51199 56260 51233 56294
rect 52063 56260 52097 56294
rect 54559 56260 54593 56294
rect 55711 56260 55745 56294
rect 55999 56260 56033 56294
rect 57823 56260 57857 56294
rect 1759 56186 1793 56220
rect 1951 56186 1985 56220
rect 2527 56186 2561 56220
rect 2911 56186 2945 56220
rect 3295 56186 3329 56220
rect 4255 56186 4289 56220
rect 4543 56186 4577 56220
rect 5215 56186 5249 56220
rect 5599 56186 5633 56220
rect 6079 56186 6113 56220
rect 6367 56186 6401 56220
rect 6943 56186 6977 56220
rect 7231 56186 7265 56220
rect 8575 56186 8609 56220
rect 10111 56186 10145 56220
rect 10399 56186 10433 56220
rect 11167 56186 11201 56220
rect 11551 56186 11585 56220
rect 11935 56186 11969 56220
rect 12703 56186 12737 56220
rect 13567 56186 13601 56220
rect 14719 56186 14753 56220
rect 15007 56186 15041 56220
rect 15487 56186 15521 56220
rect 15775 56186 15809 56220
rect 15871 56186 15905 56220
rect 16831 56186 16865 56220
rect 17119 56186 17153 56220
rect 18271 56186 18305 56220
rect 19039 56186 19073 56220
rect 20383 56186 20417 56220
rect 21055 56186 21089 56220
rect 21343 56186 21377 56220
rect 22687 56186 22721 56220
rect 22879 56186 22913 56220
rect 24127 56186 24161 56220
rect 24319 56186 24353 56220
rect 26527 56186 26561 56220
rect 26815 56186 26849 56220
rect 27487 56186 27521 56220
rect 27679 56186 27713 56220
rect 28159 56186 28193 56220
rect 28543 56186 28577 56220
rect 29311 56186 29345 56220
rect 29599 56186 29633 56220
rect 30943 56186 30977 56220
rect 32479 56186 32513 56220
rect 32959 56186 32993 56220
rect 33151 56186 33185 56220
rect 33247 56186 33281 56220
rect 34399 56186 34433 56220
rect 34687 56186 34721 56220
rect 35935 56186 35969 56220
rect 36223 56186 36257 56220
rect 36607 56186 36641 56220
rect 36895 56186 36929 56220
rect 37471 56186 37505 56220
rect 37663 56186 37697 56220
rect 38815 56186 38849 56220
rect 39871 56186 39905 56220
rect 40255 56186 40289 56220
rect 42463 56186 42497 56220
rect 42655 56186 42689 56220
rect 44287 56186 44321 56220
rect 46783 56186 46817 56220
rect 48223 56186 48257 56220
rect 48703 56186 48737 56220
rect 48895 56186 48929 56220
rect 48991 56186 49025 56220
rect 49567 56186 49601 56220
rect 49855 56186 49889 56220
rect 52639 56186 52673 56220
rect 52927 56186 52961 56220
rect 53215 56186 53249 56220
rect 53503 56186 53537 56220
rect 53695 56186 53729 56220
rect 55327 56186 55361 56220
rect 1663 55668 1697 55702
rect 4447 55668 4481 55702
rect 7615 55668 7649 55702
rect 9343 55668 9377 55702
rect 13951 55668 13985 55702
rect 20287 55668 20321 55702
rect 23551 55668 23585 55702
rect 24991 55668 25025 55702
rect 39295 55668 39329 55702
rect 40927 55668 40961 55702
rect 45631 55668 45665 55702
rect 47071 55668 47105 55702
rect 51871 55668 51905 55702
rect 56671 55668 56705 55702
rect 57727 55668 57761 55702
rect 51967 55594 52001 55628
rect 1759 55520 1793 55554
rect 4255 55520 4289 55554
rect 4543 55520 4577 55554
rect 7423 55520 7457 55554
rect 7711 55520 7745 55554
rect 9247 55520 9281 55554
rect 14047 55520 14081 55554
rect 20095 55520 20129 55554
rect 20383 55520 20417 55554
rect 23263 55520 23297 55554
rect 23455 55520 23489 55554
rect 24799 55520 24833 55554
rect 25087 55520 25121 55554
rect 27967 55520 28001 55554
rect 28255 55520 28289 55554
rect 29023 55520 29057 55554
rect 39199 55520 39233 55554
rect 40639 55520 40673 55554
rect 40831 55520 40865 55554
rect 45535 55520 45569 55554
rect 47167 55520 47201 55554
rect 49183 55520 49217 55554
rect 56383 55520 56417 55554
rect 56575 55520 56609 55554
rect 57439 55520 57473 55554
rect 57631 55520 57665 55554
rect 8959 55372 8993 55406
rect 13663 55372 13697 55406
rect 28927 55372 28961 55406
rect 38911 55372 38945 55406
rect 45247 55372 45281 55406
rect 49087 55372 49121 55406
rect 57919 55150 57953 55184
rect 27583 54854 27617 54888
rect 57631 54854 57665 54888
rect 57823 54854 57857 54888
rect 27295 54780 27329 54814
rect 25279 54706 25313 54740
rect 25663 54706 25697 54740
rect 26623 54706 26657 54740
rect 26911 54706 26945 54740
rect 57919 54336 57953 54370
rect 56575 54188 56609 54222
rect 57631 54188 57665 54222
rect 57823 54188 57857 54222
rect 58111 54188 58145 54222
rect 56383 54040 56417 54074
rect 57919 53818 57953 53852
rect 55807 53522 55841 53556
rect 55999 53522 56033 53556
rect 57823 53522 57857 53556
rect 32191 53448 32225 53482
rect 32479 53448 32513 53482
rect 2239 53374 2273 53408
rect 2623 53374 2657 53408
rect 17599 53374 17633 53408
rect 17983 53374 18017 53408
rect 39391 53374 39425 53408
rect 39583 53374 39617 53408
rect 43039 53374 43073 53408
rect 43135 53374 43169 53408
rect 57631 53374 57665 53408
rect 17695 53004 17729 53038
rect 6943 52856 6977 52890
rect 7231 52856 7265 52890
rect 37759 52338 37793 52372
rect 3103 52042 3137 52076
rect 3391 52042 3425 52076
rect 18079 52042 18113 52076
rect 18367 52042 18401 52076
rect 39775 52042 39809 52076
rect 40063 52042 40097 52076
rect 29503 51672 29537 51706
rect 10303 51450 10337 51484
rect 15775 50710 15809 50744
rect 16063 50710 16097 50744
rect 53599 50710 53633 50744
rect 53791 50710 53825 50744
rect 39487 50192 39521 50226
rect 57631 50192 57665 50226
rect 51583 50118 51617 50152
rect 39391 50044 39425 50078
rect 57535 50044 57569 50078
rect 11839 49378 11873 49412
rect 11935 49378 11969 49412
rect 15583 49378 15617 49412
rect 15679 49378 15713 49412
rect 52447 49378 52481 49412
rect 18559 49008 18593 49042
rect 3295 48860 3329 48894
rect 3583 48860 3617 48894
rect 49087 48860 49121 48894
rect 49375 48860 49409 48894
rect 22783 48712 22817 48746
rect 41311 48490 41345 48524
rect 4351 48046 4385 48080
rect 4447 48046 4481 48080
rect 52639 48046 52673 48080
rect 52831 48046 52865 48080
rect 34591 47528 34625 47562
rect 34687 47528 34721 47562
rect 6751 47010 6785 47044
rect 23647 46714 23681 46748
rect 23935 46714 23969 46748
rect 9631 46196 9665 46230
rect 9919 46196 9953 46230
rect 12607 46048 12641 46082
rect 35071 45678 35105 45712
rect 51679 45382 51713 45416
rect 51871 45382 51905 45416
rect 38815 45160 38849 45194
rect 39679 45012 39713 45046
rect 8191 44864 8225 44898
rect 8479 44864 8513 44898
rect 21055 44864 21089 44898
rect 21343 44864 21377 44898
rect 7615 44790 7649 44824
rect 53503 44938 53537 44972
rect 41215 44864 41249 44898
rect 39679 44716 39713 44750
rect 41023 44716 41057 44750
rect 11071 44050 11105 44084
rect 11359 44050 11393 44084
rect 12415 43532 12449 43566
rect 12703 43532 12737 43566
rect 50047 43532 50081 43566
rect 49951 43384 49985 43418
rect 6559 42718 6593 42752
rect 46399 42718 46433 42752
rect 46783 42718 46817 42752
rect 53983 42718 54017 42752
rect 54175 42718 54209 42752
rect 7711 42200 7745 42234
rect 7999 42200 8033 42234
rect 4735 41756 4769 41790
rect 27295 41386 27329 41420
rect 27583 41386 27617 41420
rect 8287 40942 8321 40976
rect 8575 40942 8609 40976
rect 12223 40868 12257 40902
rect 19615 40868 19649 40902
rect 19903 40868 19937 40902
rect 40543 40868 40577 40902
rect 12127 40720 12161 40754
rect 40351 40720 40385 40754
rect 45055 40054 45089 40088
rect 45247 40054 45281 40088
rect 45823 39832 45857 39866
rect 7135 39536 7169 39570
rect 23647 39536 23681 39570
rect 43807 39536 43841 39570
rect 44095 39536 44129 39570
rect 49567 39536 49601 39570
rect 49375 39462 49409 39496
rect 6751 39388 6785 39422
rect 15295 38796 15329 38830
rect 47935 38722 47969 38756
rect 48031 38722 48065 38756
rect 56959 38722 56993 38756
rect 57151 38722 57185 38756
rect 30751 38500 30785 38534
rect 14431 38204 14465 38238
rect 18271 38204 18305 38238
rect 23935 38204 23969 38238
rect 38719 38204 38753 38238
rect 29887 38130 29921 38164
rect 14239 38056 14273 38090
rect 18079 38056 18113 38090
rect 38527 38056 38561 38090
rect 32959 37464 32993 37498
rect 10975 37390 11009 37424
rect 11263 37390 11297 37424
rect 33247 37390 33281 37424
rect 57343 37390 57377 37424
rect 43999 36872 44033 36906
rect 44191 36872 44225 36906
rect 15007 36058 15041 36092
rect 15199 36058 15233 36092
rect 40063 36058 40097 36092
rect 40351 36058 40385 36092
rect 46399 36058 46433 36092
rect 46591 36058 46625 36092
rect 36031 35688 36065 35722
rect 52063 35614 52097 35648
rect 33247 35540 33281 35574
rect 33535 35540 33569 35574
rect 14815 34726 14849 34760
rect 15103 34726 15137 34760
rect 32671 34726 32705 34760
rect 32767 34726 32801 34760
rect 41503 34726 41537 34760
rect 47263 34208 47297 34242
rect 57151 33468 57185 33502
rect 57343 33468 57377 33502
rect 19039 33172 19073 33206
rect 47743 33172 47777 33206
rect 28255 33098 28289 33132
rect 42367 32876 42401 32910
rect 19039 32506 19073 32540
rect 13951 32062 13985 32096
rect 30943 32062 30977 32096
rect 34111 32062 34145 32096
rect 39871 31840 39905 31874
rect 58015 31692 58049 31726
rect 16927 30804 16961 30838
rect 17599 30730 17633 30764
rect 31807 30360 31841 30394
rect 29983 30286 30017 30320
rect 52447 29546 52481 29580
rect 52255 29472 52289 29506
rect 17791 29398 17825 29432
rect 19231 29398 19265 29432
rect 40351 29398 40385 29432
rect 50047 29398 50081 29432
rect 53695 29398 53729 29432
rect 54559 29398 54593 29432
rect 55711 29398 55745 29432
rect 14239 29176 14273 29210
rect 55711 29176 55745 29210
rect 55903 29176 55937 29210
rect 14431 29028 14465 29062
rect 46879 28954 46913 28988
rect 15295 28880 15329 28914
rect 44767 28880 44801 28914
rect 38143 28140 38177 28174
rect 38335 28140 38369 28174
rect 20383 28066 20417 28100
rect 41791 28066 41825 28100
rect 14335 27548 14369 27582
rect 55231 27548 55265 27582
rect 55423 27548 55457 27582
rect 14815 26882 14849 26916
rect 15103 26882 15137 26916
rect 28639 26734 28673 26768
rect 47263 26734 47297 26768
rect 47455 26734 47489 26768
rect 24223 26216 24257 26250
rect 39007 26216 39041 26250
rect 57343 26216 57377 26250
rect 55327 25846 55361 25880
rect 7039 25698 7073 25732
rect 7327 25698 7361 25732
rect 55519 25698 55553 25732
rect 4543 25402 4577 25436
rect 21151 25402 21185 25436
rect 21439 25402 21473 25436
rect 14623 24884 14657 24918
rect 49855 24884 49889 24918
rect 52543 24884 52577 24918
rect 11647 24070 11681 24104
rect 22879 24070 22913 24104
rect 35071 23848 35105 23882
rect 35263 23700 35297 23734
rect 12415 23552 12449 23586
rect 21727 23552 21761 23586
rect 42943 23552 42977 23586
rect 13279 22738 13313 22772
rect 42847 22738 42881 22772
rect 9151 22220 9185 22254
rect 34975 22220 35009 22254
rect 36511 22220 36545 22254
rect 20575 21702 20609 21736
rect 20863 21702 20897 21736
rect 9823 21406 9857 21440
rect 7615 21184 7649 21218
rect 7903 21184 7937 21218
rect 8191 21184 8225 21218
rect 15775 20888 15809 20922
rect 28255 20888 28289 20922
rect 37951 20444 37985 20478
rect 27103 20074 27137 20108
rect 53023 20074 53057 20108
rect 7615 19852 7649 19886
rect 7903 19852 7937 19886
rect 8191 19852 8225 19886
rect 44095 19556 44129 19590
rect 8383 18742 8417 18776
rect 7615 18520 7649 18554
rect 9343 18520 9377 18554
rect 8287 18446 8321 18480
rect 8479 18446 8513 18480
rect 8959 18446 8993 18480
rect 24415 18446 24449 18480
rect 24703 18446 24737 18480
rect 20671 18298 20705 18332
rect 51679 18224 51713 18258
rect 1759 17410 1793 17444
rect 7519 17188 7553 17222
rect 9055 17040 9089 17074
rect 8671 16892 8705 16926
rect 30463 16892 30497 16926
rect 7519 15856 7553 15890
rect 55327 15856 55361 15890
rect 55519 15856 55553 15890
rect 19231 15560 19265 15594
rect 19519 15560 19553 15594
rect 15103 14820 15137 14854
rect 18271 14746 18305 14780
rect 44383 14450 44417 14484
rect 51199 14228 51233 14262
rect 7615 14080 7649 14114
rect 15967 13858 16001 13892
rect 16255 13710 16289 13744
rect 11455 13414 11489 13448
rect 45151 13414 45185 13448
rect 56863 13192 56897 13226
rect 7615 13118 7649 13152
rect 56959 13044 56993 13078
rect 57823 12970 57857 13004
rect 57343 12526 57377 12560
rect 57631 12378 57665 12412
rect 57919 12378 57953 12412
rect 37471 12230 37505 12264
rect 37759 12230 37793 12264
rect 57727 12230 57761 12264
rect 2143 12156 2177 12190
rect 48991 12156 49025 12190
rect 49183 12156 49217 12190
rect 6559 12082 6593 12116
rect 7615 11786 7649 11820
rect 56863 11786 56897 11820
rect 56959 11786 56993 11820
rect 56575 11712 56609 11746
rect 56191 11638 56225 11672
rect 56479 11638 56513 11672
rect 56863 11638 56897 11672
rect 57247 11638 57281 11672
rect 23935 11564 23969 11598
rect 55903 11564 55937 11598
rect 57343 11416 57377 11450
rect 37951 11046 37985 11080
rect 56959 11046 56993 11080
rect 57247 11046 57281 11080
rect 56095 10972 56129 11006
rect 55999 10898 56033 10932
rect 57343 10898 57377 10932
rect 18847 10824 18881 10858
rect 19039 10824 19073 10858
rect 29407 10824 29441 10858
rect 37951 10824 37985 10858
rect 48607 10824 48641 10858
rect 48799 10824 48833 10858
rect 8095 10750 8129 10784
rect 9919 10750 9953 10784
rect 32479 10750 32513 10784
rect 54655 10750 54689 10784
rect 7615 10528 7649 10562
rect 56383 10528 56417 10562
rect 55903 10380 55937 10414
rect 56671 10380 56705 10414
rect 54751 10306 54785 10340
rect 55039 10306 55073 10340
rect 57439 10306 57473 10340
rect 39583 10232 39617 10266
rect 57359 10232 57393 10266
rect 55135 10084 55169 10118
rect 55807 10084 55841 10118
rect 56575 10084 56609 10118
rect 55231 9862 55265 9896
rect 55999 9862 56033 9896
rect 55615 9788 55649 9822
rect 56191 9788 56225 9822
rect 55903 9714 55937 9748
rect 54847 9640 54881 9674
rect 55135 9640 55169 9674
rect 57631 9640 57665 9674
rect 54367 9566 54401 9600
rect 54463 9566 54497 9600
rect 24223 9492 24257 9526
rect 24511 9492 24545 9526
rect 50335 9418 50369 9452
rect 52639 9418 52673 9452
rect 7519 9196 7553 9230
rect 8191 9196 8225 9230
rect 39583 9122 39617 9156
rect 49951 9122 49985 9156
rect 4735 8900 4769 8934
rect 54655 9048 54689 9082
rect 55423 9048 55457 9082
rect 53407 8974 53441 9008
rect 56575 8974 56609 9008
rect 57247 8974 57281 9008
rect 50719 8900 50753 8934
rect 52159 8900 52193 8934
rect 55039 8900 55073 8934
rect 55327 8900 55361 8934
rect 8095 8826 8129 8860
rect 53311 8752 53345 8786
rect 54559 8752 54593 8786
rect 2047 8530 2081 8564
rect 12031 8530 12065 8564
rect 47743 8530 47777 8564
rect 47839 8530 47873 8564
rect 52543 8530 52577 8564
rect 9343 8456 9377 8490
rect 9439 8456 9473 8490
rect 46015 8456 46049 8490
rect 1759 8382 1793 8416
rect 3295 8382 3329 8416
rect 4543 8382 4577 8416
rect 2239 8308 2273 8342
rect 2527 8308 2561 8342
rect 5503 8308 5537 8342
rect 5791 8308 5825 8342
rect 10591 8382 10625 8416
rect 12815 8382 12849 8416
rect 13663 8382 13697 8416
rect 37951 8382 37985 8416
rect 12607 8308 12641 8342
rect 16175 8308 16209 8342
rect 25087 8308 25121 8342
rect 1663 8234 1697 8268
rect 2431 8234 2465 8268
rect 3199 8234 3233 8268
rect 4447 8234 4481 8268
rect 7807 8234 7841 8268
rect 7903 8234 7937 8268
rect 9343 8234 9377 8268
rect 9727 8234 9761 8268
rect 9823 8234 9857 8268
rect 10495 8234 10529 8268
rect 11263 8234 11297 8268
rect 11359 8234 11393 8268
rect 12127 8234 12161 8268
rect 12895 8234 12929 8268
rect 13567 8234 13601 8268
rect 16255 8234 16289 8268
rect 16927 8234 16961 8268
rect 17023 8234 17057 8268
rect 47743 8382 47777 8416
rect 48127 8382 48161 8416
rect 48703 8382 48737 8416
rect 48895 8382 48929 8416
rect 50527 8308 50561 8342
rect 50719 8308 50753 8342
rect 52927 8308 52961 8342
rect 53215 8308 53249 8342
rect 55231 8308 55265 8342
rect 55999 8308 56033 8342
rect 57151 8308 57185 8342
rect 25087 8160 25121 8194
rect 29791 8160 29825 8194
rect 37951 8160 37985 8194
rect 48223 8234 48257 8268
rect 48991 8234 49025 8268
rect 49663 8234 49697 8268
rect 49759 8234 49793 8268
rect 52447 8234 52481 8268
rect 53311 8234 53345 8268
rect 53983 8234 54017 8268
rect 54079 8234 54113 8268
rect 30943 8086 30977 8120
rect 34399 8086 34433 8120
rect 35071 8086 35105 8120
rect 46207 8086 46241 8120
rect 52159 8086 52193 8120
rect 3679 7864 3713 7898
rect 8479 7864 8513 7898
rect 12031 7864 12065 7898
rect 25951 7864 25985 7898
rect 29119 7864 29153 7898
rect 37087 7864 37121 7898
rect 44479 7864 44513 7898
rect 45247 7864 45281 7898
rect 5311 7790 5345 7824
rect 28927 7790 28961 7824
rect 3295 7716 3329 7750
rect 4063 7716 4097 7750
rect 4831 7716 4865 7750
rect 5599 7716 5633 7750
rect 1567 7642 1601 7676
rect 2239 7568 2273 7602
rect 2527 7568 2561 7602
rect 9151 7716 9185 7750
rect 9439 7716 9473 7750
rect 9919 7716 9953 7750
rect 10207 7716 10241 7750
rect 12319 7716 12353 7750
rect 13183 7716 13217 7750
rect 15583 7716 15617 7750
rect 15775 7716 15809 7750
rect 19327 7716 19361 7750
rect 20959 7716 20993 7750
rect 23935 7716 23969 7750
rect 24703 7716 24737 7750
rect 25471 7716 25505 7750
rect 26143 7716 26177 7750
rect 28255 7716 28289 7750
rect 10975 7642 11009 7676
rect 27967 7642 28001 7676
rect 13663 7568 13697 7602
rect 13951 7568 13985 7602
rect 19327 7568 19361 7602
rect 27007 7568 27041 7602
rect 29407 7716 29441 7750
rect 30175 7716 30209 7750
rect 30847 7716 30881 7750
rect 31135 7716 31169 7750
rect 31423 7716 31457 7750
rect 34015 7716 34049 7750
rect 34303 7716 34337 7750
rect 34591 7716 34625 7750
rect 36127 7716 36161 7750
rect 36895 7716 36929 7750
rect 33823 7568 33857 7602
rect 8383 7494 8417 7528
rect 9359 7494 9393 7528
rect 13871 7494 13905 7528
rect 28927 7494 28961 7528
rect 35359 7568 35393 7602
rect 34015 7494 34049 7528
rect 46687 7790 46721 7824
rect 46783 7790 46817 7824
rect 38815 7716 38849 7750
rect 39583 7716 39617 7750
rect 40351 7716 40385 7750
rect 41119 7716 41153 7750
rect 41887 7716 41921 7750
rect 42655 7716 42689 7750
rect 44767 7716 44801 7750
rect 45535 7716 45569 7750
rect 45823 7716 45857 7750
rect 47935 7716 47969 7750
rect 49375 7716 49409 7750
rect 50143 7716 50177 7750
rect 51007 7716 51041 7750
rect 51583 7716 51617 7750
rect 51775 7716 51809 7750
rect 53407 7716 53441 7750
rect 48991 7642 49025 7676
rect 49279 7642 49313 7676
rect 51103 7642 51137 7676
rect 53119 7642 53153 7676
rect 53311 7642 53345 7676
rect 55135 7642 55169 7676
rect 55807 7642 55841 7676
rect 56575 7642 56609 7676
rect 57343 7642 57377 7676
rect 44095 7568 44129 7602
rect 45823 7568 45857 7602
rect 46015 7568 46049 7602
rect 46303 7568 46337 7602
rect 46687 7568 46721 7602
rect 47071 7568 47105 7602
rect 47839 7568 47873 7602
rect 52639 7568 52673 7602
rect 37087 7494 37121 7528
rect 2431 7420 2465 7454
rect 3199 7420 3233 7454
rect 3967 7420 4001 7454
rect 4735 7420 4769 7454
rect 5503 7420 5537 7454
rect 7615 7420 7649 7454
rect 10111 7420 10145 7454
rect 10879 7420 10913 7454
rect 12415 7420 12449 7454
rect 13087 7420 13121 7454
rect 15871 7420 15905 7454
rect 20863 7420 20897 7454
rect 23839 7420 23873 7454
rect 24607 7420 24641 7454
rect 25375 7420 25409 7454
rect 26239 7420 26273 7454
rect 26911 7420 26945 7454
rect 28351 7420 28385 7454
rect 29311 7420 29345 7454
rect 30079 7420 30113 7454
rect 31231 7420 31265 7454
rect 33727 7420 33761 7454
rect 34495 7420 34529 7454
rect 35263 7420 35297 7454
rect 36031 7420 36065 7454
rect 36799 7420 36833 7454
rect 38719 7420 38753 7454
rect 39487 7420 39521 7454
rect 40255 7420 40289 7454
rect 41023 7420 41057 7454
rect 41791 7420 41825 7454
rect 42559 7420 42593 7454
rect 43999 7420 44033 7454
rect 44863 7420 44897 7454
rect 45631 7420 45665 7454
rect 46399 7420 46433 7454
rect 47167 7420 47201 7454
rect 47647 7420 47681 7454
rect 50047 7420 50081 7454
rect 51871 7420 51905 7454
rect 52543 7420 52577 7454
rect 5215 7198 5249 7232
rect 7519 7198 7553 7232
rect 25375 7124 25409 7158
rect 27119 7124 27153 7158
rect 31327 7124 31361 7158
rect 31903 7124 31937 7158
rect 41423 7124 41457 7158
rect 42959 7124 42993 7158
rect 51679 7124 51713 7158
rect 5023 7050 5057 7084
rect 5311 7050 5345 7084
rect 6559 7050 6593 7084
rect 6847 7050 6881 7084
rect 11935 7050 11969 7084
rect 12223 7050 12257 7084
rect 20095 7050 20129 7084
rect 21151 7050 21185 7084
rect 21631 7050 21665 7084
rect 21919 7050 21953 7084
rect 22687 7050 22721 7084
rect 24223 7050 24257 7084
rect 26431 7050 26465 7084
rect 27199 7050 27233 7084
rect 28735 7050 28769 7084
rect 29503 7050 29537 7084
rect 30943 7050 30977 7084
rect 31615 7050 31649 7084
rect 32191 7050 32225 7084
rect 32479 7050 32513 7084
rect 32959 7050 32993 7084
rect 33247 7050 33281 7084
rect 34783 7050 34817 7084
rect 36991 7050 37025 7084
rect 39295 7050 39329 7084
rect 42271 7050 42305 7084
rect 44287 7050 44321 7084
rect 44479 7050 44513 7084
rect 48319 7050 48353 7084
rect 50047 7050 50081 7084
rect 50239 7050 50273 7084
rect 51967 7050 52001 7084
rect 1663 6976 1697 7010
rect 2527 6976 2561 7010
rect 7615 6976 7649 7010
rect 9823 6976 9857 7010
rect 10015 6976 10049 7010
rect 11263 6976 11297 7010
rect 12703 6976 12737 7010
rect 36223 6976 36257 7010
rect 41215 6976 41249 7010
rect 41503 6976 41537 7010
rect 43039 6976 43073 7010
rect 43807 6976 43841 7010
rect 45263 6976 45297 7010
rect 49087 6976 49121 7010
rect 54079 6976 54113 7010
rect 54751 6976 54785 7010
rect 55519 6976 55553 7010
rect 57823 6976 57857 7010
rect 4447 6902 4481 6936
rect 4543 6902 4577 6936
rect 5983 6902 6017 6936
rect 6079 6902 6113 6936
rect 6751 6902 6785 6936
rect 8287 6902 8321 6936
rect 8383 6902 8417 6936
rect 9727 6902 9761 6936
rect 10495 6902 10529 6936
rect 10591 6902 10625 6936
rect 13567 6902 13601 6936
rect 13663 6902 13697 6936
rect 15007 6902 15041 6936
rect 15103 6902 15137 6936
rect 15775 6902 15809 6936
rect 15871 6902 15905 6936
rect 17215 6902 17249 6936
rect 17311 6902 17345 6936
rect 17791 6902 17825 6936
rect 17983 6902 18017 6936
rect 18079 6902 18113 6936
rect 18751 6902 18785 6936
rect 18847 6902 18881 6936
rect 20287 6902 20321 6936
rect 20383 6902 20417 6936
rect 21055 6902 21089 6936
rect 21823 6902 21857 6936
rect 22591 6902 22625 6936
rect 23359 6902 23393 6936
rect 23455 6902 23489 6936
rect 24127 6902 24161 6936
rect 25567 6902 25601 6936
rect 25663 6902 25697 6936
rect 26335 6902 26369 6936
rect 27871 6902 27905 6936
rect 27967 6902 28001 6936
rect 28639 6902 28673 6936
rect 29423 6902 29457 6936
rect 30847 6902 30881 6936
rect 31711 6902 31745 6936
rect 32383 6902 32417 6936
rect 33151 6902 33185 6936
rect 33919 6902 33953 6936
rect 34015 6902 34049 6936
rect 34687 6902 34721 6936
rect 36127 6902 36161 6936
rect 36895 6902 36929 6936
rect 37663 6902 37697 6936
rect 37759 6902 37793 6936
rect 38431 6902 38465 6936
rect 38527 6902 38561 6936
rect 39199 6902 39233 6936
rect 39967 6902 40001 6936
rect 40063 6902 40097 6936
rect 42175 6902 42209 6936
rect 43711 6902 43745 6936
rect 44575 6902 44609 6936
rect 45343 6902 45377 6936
rect 46687 6902 46721 6936
rect 46783 6902 46817 6936
rect 47455 6902 47489 6936
rect 47551 6902 47585 6936
rect 48223 6902 48257 6936
rect 48991 6902 49025 6936
rect 50335 6902 50369 6936
rect 52063 6902 52097 6936
rect 52735 6902 52769 6936
rect 52831 6902 52865 6936
rect 8095 6828 8129 6862
rect 10015 6828 10049 6862
rect 10303 6828 10337 6862
rect 18559 6754 18593 6788
rect 33727 6754 33761 6788
rect 46399 6754 46433 6788
rect 47167 6754 47201 6788
rect 6847 6532 6881 6566
rect 13567 6532 13601 6566
rect 28735 6532 28769 6566
rect 36895 6532 36929 6566
rect 44575 6532 44609 6566
rect 51295 6532 51329 6566
rect 7615 6458 7649 6492
rect 18175 6458 18209 6492
rect 5695 6384 5729 6418
rect 7135 6384 7169 6418
rect 13855 6384 13889 6418
rect 14719 6384 14753 6418
rect 15103 6384 15137 6418
rect 15487 6384 15521 6418
rect 16255 6384 16289 6418
rect 17599 6384 17633 6418
rect 1567 6310 1601 6344
rect 2335 6310 2369 6344
rect 3199 6310 3233 6344
rect 3967 6310 4001 6344
rect 4735 6310 4769 6344
rect 9439 6310 9473 6344
rect 10207 6310 10241 6344
rect 10975 6310 11009 6344
rect 12223 6310 12257 6344
rect 13087 6310 13121 6344
rect 27775 6458 27809 6492
rect 18463 6384 18497 6418
rect 19711 6384 19745 6418
rect 19999 6384 20033 6418
rect 24511 6384 24545 6418
rect 28447 6458 28481 6492
rect 27967 6384 28001 6418
rect 28255 6384 28289 6418
rect 19231 6310 19265 6344
rect 20687 6310 20721 6344
rect 25663 6310 25697 6344
rect 26815 6310 26849 6344
rect 27775 6310 27809 6344
rect 36223 6458 36257 6492
rect 29023 6384 29057 6418
rect 30367 6384 30401 6418
rect 30655 6384 30689 6418
rect 31903 6384 31937 6418
rect 32095 6384 32129 6418
rect 32383 6384 32417 6418
rect 34303 6384 34337 6418
rect 34687 6384 34721 6418
rect 34975 6384 35009 6418
rect 36031 6384 36065 6418
rect 29695 6310 29729 6344
rect 31231 6310 31265 6344
rect 32767 6310 32801 6344
rect 17695 6236 17729 6270
rect 18175 6236 18209 6270
rect 20767 6236 20801 6270
rect 21535 6236 21569 6270
rect 22975 6236 23009 6270
rect 23743 6236 23777 6270
rect 28447 6236 28481 6270
rect 29599 6236 29633 6270
rect 17407 6162 17441 6196
rect 33247 6236 33281 6270
rect 33439 6236 33473 6270
rect 33727 6236 33761 6270
rect 36031 6236 36065 6270
rect 37183 6384 37217 6418
rect 41311 6384 41345 6418
rect 44095 6384 44129 6418
rect 44767 6384 44801 6418
rect 50911 6384 50945 6418
rect 51583 6384 51617 6418
rect 52159 6384 52193 6418
rect 52351 6384 52385 6418
rect 36319 6310 36353 6344
rect 38911 6310 38945 6344
rect 40351 6310 40385 6344
rect 41887 6310 41921 6344
rect 45535 6310 45569 6344
rect 46975 6310 47009 6344
rect 47743 6310 47777 6344
rect 49183 6310 49217 6344
rect 49951 6310 49985 6344
rect 53311 6310 53345 6344
rect 54463 6310 54497 6344
rect 55231 6310 55265 6344
rect 55999 6310 56033 6344
rect 57055 6310 57089 6344
rect 57823 6310 57857 6344
rect 36223 6236 36257 6270
rect 42463 6236 42497 6270
rect 42751 6236 42785 6270
rect 43711 6236 43745 6270
rect 43999 6236 44033 6270
rect 46303 6236 46337 6270
rect 46111 6162 46145 6196
rect 5599 6088 5633 6122
rect 7039 6088 7073 6122
rect 13951 6088 13985 6122
rect 14623 6088 14657 6122
rect 15391 6088 15425 6122
rect 16159 6088 16193 6122
rect 18367 6088 18401 6122
rect 19135 6088 19169 6122
rect 19903 6088 19937 6122
rect 21439 6088 21473 6122
rect 22879 6088 22913 6122
rect 23647 6088 23681 6122
rect 24415 6088 24449 6122
rect 28159 6088 28193 6122
rect 28927 6088 28961 6122
rect 29599 6088 29633 6122
rect 30559 6088 30593 6122
rect 32191 6088 32225 6122
rect 32767 6088 32801 6122
rect 33535 6088 33569 6122
rect 34207 6088 34241 6122
rect 35071 6088 35105 6122
rect 37279 6088 37313 6122
rect 41215 6088 41249 6122
rect 42847 6088 42881 6122
rect 44863 6088 44897 6122
rect 50815 6088 50849 6122
rect 51679 6088 51713 6122
rect 52447 6088 52481 6122
rect 55039 5866 55073 5900
rect 55423 5866 55457 5900
rect 5791 5718 5825 5752
rect 6079 5718 6113 5752
rect 1567 5644 1601 5678
rect 2911 5644 2945 5678
rect 4447 5644 4481 5678
rect 5215 5644 5249 5678
rect 6847 5644 6881 5678
rect 7615 5644 7649 5678
rect 8383 5644 8417 5678
rect 9631 5644 9665 5678
rect 10399 5644 10433 5678
rect 11167 5644 11201 5678
rect 12607 5644 12641 5678
rect 13375 5644 13409 5678
rect 15007 5644 15041 5678
rect 15871 5644 15905 5678
rect 16543 5644 16577 5678
rect 17407 5644 17441 5678
rect 18751 5644 18785 5678
rect 20191 5644 20225 5678
rect 20959 5644 20993 5678
rect 21727 5644 21761 5678
rect 22495 5644 22529 5678
rect 23263 5644 23297 5678
rect 24031 5644 24065 5678
rect 25471 5644 25505 5678
rect 26239 5644 26273 5678
rect 27007 5644 27041 5678
rect 27775 5644 27809 5678
rect 28543 5644 28577 5678
rect 29311 5644 29345 5678
rect 30751 5644 30785 5678
rect 31519 5644 31553 5678
rect 32287 5644 32321 5678
rect 33151 5644 33185 5678
rect 33823 5644 33857 5678
rect 34687 5644 34721 5678
rect 36031 5644 36065 5678
rect 36799 5644 36833 5678
rect 37567 5644 37601 5678
rect 38335 5644 38369 5678
rect 39103 5644 39137 5678
rect 39871 5644 39905 5678
rect 41311 5644 41345 5678
rect 42079 5644 42113 5678
rect 42847 5644 42881 5678
rect 43615 5644 43649 5678
rect 44383 5644 44417 5678
rect 45151 5644 45185 5678
rect 46591 5644 46625 5678
rect 47359 5644 47393 5678
rect 48127 5644 48161 5678
rect 48991 5644 49025 5678
rect 49663 5644 49697 5678
rect 50527 5644 50561 5678
rect 52159 5644 52193 5678
rect 52927 5644 52961 5678
rect 53695 5644 53729 5678
rect 54463 5644 54497 5678
rect 55999 5644 56033 5678
rect 57439 5644 57473 5678
rect 5983 5570 6017 5604
rect 12127 5422 12161 5456
rect 7519 5200 7553 5234
rect 7711 5200 7745 5234
rect 8383 5126 8417 5160
rect 1567 4978 1601 5012
rect 2335 4978 2369 5012
rect 3103 4978 3137 5012
rect 4159 4978 4193 5012
rect 5407 4978 5441 5012
rect 6943 4978 6977 5012
rect 9247 4978 9281 5012
rect 10111 4978 10145 5012
rect 10879 4978 10913 5012
rect 12223 4978 12257 5012
rect 12991 4978 13025 5012
rect 13951 4978 13985 5012
rect 14719 4978 14753 5012
rect 15487 4978 15521 5012
rect 16351 4978 16385 5012
rect 17503 4978 17537 5012
rect 18271 4978 18305 5012
rect 19039 4978 19073 5012
rect 19807 4978 19841 5012
rect 20575 4978 20609 5012
rect 21343 4978 21377 5012
rect 22783 4978 22817 5012
rect 23551 4978 23585 5012
rect 24319 4978 24353 5012
rect 25087 4978 25121 5012
rect 25855 4978 25889 5012
rect 26623 4978 26657 5012
rect 28063 4978 28097 5012
rect 28927 4978 28961 5012
rect 29599 4978 29633 5012
rect 30367 4978 30401 5012
rect 31135 4978 31169 5012
rect 31903 4978 31937 5012
rect 33343 4978 33377 5012
rect 34111 4978 34145 5012
rect 34879 4978 34913 5012
rect 35647 4978 35681 5012
rect 36415 4978 36449 5012
rect 37183 4978 37217 5012
rect 38623 4978 38657 5012
rect 39391 4978 39425 5012
rect 40159 4978 40193 5012
rect 40927 4978 40961 5012
rect 41695 4978 41729 5012
rect 42463 4978 42497 5012
rect 43903 4978 43937 5012
rect 44767 4978 44801 5012
rect 45439 4978 45473 5012
rect 46207 4978 46241 5012
rect 46975 4978 47009 5012
rect 47743 4978 47777 5012
rect 49375 4978 49409 5012
rect 50431 4978 50465 5012
rect 51103 4978 51137 5012
rect 51871 4978 51905 5012
rect 52639 4978 52673 5012
rect 54463 4978 54497 5012
rect 55615 4978 55649 5012
rect 56383 4978 56417 5012
rect 57055 4978 57089 5012
rect 57727 4756 57761 4790
rect 57823 4756 57857 4790
rect 15775 4534 15809 4568
rect 44095 4534 44129 4568
rect 16543 4460 16577 4494
rect 17311 4460 17345 4494
rect 44287 4386 44321 4420
rect 1567 4312 1601 4346
rect 2335 4312 2369 4346
rect 3103 4312 3137 4346
rect 4351 4312 4385 4346
rect 5119 4312 5153 4346
rect 5887 4312 5921 4346
rect 6655 4312 6689 4346
rect 7423 4312 7457 4346
rect 8191 4312 8225 4346
rect 9631 4312 9665 4346
rect 10399 4312 10433 4346
rect 11167 4312 11201 4346
rect 11935 4312 11969 4346
rect 12703 4312 12737 4346
rect 13567 4312 13601 4346
rect 15487 4312 15521 4346
rect 16255 4312 16289 4346
rect 17023 4312 17057 4346
rect 17791 4312 17825 4346
rect 18559 4312 18593 4346
rect 20287 4312 20321 4346
rect 21055 4312 21089 4346
rect 21823 4312 21857 4346
rect 23263 4312 23297 4346
rect 24031 4312 24065 4346
rect 25471 4312 25505 4346
rect 26239 4312 26273 4346
rect 27007 4312 27041 4346
rect 28351 4312 28385 4346
rect 29119 4312 29153 4346
rect 30943 4312 30977 4346
rect 31711 4312 31745 4346
rect 32767 4312 32801 4346
rect 33919 4312 33953 4346
rect 34687 4312 34721 4346
rect 36031 4312 36065 4346
rect 36799 4312 36833 4346
rect 37567 4312 37601 4346
rect 39007 4312 39041 4346
rect 39775 4312 39809 4346
rect 41983 4312 42017 4346
rect 42751 4312 42785 4346
rect 43519 4312 43553 4346
rect 44959 4312 44993 4346
rect 46783 4312 46817 4346
rect 47551 4312 47585 4346
rect 48319 4312 48353 4346
rect 49087 4312 49121 4346
rect 49855 4312 49889 4346
rect 50623 4312 50657 4346
rect 51871 4312 51905 4346
rect 52639 4312 52673 4346
rect 53407 4312 53441 4346
rect 54175 4312 54209 4346
rect 55615 4312 55649 4346
rect 57247 4312 57281 4346
rect 22783 4238 22817 4272
rect 55135 4164 55169 4198
rect 19327 3868 19361 3902
rect 10687 3794 10721 3828
rect 1567 3646 1601 3680
rect 2335 3646 2369 3680
rect 3103 3646 3137 3680
rect 3871 3646 3905 3680
rect 4639 3646 4673 3680
rect 5599 3646 5633 3680
rect 6943 3646 6977 3680
rect 7711 3646 7745 3680
rect 8479 3646 8513 3680
rect 9247 3646 9281 3680
rect 10015 3646 10049 3680
rect 24223 3794 24257 3828
rect 15487 3720 15521 3754
rect 10783 3646 10817 3680
rect 12991 3646 13025 3680
rect 13663 3646 13697 3680
rect 14431 3646 14465 3680
rect 15199 3646 15233 3680
rect 15967 3646 16001 3680
rect 17503 3646 17537 3680
rect 18271 3646 18305 3680
rect 19039 3646 19073 3680
rect 19807 3646 19841 3680
rect 20575 3646 20609 3680
rect 21343 3646 21377 3680
rect 22783 3646 22817 3680
rect 23551 3646 23585 3680
rect 24319 3646 24353 3680
rect 25087 3646 25121 3680
rect 25855 3646 25889 3680
rect 26623 3646 26657 3680
rect 28063 3646 28097 3680
rect 28831 3646 28865 3680
rect 29599 3646 29633 3680
rect 30367 3646 30401 3680
rect 31135 3646 31169 3680
rect 31903 3646 31937 3680
rect 33343 3646 33377 3680
rect 34111 3646 34145 3680
rect 34879 3646 34913 3680
rect 35647 3646 35681 3680
rect 36415 3646 36449 3680
rect 37183 3646 37217 3680
rect 38623 3646 38657 3680
rect 39391 3646 39425 3680
rect 40159 3646 40193 3680
rect 40927 3646 40961 3680
rect 41695 3646 41729 3680
rect 42463 3646 42497 3680
rect 43903 3646 43937 3680
rect 44671 3646 44705 3680
rect 45439 3646 45473 3680
rect 46207 3646 46241 3680
rect 46975 3646 47009 3680
rect 47743 3646 47777 3680
rect 49183 3646 49217 3680
rect 50527 3646 50561 3680
rect 51199 3646 51233 3680
rect 51967 3646 52001 3680
rect 52735 3646 52769 3680
rect 54463 3646 54497 3680
rect 55231 3646 55265 3680
rect 55999 3646 56033 3680
rect 56767 3646 56801 3680
rect 57535 3646 57569 3680
rect 10687 3572 10721 3606
rect 12415 3572 12449 3606
rect 24223 3572 24257 3606
rect 14719 3498 14753 3532
rect 17791 3424 17825 3458
rect 20863 3424 20897 3458
rect 12703 3202 12737 3236
rect 14047 3202 14081 3236
rect 15391 3202 15425 3236
rect 16831 3202 16865 3236
rect 19135 3202 19169 3236
rect 19327 3202 19361 3236
rect 48511 3202 48545 3236
rect 13279 3128 13313 3162
rect 18847 3128 18881 3162
rect 20767 3128 20801 3162
rect 35359 3128 35393 3162
rect 35647 3128 35681 3162
rect 12703 3054 12737 3088
rect 1567 2980 1601 3014
rect 2335 2980 2369 3014
rect 3103 2980 3137 3014
rect 4927 2980 4961 3014
rect 5695 2980 5729 3014
rect 7039 2980 7073 3014
rect 7807 2980 7841 3014
rect 9727 2980 9761 3014
rect 10591 2980 10625 3014
rect 12991 2980 13025 3014
rect 13759 2980 13793 3014
rect 15103 2980 15137 3014
rect 16639 2980 16673 3014
rect 17791 2980 17825 3014
rect 18559 2980 18593 3014
rect 20479 2980 20513 3014
rect 21247 2980 21281 3014
rect 23167 2980 23201 3014
rect 23935 2980 23969 3014
rect 25855 2980 25889 3014
rect 26623 2980 26657 3014
rect 28543 2980 28577 3014
rect 29311 2980 29345 3014
rect 31231 2980 31265 3014
rect 31999 2980 32033 3014
rect 33919 2980 33953 3014
rect 34687 2980 34721 3014
rect 36607 2980 36641 3014
rect 37375 2980 37409 3014
rect 39295 2980 39329 3014
rect 40063 2980 40097 3014
rect 41983 2980 42017 3014
rect 42751 2980 42785 3014
rect 44671 2980 44705 3014
rect 45439 2980 45473 3014
rect 47359 2980 47393 3014
rect 48127 2980 48161 3014
rect 21535 2906 21569 2940
rect 46399 2832 46433 2866
rect 51775 3054 51809 3088
rect 56767 3054 56801 3088
rect 56959 3054 56993 3088
rect 50047 2980 50081 3014
rect 50815 2980 50849 3014
rect 52735 2980 52769 3014
rect 53503 2980 53537 3014
rect 55423 2980 55457 3014
rect 56191 2980 56225 3014
rect 22207 2758 22241 2792
rect 43711 2758 43745 2792
rect 48511 2758 48545 2792
rect 54463 2758 54497 2792
<< metal1 >>
rect 43984 57361 43990 57413
rect 44042 57401 44048 57413
rect 54544 57401 54550 57413
rect 44042 57373 54550 57401
rect 44042 57361 44048 57373
rect 54544 57361 54550 57373
rect 54602 57361 54608 57413
rect 1152 57302 58848 57324
rect 1152 57250 4294 57302
rect 4346 57250 4358 57302
rect 4410 57250 4422 57302
rect 4474 57250 4486 57302
rect 4538 57250 35014 57302
rect 35066 57250 35078 57302
rect 35130 57250 35142 57302
rect 35194 57250 35206 57302
rect 35258 57250 58848 57302
rect 1152 57228 58848 57250
rect 16624 57139 16630 57191
rect 16682 57179 16688 57191
rect 56755 57182 56813 57188
rect 56755 57179 56767 57182
rect 16682 57151 56767 57179
rect 16682 57139 16688 57151
rect 56755 57148 56767 57151
rect 56801 57148 56813 57182
rect 56755 57142 56813 57148
rect 1744 56991 1750 57043
rect 1802 57031 1808 57043
rect 1802 57003 2846 57031
rect 1802 56991 1808 57003
rect 208 56917 214 56969
rect 266 56957 272 56969
rect 2818 56966 2846 57003
rect 3280 56991 3286 57043
rect 3338 57031 3344 57043
rect 3338 57003 5822 57031
rect 3338 56991 3344 57003
rect 1939 56960 1997 56966
rect 1939 56957 1951 56960
rect 266 56929 1951 56957
rect 266 56917 272 56929
rect 1939 56926 1951 56929
rect 1985 56926 1997 56960
rect 1939 56920 1997 56926
rect 2803 56960 2861 56966
rect 2803 56926 2815 56960
rect 2849 56926 2861 56960
rect 2803 56920 2861 56926
rect 4912 56917 4918 56969
rect 4970 56957 4976 56969
rect 5794 56966 5822 57003
rect 9616 56991 9622 57043
rect 9674 57031 9680 57043
rect 9907 57034 9965 57040
rect 9907 57031 9919 57034
rect 9674 57003 9919 57031
rect 9674 56991 9680 57003
rect 9907 57000 9919 57003
rect 9953 57000 9965 57034
rect 9907 56994 9965 57000
rect 11248 56991 11254 57043
rect 11306 57031 11312 57043
rect 13939 57034 13997 57040
rect 11306 57003 11486 57031
rect 11306 56991 11312 57003
rect 5299 56960 5357 56966
rect 5299 56957 5311 56960
rect 4970 56929 5311 56957
rect 4970 56917 4976 56929
rect 5299 56926 5311 56929
rect 5345 56926 5357 56960
rect 5299 56920 5357 56926
rect 5779 56960 5837 56966
rect 5779 56926 5791 56960
rect 5825 56926 5837 56960
rect 5779 56920 5837 56926
rect 6448 56917 6454 56969
rect 6506 56957 6512 56969
rect 7411 56960 7469 56966
rect 7411 56957 7423 56960
rect 6506 56929 7423 56957
rect 6506 56917 6512 56929
rect 7411 56926 7423 56929
rect 7457 56926 7469 56960
rect 8080 56957 8086 56969
rect 8041 56929 8086 56957
rect 7411 56920 7469 56926
rect 8080 56917 8086 56929
rect 8138 56917 8144 56969
rect 11458 56966 11486 57003
rect 13939 57000 13951 57034
rect 13985 57031 13997 57034
rect 16432 57031 16438 57043
rect 13985 57003 16438 57031
rect 13985 57000 13997 57003
rect 13939 56994 13997 57000
rect 16432 56991 16438 57003
rect 16490 56991 16496 57043
rect 29104 56991 29110 57043
rect 29162 57031 29168 57043
rect 32563 57034 32621 57040
rect 32563 57031 32575 57034
rect 29162 57003 32575 57031
rect 29162 56991 29168 57003
rect 32563 57000 32575 57003
rect 32609 57000 32621 57034
rect 32563 56994 32621 57000
rect 39472 56991 39478 57043
rect 39530 57031 39536 57043
rect 43792 57031 43798 57043
rect 39530 57003 43798 57031
rect 39530 56991 39536 57003
rect 43792 56991 43798 57003
rect 43850 56991 43856 57043
rect 44080 56991 44086 57043
rect 44138 57031 44144 57043
rect 52048 57031 52054 57043
rect 44138 57003 52054 57031
rect 44138 56991 44144 57003
rect 52048 56991 52054 57003
rect 52106 56991 52112 57043
rect 11443 56960 11501 56966
rect 11443 56926 11455 56960
rect 11489 56926 11501 56960
rect 11443 56920 11501 56926
rect 12784 56917 12790 56969
rect 12842 56957 12848 56969
rect 13171 56960 13229 56966
rect 13171 56957 13183 56960
rect 12842 56929 13183 56957
rect 12842 56917 12848 56929
rect 13171 56926 13183 56929
rect 13217 56926 13229 56960
rect 13171 56920 13229 56926
rect 14416 56917 14422 56969
rect 14474 56957 14480 56969
rect 15091 56960 15149 56966
rect 15091 56957 15103 56960
rect 14474 56929 15103 56957
rect 14474 56917 14480 56929
rect 15091 56926 15103 56929
rect 15137 56926 15149 56960
rect 15091 56920 15149 56926
rect 15952 56917 15958 56969
rect 16010 56957 16016 56969
rect 16339 56960 16397 56966
rect 16339 56957 16351 56960
rect 16010 56929 16351 56957
rect 16010 56917 16016 56929
rect 16339 56926 16351 56929
rect 16385 56926 16397 56960
rect 16339 56920 16397 56926
rect 17488 56917 17494 56969
rect 17546 56957 17552 56969
rect 18163 56960 18221 56966
rect 18163 56957 18175 56960
rect 17546 56929 18175 56957
rect 17546 56917 17552 56929
rect 18163 56926 18175 56929
rect 18209 56926 18221 56960
rect 18163 56920 18221 56926
rect 19120 56917 19126 56969
rect 19178 56957 19184 56969
rect 19507 56960 19565 56966
rect 19507 56957 19519 56960
rect 19178 56929 19519 56957
rect 19178 56917 19184 56929
rect 19507 56926 19519 56929
rect 19553 56926 19565 56960
rect 19507 56920 19565 56926
rect 20656 56917 20662 56969
rect 20714 56957 20720 56969
rect 21043 56960 21101 56966
rect 21043 56957 21055 56960
rect 20714 56929 21055 56957
rect 20714 56917 20720 56929
rect 21043 56926 21055 56929
rect 21089 56926 21101 56960
rect 21043 56920 21101 56926
rect 22003 56960 22061 56966
rect 22003 56926 22015 56960
rect 22049 56957 22061 56960
rect 22288 56957 22294 56969
rect 22049 56929 22294 56957
rect 22049 56926 22061 56929
rect 22003 56920 22061 56926
rect 22288 56917 22294 56929
rect 22346 56917 22352 56969
rect 23824 56917 23830 56969
rect 23882 56957 23888 56969
rect 24211 56960 24269 56966
rect 24211 56957 24223 56960
rect 23882 56929 24223 56957
rect 23882 56917 23888 56929
rect 24211 56926 24223 56929
rect 24257 56926 24269 56960
rect 24211 56920 24269 56926
rect 25456 56917 25462 56969
rect 25514 56957 25520 56969
rect 25939 56960 25997 56966
rect 25939 56957 25951 56960
rect 25514 56929 25951 56957
rect 25514 56917 25520 56929
rect 25939 56926 25951 56929
rect 25985 56926 25997 56960
rect 25939 56920 25997 56926
rect 26992 56917 26998 56969
rect 27050 56957 27056 56969
rect 27379 56960 27437 56966
rect 27379 56957 27391 56960
rect 27050 56929 27391 56957
rect 27050 56917 27056 56929
rect 27379 56926 27391 56929
rect 27425 56926 27437 56960
rect 28624 56957 28630 56969
rect 28585 56929 28630 56957
rect 27379 56920 27437 56926
rect 28624 56917 28630 56929
rect 28682 56917 28688 56969
rect 30256 56957 30262 56969
rect 30217 56929 30262 56957
rect 30256 56917 30262 56929
rect 30314 56917 30320 56969
rect 31696 56957 31702 56969
rect 31657 56929 31702 56957
rect 31696 56917 31702 56929
rect 31754 56917 31760 56969
rect 33328 56917 33334 56969
rect 33386 56957 33392 56969
rect 34291 56960 34349 56966
rect 34291 56957 34303 56960
rect 33386 56929 34303 56957
rect 33386 56917 33392 56929
rect 34291 56926 34303 56929
rect 34337 56926 34349 56960
rect 34864 56957 34870 56969
rect 34825 56929 34870 56957
rect 34291 56920 34349 56926
rect 34864 56917 34870 56929
rect 34922 56917 34928 56969
rect 38032 56957 38038 56969
rect 37993 56929 38038 56957
rect 38032 56917 38038 56929
rect 38090 56917 38096 56969
rect 38128 56917 38134 56969
rect 38186 56957 38192 56969
rect 38186 56929 40862 56957
rect 38186 56917 38192 56929
rect 1744 56883 1750 56895
rect 1705 56855 1750 56883
rect 1744 56843 1750 56855
rect 1802 56843 1808 56895
rect 2611 56886 2669 56892
rect 2611 56852 2623 56886
rect 2657 56883 2669 56886
rect 3568 56883 3574 56895
rect 2657 56855 3574 56883
rect 2657 56852 2669 56855
rect 2611 56846 2669 56852
rect 3568 56843 3574 56855
rect 3626 56843 3632 56895
rect 5104 56883 5110 56895
rect 5065 56855 5110 56883
rect 5104 56843 5110 56855
rect 5162 56843 5168 56895
rect 7219 56886 7277 56892
rect 7219 56852 7231 56886
rect 7265 56883 7277 56886
rect 8272 56883 8278 56895
rect 7265 56855 8278 56883
rect 7265 56852 7277 56855
rect 7219 56846 7277 56852
rect 8272 56843 8278 56855
rect 8330 56843 8336 56895
rect 11248 56883 11254 56895
rect 11209 56855 11254 56883
rect 11248 56843 11254 56855
rect 11306 56843 11312 56895
rect 12976 56883 12982 56895
rect 12937 56855 12982 56883
rect 12976 56843 12982 56855
rect 13034 56843 13040 56895
rect 14035 56886 14093 56892
rect 14035 56852 14047 56886
rect 14081 56883 14093 56886
rect 15568 56883 15574 56895
rect 14081 56855 15574 56883
rect 14081 56852 14093 56855
rect 14035 56846 14093 56852
rect 15568 56843 15574 56855
rect 15626 56843 15632 56895
rect 16144 56883 16150 56895
rect 16105 56855 16150 56883
rect 16144 56843 16150 56855
rect 16202 56843 16208 56895
rect 17968 56883 17974 56895
rect 17929 56855 17974 56883
rect 17968 56843 17974 56855
rect 18026 56843 18032 56895
rect 19312 56883 19318 56895
rect 19273 56855 19318 56883
rect 19312 56843 19318 56855
rect 19370 56843 19376 56895
rect 20848 56883 20854 56895
rect 20809 56855 20854 56883
rect 20848 56843 20854 56855
rect 20906 56843 20912 56895
rect 24019 56886 24077 56892
rect 24019 56883 24031 56886
rect 22306 56855 24031 56883
rect 22306 56821 22334 56855
rect 24019 56852 24031 56855
rect 24065 56852 24077 56886
rect 24019 56846 24077 56852
rect 25168 56843 25174 56895
rect 25226 56883 25232 56895
rect 27187 56886 27245 56892
rect 27187 56883 27199 56886
rect 25226 56855 27199 56883
rect 25226 56843 25232 56855
rect 27187 56852 27199 56855
rect 27233 56852 27245 56886
rect 30064 56883 30070 56895
rect 30025 56855 30070 56883
rect 27187 56846 27245 56852
rect 30064 56843 30070 56855
rect 30122 56843 30128 56895
rect 32656 56883 32662 56895
rect 32617 56855 32662 56883
rect 32656 56843 32662 56855
rect 32714 56843 32720 56895
rect 34099 56886 34157 56892
rect 34099 56852 34111 56886
rect 34145 56852 34157 56886
rect 34099 56846 34157 56852
rect 22288 56769 22294 56821
rect 22346 56769 22352 56821
rect 25552 56769 25558 56821
rect 25610 56809 25616 56821
rect 34114 56809 34142 56846
rect 36496 56843 36502 56895
rect 36554 56883 36560 56895
rect 36979 56886 37037 56892
rect 36979 56883 36991 56886
rect 36554 56855 36991 56883
rect 36554 56843 36560 56855
rect 36979 56852 36991 56855
rect 37025 56852 37037 56886
rect 36979 56846 37037 56852
rect 39664 56843 39670 56895
rect 39722 56883 39728 56895
rect 40051 56886 40109 56892
rect 40051 56883 40063 56886
rect 39722 56855 40063 56883
rect 39722 56843 39728 56855
rect 40051 56852 40063 56855
rect 40097 56852 40109 56886
rect 40051 56846 40109 56852
rect 40723 56886 40781 56892
rect 40723 56852 40735 56886
rect 40769 56852 40781 56886
rect 40834 56883 40862 56929
rect 41200 56917 41206 56969
rect 41258 56957 41264 56969
rect 41971 56960 42029 56966
rect 41971 56957 41983 56960
rect 41258 56929 41983 56957
rect 41258 56917 41264 56929
rect 41971 56926 41983 56929
rect 42017 56926 42029 56960
rect 41971 56920 42029 56926
rect 47536 56917 47542 56969
rect 47594 56957 47600 56969
rect 47594 56929 47639 56957
rect 47594 56917 47600 56929
rect 52240 56917 52246 56969
rect 52298 56957 52304 56969
rect 52723 56960 52781 56966
rect 52723 56957 52735 56960
rect 52298 56929 52735 56957
rect 52298 56917 52304 56929
rect 52723 56926 52735 56929
rect 52769 56926 52781 56960
rect 52723 56920 52781 56926
rect 40834 56855 41342 56883
rect 40723 56846 40781 56852
rect 25610 56781 34142 56809
rect 40531 56812 40589 56818
rect 25610 56769 25616 56781
rect 40531 56778 40543 56812
rect 40577 56809 40589 56812
rect 40738 56809 40766 56846
rect 41200 56809 41206 56821
rect 40577 56781 41206 56809
rect 40577 56778 40589 56781
rect 40531 56772 40589 56778
rect 41200 56769 41206 56781
rect 41258 56769 41264 56821
rect 41314 56809 41342 56855
rect 42832 56843 42838 56895
rect 42890 56883 42896 56895
rect 43219 56886 43277 56892
rect 43219 56883 43231 56886
rect 42890 56855 43231 56883
rect 42890 56843 42896 56855
rect 43219 56852 43231 56855
rect 43265 56852 43277 56886
rect 43219 56846 43277 56852
rect 44368 56843 44374 56895
rect 44426 56883 44432 56895
rect 45043 56886 45101 56892
rect 45043 56883 45055 56886
rect 44426 56855 45055 56883
rect 44426 56843 44432 56855
rect 45043 56852 45055 56855
rect 45089 56852 45101 56886
rect 45043 56846 45101 56852
rect 45904 56843 45910 56895
rect 45962 56883 45968 56895
rect 46291 56886 46349 56892
rect 46291 56883 46303 56886
rect 45962 56855 46303 56883
rect 45962 56843 45968 56855
rect 46291 56852 46303 56855
rect 46337 56852 46349 56886
rect 46291 56846 46349 56852
rect 48979 56886 49037 56892
rect 48979 56852 48991 56886
rect 49025 56883 49037 56886
rect 49072 56883 49078 56895
rect 49025 56855 49078 56883
rect 49025 56852 49037 56855
rect 48979 56846 49037 56852
rect 49072 56843 49078 56855
rect 49130 56843 49136 56895
rect 50704 56843 50710 56895
rect 50762 56883 50768 56895
rect 51091 56886 51149 56892
rect 51091 56883 51103 56886
rect 50762 56855 51103 56883
rect 50762 56843 50768 56855
rect 51091 56852 51103 56855
rect 51137 56852 51149 56886
rect 51091 56846 51149 56852
rect 53872 56843 53878 56895
rect 53930 56883 53936 56895
rect 54259 56886 54317 56892
rect 54259 56883 54271 56886
rect 53930 56855 54271 56883
rect 53930 56843 53936 56855
rect 54259 56852 54271 56855
rect 54305 56852 54317 56886
rect 54259 56846 54317 56852
rect 55408 56843 55414 56895
rect 55466 56883 55472 56895
rect 55795 56886 55853 56892
rect 55795 56883 55807 56886
rect 55466 56855 55807 56883
rect 55466 56843 55472 56855
rect 55795 56852 55807 56855
rect 55841 56852 55853 56886
rect 57040 56883 57046 56895
rect 57001 56855 57046 56883
rect 55795 56846 55853 56852
rect 57040 56843 57046 56855
rect 57098 56843 57104 56895
rect 55312 56809 55318 56821
rect 41314 56781 55318 56809
rect 55312 56769 55318 56781
rect 55370 56769 55376 56821
rect 9712 56695 9718 56747
rect 9770 56735 9776 56747
rect 9811 56738 9869 56744
rect 9811 56735 9823 56738
rect 9770 56707 9823 56735
rect 9770 56695 9776 56707
rect 9811 56704 9823 56707
rect 9857 56704 9869 56738
rect 36688 56735 36694 56747
rect 36649 56707 36694 56735
rect 9811 56698 9869 56704
rect 36688 56695 36694 56707
rect 36746 56695 36752 56747
rect 39760 56735 39766 56747
rect 39721 56707 39766 56735
rect 39760 56695 39766 56707
rect 39818 56695 39824 56747
rect 40816 56735 40822 56747
rect 40777 56707 40822 56735
rect 40816 56695 40822 56707
rect 40874 56695 40880 56747
rect 42928 56735 42934 56747
rect 42889 56707 42934 56735
rect 42928 56695 42934 56707
rect 42986 56695 42992 56747
rect 44752 56735 44758 56747
rect 44713 56707 44758 56735
rect 44752 56695 44758 56707
rect 44810 56695 44816 56747
rect 46003 56738 46061 56744
rect 46003 56704 46015 56738
rect 46049 56735 46061 56738
rect 46096 56735 46102 56747
rect 46049 56707 46102 56735
rect 46049 56704 46061 56707
rect 46003 56698 46061 56704
rect 46096 56695 46102 56707
rect 46154 56695 46160 56747
rect 48688 56735 48694 56747
rect 48649 56707 48694 56735
rect 48688 56695 48694 56707
rect 48746 56695 48752 56747
rect 50800 56735 50806 56747
rect 50761 56707 50806 56735
rect 50800 56695 50806 56707
rect 50858 56695 50864 56747
rect 53968 56735 53974 56747
rect 53929 56707 53974 56735
rect 53968 56695 53974 56707
rect 54026 56695 54032 56747
rect 55504 56735 55510 56747
rect 55465 56707 55510 56735
rect 55504 56695 55510 56707
rect 55562 56695 55568 56747
rect 1152 56636 58848 56658
rect 1152 56584 19654 56636
rect 19706 56584 19718 56636
rect 19770 56584 19782 56636
rect 19834 56584 19846 56636
rect 19898 56584 50374 56636
rect 50426 56584 50438 56636
rect 50490 56584 50502 56636
rect 50554 56584 50566 56636
rect 50618 56584 58848 56636
rect 1152 56562 58848 56584
rect 688 56473 694 56525
rect 746 56513 752 56525
rect 1651 56516 1709 56522
rect 1651 56513 1663 56516
rect 746 56485 1663 56513
rect 746 56473 752 56485
rect 1651 56482 1663 56485
rect 1697 56482 1709 56516
rect 1651 56476 1709 56482
rect 2224 56473 2230 56525
rect 2282 56513 2288 56525
rect 2419 56516 2477 56522
rect 2419 56513 2431 56516
rect 2282 56485 2431 56513
rect 2282 56473 2288 56485
rect 2419 56482 2431 56485
rect 2465 56482 2477 56516
rect 2419 56476 2477 56482
rect 2800 56473 2806 56525
rect 2858 56513 2864 56525
rect 3187 56516 3245 56522
rect 3187 56513 3199 56516
rect 2858 56485 3199 56513
rect 2858 56473 2864 56485
rect 3187 56482 3199 56485
rect 3233 56482 3245 56516
rect 3187 56476 3245 56482
rect 3856 56473 3862 56525
rect 3914 56513 3920 56525
rect 4435 56516 4493 56522
rect 4435 56513 4447 56516
rect 3914 56485 4447 56513
rect 3914 56473 3920 56485
rect 4435 56482 4447 56485
rect 4481 56482 4493 56516
rect 4435 56476 4493 56482
rect 5392 56473 5398 56525
rect 5450 56513 5456 56525
rect 5491 56516 5549 56522
rect 5491 56513 5503 56516
rect 5450 56485 5503 56513
rect 5450 56473 5456 56485
rect 5491 56482 5503 56485
rect 5537 56482 5549 56516
rect 5491 56476 5549 56482
rect 5968 56473 5974 56525
rect 6026 56513 6032 56525
rect 6259 56516 6317 56522
rect 6259 56513 6271 56516
rect 6026 56485 6271 56513
rect 6026 56473 6032 56485
rect 6259 56482 6271 56485
rect 6305 56482 6317 56516
rect 6259 56476 6317 56482
rect 7024 56473 7030 56525
rect 7082 56513 7088 56525
rect 7123 56516 7181 56522
rect 7123 56513 7135 56516
rect 7082 56485 7135 56513
rect 7082 56473 7088 56485
rect 7123 56482 7135 56485
rect 7169 56482 7181 56516
rect 7123 56476 7181 56482
rect 8467 56516 8525 56522
rect 8467 56482 8479 56516
rect 8513 56513 8525 56516
rect 8560 56513 8566 56525
rect 8513 56485 8566 56513
rect 8513 56482 8525 56485
rect 8467 56476 8525 56482
rect 8560 56473 8566 56485
rect 8618 56473 8624 56525
rect 10192 56473 10198 56525
rect 10250 56513 10256 56525
rect 10291 56516 10349 56522
rect 10291 56513 10303 56516
rect 10250 56485 10303 56513
rect 10250 56473 10256 56485
rect 10291 56482 10303 56485
rect 10337 56482 10349 56516
rect 10291 56476 10349 56482
rect 10672 56473 10678 56525
rect 10730 56513 10736 56525
rect 11059 56516 11117 56522
rect 11059 56513 11071 56516
rect 10730 56485 11071 56513
rect 10730 56473 10736 56485
rect 11059 56482 11071 56485
rect 11105 56482 11117 56516
rect 11059 56476 11117 56482
rect 11728 56473 11734 56525
rect 11786 56513 11792 56525
rect 11827 56516 11885 56522
rect 11827 56513 11839 56516
rect 11786 56485 11839 56513
rect 11786 56473 11792 56485
rect 11827 56482 11839 56485
rect 11873 56482 11885 56516
rect 11827 56476 11885 56482
rect 12304 56473 12310 56525
rect 12362 56513 12368 56525
rect 12595 56516 12653 56522
rect 12595 56513 12607 56516
rect 12362 56485 12607 56513
rect 12362 56473 12368 56485
rect 12595 56482 12607 56485
rect 12641 56482 12653 56516
rect 12595 56476 12653 56482
rect 13360 56473 13366 56525
rect 13418 56513 13424 56525
rect 13459 56516 13517 56522
rect 13459 56513 13471 56516
rect 13418 56485 13471 56513
rect 13418 56473 13424 56485
rect 13459 56482 13471 56485
rect 13505 56482 13517 56516
rect 13459 56476 13517 56482
rect 14896 56473 14902 56525
rect 14954 56513 14960 56525
rect 15091 56516 15149 56522
rect 15091 56513 15103 56516
rect 14954 56485 15103 56513
rect 14954 56473 14960 56485
rect 15091 56482 15103 56485
rect 15137 56482 15149 56516
rect 15091 56476 15149 56482
rect 17008 56473 17014 56525
rect 17066 56513 17072 56525
rect 17203 56516 17261 56522
rect 17203 56513 17215 56516
rect 17066 56485 17215 56513
rect 17066 56473 17072 56485
rect 17203 56482 17215 56485
rect 17249 56482 17261 56516
rect 17203 56476 17261 56482
rect 18064 56473 18070 56525
rect 18122 56513 18128 56525
rect 18163 56516 18221 56522
rect 18163 56513 18175 56516
rect 18122 56485 18175 56513
rect 18122 56473 18128 56485
rect 18163 56482 18175 56485
rect 18209 56482 18221 56516
rect 18163 56476 18221 56482
rect 18544 56473 18550 56525
rect 18602 56513 18608 56525
rect 18931 56516 18989 56522
rect 18931 56513 18943 56516
rect 18602 56485 18943 56513
rect 18602 56473 18608 56485
rect 18931 56482 18943 56485
rect 18977 56482 18989 56516
rect 18931 56476 18989 56482
rect 19984 56473 19990 56525
rect 20042 56513 20048 56525
rect 20275 56516 20333 56522
rect 20275 56513 20287 56516
rect 20042 56485 20287 56513
rect 20042 56473 20048 56485
rect 20275 56482 20287 56485
rect 20321 56482 20333 56516
rect 20275 56476 20333 56482
rect 21232 56473 21238 56525
rect 21290 56513 21296 56525
rect 21427 56516 21485 56522
rect 21427 56513 21439 56516
rect 21290 56485 21439 56513
rect 21290 56473 21296 56485
rect 21427 56482 21439 56485
rect 21473 56482 21485 56516
rect 21427 56476 21485 56482
rect 21712 56473 21718 56525
rect 21770 56513 21776 56525
rect 22099 56516 22157 56522
rect 22099 56513 22111 56516
rect 21770 56485 22111 56513
rect 21770 56473 21776 56485
rect 22099 56482 22111 56485
rect 22145 56482 22157 56516
rect 22099 56476 22157 56482
rect 22768 56473 22774 56525
rect 22826 56513 22832 56525
rect 22963 56516 23021 56522
rect 22963 56513 22975 56516
rect 22826 56485 22975 56513
rect 22826 56473 22832 56485
rect 22963 56482 22975 56485
rect 23009 56482 23021 56516
rect 24400 56513 24406 56525
rect 24361 56485 24406 56513
rect 22963 56476 23021 56482
rect 24400 56473 24406 56485
rect 24458 56473 24464 56525
rect 25936 56473 25942 56525
rect 25994 56513 26000 56525
rect 26035 56516 26093 56522
rect 26035 56513 26047 56516
rect 25994 56485 26047 56513
rect 25994 56473 26000 56485
rect 26035 56482 26047 56485
rect 26081 56482 26093 56516
rect 26035 56476 26093 56482
rect 26512 56473 26518 56525
rect 26570 56513 26576 56525
rect 26899 56516 26957 56522
rect 26899 56513 26911 56516
rect 26570 56485 26911 56513
rect 26570 56473 26576 56485
rect 26899 56482 26911 56485
rect 26945 56482 26957 56516
rect 26899 56476 26957 56482
rect 27568 56473 27574 56525
rect 27626 56513 27632 56525
rect 27763 56516 27821 56522
rect 27763 56513 27775 56516
rect 27626 56485 27775 56513
rect 27626 56473 27632 56485
rect 27763 56482 27775 56485
rect 27809 56482 27821 56516
rect 27763 56476 27821 56482
rect 28048 56473 28054 56525
rect 28106 56513 28112 56525
rect 28435 56516 28493 56522
rect 28435 56513 28447 56516
rect 28106 56485 28447 56513
rect 28106 56473 28112 56485
rect 28435 56482 28447 56485
rect 28481 56482 28493 56516
rect 29680 56513 29686 56525
rect 29641 56485 29686 56513
rect 28435 56476 28493 56482
rect 29680 56473 29686 56485
rect 29738 56473 29744 56525
rect 30640 56473 30646 56525
rect 30698 56513 30704 56525
rect 30835 56516 30893 56522
rect 30835 56513 30847 56516
rect 30698 56485 30847 56513
rect 30698 56473 30704 56485
rect 30835 56482 30847 56485
rect 30881 56482 30893 56516
rect 30835 56476 30893 56482
rect 31216 56473 31222 56525
rect 31274 56513 31280 56525
rect 31603 56516 31661 56522
rect 31603 56513 31615 56516
rect 31274 56485 31615 56513
rect 31274 56473 31280 56485
rect 31603 56482 31615 56485
rect 31649 56482 31661 56516
rect 31603 56476 31661 56482
rect 32272 56473 32278 56525
rect 32330 56513 32336 56525
rect 32371 56516 32429 56522
rect 32371 56513 32383 56516
rect 32330 56485 32383 56513
rect 32330 56473 32336 56485
rect 32371 56482 32383 56485
rect 32417 56482 32429 56516
rect 32371 56476 32429 56482
rect 33808 56473 33814 56525
rect 33866 56513 33872 56525
rect 33907 56516 33965 56522
rect 33907 56513 33919 56516
rect 33866 56485 33919 56513
rect 33866 56473 33872 56485
rect 33907 56482 33919 56485
rect 33953 56482 33965 56516
rect 33907 56476 33965 56482
rect 34576 56473 34582 56525
rect 34634 56513 34640 56525
rect 34771 56516 34829 56522
rect 34771 56513 34783 56516
rect 34634 56485 34783 56513
rect 34634 56473 34640 56485
rect 34771 56482 34783 56485
rect 34817 56482 34829 56516
rect 34771 56476 34829 56482
rect 35440 56473 35446 56525
rect 35498 56513 35504 56525
rect 36115 56516 36173 56522
rect 36115 56513 36127 56516
rect 35498 56485 36127 56513
rect 35498 56473 35504 56485
rect 36115 56482 36127 56485
rect 36161 56482 36173 56516
rect 36115 56476 36173 56482
rect 36208 56473 36214 56525
rect 36266 56513 36272 56525
rect 36979 56516 37037 56522
rect 36979 56513 36991 56516
rect 36266 56485 36991 56513
rect 36266 56473 36272 56485
rect 36979 56482 36991 56485
rect 37025 56482 37037 56516
rect 36979 56476 37037 56482
rect 37552 56473 37558 56525
rect 37610 56513 37616 56525
rect 37747 56516 37805 56522
rect 37747 56513 37759 56516
rect 37610 56485 37759 56513
rect 37610 56473 37616 56485
rect 37747 56482 37759 56485
rect 37793 56482 37805 56516
rect 37747 56476 37805 56482
rect 38608 56473 38614 56525
rect 38666 56513 38672 56525
rect 38707 56516 38765 56522
rect 38707 56513 38719 56516
rect 38666 56485 38719 56513
rect 38666 56473 38672 56485
rect 38707 56482 38719 56485
rect 38753 56482 38765 56516
rect 40144 56513 40150 56525
rect 40105 56485 40150 56513
rect 38707 56476 38765 56482
rect 40144 56473 40150 56485
rect 40202 56473 40208 56525
rect 41776 56473 41782 56525
rect 41834 56513 41840 56525
rect 41875 56516 41933 56522
rect 41875 56513 41887 56516
rect 41834 56485 41887 56513
rect 41834 56473 41840 56485
rect 41875 56482 41887 56485
rect 41921 56482 41933 56516
rect 41875 56476 41933 56482
rect 42256 56473 42262 56525
rect 42314 56513 42320 56525
rect 42739 56516 42797 56522
rect 42739 56513 42751 56516
rect 42314 56485 42751 56513
rect 42314 56473 42320 56485
rect 42739 56482 42751 56485
rect 42785 56482 42797 56516
rect 42739 56476 42797 56482
rect 43312 56473 43318 56525
rect 43370 56513 43376 56525
rect 43411 56516 43469 56522
rect 43411 56513 43423 56516
rect 43370 56485 43423 56513
rect 43370 56473 43376 56485
rect 43411 56482 43423 56485
rect 43457 56482 43469 56516
rect 43411 56476 43469 56482
rect 43888 56473 43894 56525
rect 43946 56513 43952 56525
rect 44179 56516 44237 56522
rect 44179 56513 44191 56516
rect 43946 56485 44191 56513
rect 43946 56473 43952 56485
rect 44179 56482 44191 56485
rect 44225 56482 44237 56516
rect 44179 56476 44237 56482
rect 44944 56473 44950 56525
rect 45002 56513 45008 56525
rect 45043 56516 45101 56522
rect 45043 56513 45055 56516
rect 45002 56485 45055 56513
rect 45002 56473 45008 56485
rect 45043 56482 45055 56485
rect 45089 56482 45101 56516
rect 45043 56476 45101 56482
rect 46480 56473 46486 56525
rect 46538 56513 46544 56525
rect 46675 56516 46733 56522
rect 46675 56513 46687 56516
rect 46538 56485 46687 56513
rect 46538 56473 46544 56485
rect 46675 56482 46687 56485
rect 46721 56482 46733 56516
rect 46675 56476 46733 56482
rect 48016 56473 48022 56525
rect 48074 56513 48080 56525
rect 48115 56516 48173 56522
rect 48115 56513 48127 56516
rect 48074 56485 48127 56513
rect 48074 56473 48080 56485
rect 48115 56482 48127 56485
rect 48161 56482 48173 56516
rect 48115 56476 48173 56482
rect 49648 56473 49654 56525
rect 49706 56513 49712 56525
rect 49747 56516 49805 56522
rect 49747 56513 49759 56516
rect 49706 56485 49759 56513
rect 49706 56473 49712 56485
rect 49747 56482 49759 56485
rect 49793 56482 49805 56516
rect 49747 56476 49805 56482
rect 50128 56473 50134 56525
rect 50186 56513 50192 56525
rect 50515 56516 50573 56522
rect 50515 56513 50527 56516
rect 50186 56485 50527 56513
rect 50186 56473 50192 56485
rect 50515 56482 50527 56485
rect 50561 56482 50573 56516
rect 50515 56476 50573 56482
rect 51280 56473 51286 56525
rect 51338 56513 51344 56525
rect 51955 56516 52013 56522
rect 51955 56513 51967 56516
rect 51338 56485 51967 56513
rect 51338 56473 51344 56485
rect 51955 56482 51967 56485
rect 52001 56482 52013 56516
rect 51955 56476 52013 56482
rect 52816 56473 52822 56525
rect 52874 56513 52880 56525
rect 53011 56516 53069 56522
rect 53011 56513 53023 56516
rect 52874 56485 53023 56513
rect 52874 56473 52880 56485
rect 53011 56482 53023 56485
rect 53057 56482 53069 56516
rect 53011 56476 53069 56482
rect 53296 56473 53302 56525
rect 53354 56513 53360 56525
rect 53779 56516 53837 56522
rect 53779 56513 53791 56516
rect 53354 56485 53791 56513
rect 53354 56473 53360 56485
rect 53779 56482 53791 56485
rect 53825 56482 53837 56516
rect 53779 56476 53837 56482
rect 54352 56473 54358 56525
rect 54410 56513 54416 56525
rect 54451 56516 54509 56522
rect 54451 56513 54463 56516
rect 54410 56485 54463 56513
rect 54410 56473 54416 56485
rect 54451 56482 54463 56485
rect 54497 56482 54509 56516
rect 54451 56476 54509 56482
rect 54928 56473 54934 56525
rect 54986 56513 54992 56525
rect 55219 56516 55277 56522
rect 55219 56513 55231 56516
rect 54986 56485 55231 56513
rect 54986 56473 54992 56485
rect 55219 56482 55231 56485
rect 55265 56482 55277 56516
rect 55219 56476 55277 56482
rect 55984 56473 55990 56525
rect 56042 56513 56048 56525
rect 56083 56516 56141 56522
rect 56083 56513 56095 56516
rect 56042 56485 56095 56513
rect 56042 56473 56048 56485
rect 56083 56482 56095 56485
rect 56129 56482 56141 56516
rect 56083 56476 56141 56482
rect 16528 56399 16534 56451
rect 16586 56439 16592 56451
rect 48688 56439 48694 56451
rect 16586 56411 48694 56439
rect 16586 56399 16592 56411
rect 48688 56399 48694 56411
rect 48746 56399 48752 56451
rect 50323 56442 50381 56448
rect 50323 56408 50335 56442
rect 50369 56439 50381 56442
rect 51187 56442 51245 56448
rect 51187 56439 51199 56442
rect 50369 56411 51199 56439
rect 50369 56408 50381 56411
rect 50323 56402 50381 56408
rect 51187 56408 51199 56411
rect 51233 56439 51245 56442
rect 55120 56439 55126 56451
rect 51233 56411 55126 56439
rect 51233 56408 51245 56411
rect 51187 56402 51245 56408
rect 55120 56399 55126 56411
rect 55178 56399 55184 56451
rect 15280 56325 15286 56377
rect 15338 56365 15344 56377
rect 22195 56368 22253 56374
rect 22195 56365 22207 56368
rect 15338 56337 22207 56365
rect 15338 56325 15344 56337
rect 22195 56334 22207 56337
rect 22241 56334 22253 56368
rect 22195 56328 22253 56334
rect 31411 56368 31469 56374
rect 31411 56334 31423 56368
rect 31457 56365 31469 56368
rect 31699 56368 31757 56374
rect 31699 56365 31711 56368
rect 31457 56337 31711 56365
rect 31457 56334 31469 56337
rect 31411 56328 31469 56334
rect 31699 56334 31711 56337
rect 31745 56365 31757 56368
rect 39472 56365 39478 56377
rect 31745 56337 39478 56365
rect 31745 56334 31757 56337
rect 31699 56328 31757 56334
rect 39472 56325 39478 56337
rect 39530 56325 39536 56377
rect 39568 56325 39574 56377
rect 39626 56365 39632 56377
rect 41971 56368 42029 56374
rect 41971 56365 41983 56368
rect 39626 56337 41983 56365
rect 39626 56325 39632 56337
rect 41971 56334 41983 56337
rect 42017 56334 42029 56368
rect 41971 56328 42029 56334
rect 42448 56325 42454 56377
rect 42506 56365 42512 56377
rect 43507 56368 43565 56374
rect 43507 56365 43519 56368
rect 42506 56337 43519 56365
rect 42506 56325 42512 56337
rect 43507 56334 43519 56337
rect 43553 56334 43565 56368
rect 43507 56328 43565 56334
rect 43888 56325 43894 56377
rect 43946 56365 43952 56377
rect 55504 56365 55510 56377
rect 43946 56337 55510 56365
rect 43946 56325 43952 56337
rect 55504 56325 55510 56337
rect 55562 56325 55568 56377
rect 6736 56251 6742 56303
rect 6794 56291 6800 56303
rect 26131 56294 26189 56300
rect 26131 56291 26143 56294
rect 6794 56263 26143 56291
rect 6794 56251 6800 56263
rect 26131 56260 26143 56263
rect 26177 56260 26189 56294
rect 26131 56254 26189 56260
rect 30256 56251 30262 56303
rect 30314 56291 30320 56303
rect 34003 56294 34061 56300
rect 34003 56291 34015 56294
rect 30314 56263 34015 56291
rect 30314 56251 30320 56263
rect 34003 56260 34015 56263
rect 34049 56260 34061 56294
rect 34003 56254 34061 56260
rect 41296 56251 41302 56303
rect 41354 56291 41360 56303
rect 45139 56294 45197 56300
rect 45139 56291 45151 56294
rect 41354 56263 45151 56291
rect 41354 56251 41360 56263
rect 45139 56260 45151 56263
rect 45185 56260 45197 56294
rect 45139 56254 45197 56260
rect 50611 56294 50669 56300
rect 50611 56260 50623 56294
rect 50657 56291 50669 56294
rect 51187 56294 51245 56300
rect 51187 56291 51199 56294
rect 50657 56263 51199 56291
rect 50657 56260 50669 56263
rect 50611 56254 50669 56260
rect 51187 56260 51199 56263
rect 51233 56260 51245 56294
rect 52048 56291 52054 56303
rect 52009 56263 52054 56291
rect 51187 56254 51245 56260
rect 52048 56251 52054 56263
rect 52106 56251 52112 56303
rect 54544 56291 54550 56303
rect 52162 56263 53822 56291
rect 54505 56263 54550 56291
rect 1747 56220 1805 56226
rect 1747 56186 1759 56220
rect 1793 56217 1805 56220
rect 1936 56217 1942 56229
rect 1793 56189 1942 56217
rect 1793 56186 1805 56189
rect 1747 56180 1805 56186
rect 1936 56177 1942 56189
rect 1994 56177 2000 56229
rect 2512 56217 2518 56229
rect 2473 56189 2518 56217
rect 2512 56177 2518 56189
rect 2570 56177 2576 56229
rect 2896 56217 2902 56229
rect 2857 56189 2902 56217
rect 2896 56177 2902 56189
rect 2954 56217 2960 56229
rect 3283 56220 3341 56226
rect 3283 56217 3295 56220
rect 2954 56189 3295 56217
rect 2954 56177 2960 56189
rect 3283 56186 3295 56189
rect 3329 56186 3341 56220
rect 3283 56180 3341 56186
rect 4243 56220 4301 56226
rect 4243 56186 4255 56220
rect 4289 56217 4301 56220
rect 4531 56220 4589 56226
rect 4531 56217 4543 56220
rect 4289 56189 4543 56217
rect 4289 56186 4301 56189
rect 4243 56180 4301 56186
rect 4531 56186 4543 56189
rect 4577 56217 4589 56220
rect 4720 56217 4726 56229
rect 4577 56189 4726 56217
rect 4577 56186 4589 56189
rect 4531 56180 4589 56186
rect 4720 56177 4726 56189
rect 4778 56177 4784 56229
rect 5200 56217 5206 56229
rect 5161 56189 5206 56217
rect 5200 56177 5206 56189
rect 5258 56217 5264 56229
rect 5587 56220 5645 56226
rect 5587 56217 5599 56220
rect 5258 56189 5599 56217
rect 5258 56177 5264 56189
rect 5587 56186 5599 56189
rect 5633 56186 5645 56220
rect 5587 56180 5645 56186
rect 6067 56220 6125 56226
rect 6067 56186 6079 56220
rect 6113 56217 6125 56220
rect 6352 56217 6358 56229
rect 6113 56189 6358 56217
rect 6113 56186 6125 56189
rect 6067 56180 6125 56186
rect 6352 56177 6358 56189
rect 6410 56177 6416 56229
rect 6931 56220 6989 56226
rect 6931 56186 6943 56220
rect 6977 56217 6989 56220
rect 7216 56217 7222 56229
rect 6977 56189 7222 56217
rect 6977 56186 6989 56189
rect 6931 56180 6989 56186
rect 7216 56177 7222 56189
rect 7274 56217 7280 56229
rect 7274 56189 7367 56217
rect 7274 56177 7280 56189
rect 8560 56177 8566 56229
rect 8618 56217 8624 56229
rect 10099 56220 10157 56226
rect 8618 56189 8663 56217
rect 8618 56177 8624 56189
rect 10099 56186 10111 56220
rect 10145 56217 10157 56220
rect 10387 56220 10445 56226
rect 10387 56217 10399 56220
rect 10145 56189 10399 56217
rect 10145 56186 10157 56189
rect 10099 56180 10157 56186
rect 10387 56186 10399 56189
rect 10433 56217 10445 56220
rect 10576 56217 10582 56229
rect 10433 56189 10582 56217
rect 10433 56186 10445 56189
rect 10387 56180 10445 56186
rect 10576 56177 10582 56189
rect 10634 56177 10640 56229
rect 11152 56217 11158 56229
rect 11113 56189 11158 56217
rect 11152 56177 11158 56189
rect 11210 56177 11216 56229
rect 11536 56217 11542 56229
rect 11497 56189 11542 56217
rect 11536 56177 11542 56189
rect 11594 56217 11600 56229
rect 11923 56220 11981 56226
rect 11923 56217 11935 56220
rect 11594 56189 11935 56217
rect 11594 56177 11600 56189
rect 11923 56186 11935 56189
rect 11969 56186 11981 56220
rect 12688 56217 12694 56229
rect 12649 56189 12694 56217
rect 11923 56180 11981 56186
rect 12688 56177 12694 56189
rect 12746 56177 12752 56229
rect 13552 56177 13558 56229
rect 13610 56217 13616 56229
rect 14704 56217 14710 56229
rect 13610 56189 13655 56217
rect 14665 56189 14710 56217
rect 13610 56177 13616 56189
rect 14704 56177 14710 56189
rect 14762 56217 14768 56229
rect 14995 56220 15053 56226
rect 14995 56217 15007 56220
rect 14762 56189 15007 56217
rect 14762 56177 14768 56189
rect 14995 56186 15007 56189
rect 15041 56186 15053 56220
rect 15472 56217 15478 56229
rect 15433 56189 15478 56217
rect 14995 56180 15053 56186
rect 15472 56177 15478 56189
rect 15530 56217 15536 56229
rect 15763 56220 15821 56226
rect 15763 56217 15775 56220
rect 15530 56189 15775 56217
rect 15530 56177 15536 56189
rect 15763 56186 15775 56189
rect 15809 56186 15821 56220
rect 15763 56180 15821 56186
rect 15859 56220 15917 56226
rect 15859 56186 15871 56220
rect 15905 56186 15917 56220
rect 15859 56180 15917 56186
rect 15376 56103 15382 56155
rect 15434 56143 15440 56155
rect 15874 56143 15902 56180
rect 15952 56177 15958 56229
rect 16010 56217 16016 56229
rect 16819 56220 16877 56226
rect 16819 56217 16831 56220
rect 16010 56189 16831 56217
rect 16010 56177 16016 56189
rect 16819 56186 16831 56189
rect 16865 56217 16877 56220
rect 17107 56220 17165 56226
rect 17107 56217 17119 56220
rect 16865 56189 17119 56217
rect 16865 56186 16877 56189
rect 16819 56180 16877 56186
rect 17107 56186 17119 56189
rect 17153 56186 17165 56220
rect 18256 56217 18262 56229
rect 18217 56189 18262 56217
rect 17107 56180 17165 56186
rect 18256 56177 18262 56189
rect 18314 56177 18320 56229
rect 19024 56217 19030 56229
rect 18985 56189 19030 56217
rect 19024 56177 19030 56189
rect 19082 56177 19088 56229
rect 20371 56220 20429 56226
rect 20371 56186 20383 56220
rect 20417 56217 20429 56220
rect 20560 56217 20566 56229
rect 20417 56189 20566 56217
rect 20417 56186 20429 56189
rect 20371 56180 20429 56186
rect 20560 56177 20566 56189
rect 20618 56177 20624 56229
rect 21040 56217 21046 56229
rect 21001 56189 21046 56217
rect 21040 56177 21046 56189
rect 21098 56217 21104 56229
rect 21331 56220 21389 56226
rect 21331 56217 21343 56220
rect 21098 56189 21343 56217
rect 21098 56177 21104 56189
rect 21331 56186 21343 56189
rect 21377 56186 21389 56220
rect 21331 56180 21389 56186
rect 22675 56220 22733 56226
rect 22675 56186 22687 56220
rect 22721 56217 22733 56220
rect 22864 56217 22870 56229
rect 22721 56189 22870 56217
rect 22721 56186 22733 56189
rect 22675 56180 22733 56186
rect 22864 56177 22870 56189
rect 22922 56177 22928 56229
rect 24115 56220 24173 56226
rect 24115 56186 24127 56220
rect 24161 56217 24173 56220
rect 24304 56217 24310 56229
rect 24161 56189 24310 56217
rect 24161 56186 24173 56189
rect 24115 56180 24173 56186
rect 24304 56177 24310 56189
rect 24362 56177 24368 56229
rect 26512 56217 26518 56229
rect 26473 56189 26518 56217
rect 26512 56177 26518 56189
rect 26570 56217 26576 56229
rect 26803 56220 26861 56226
rect 26803 56217 26815 56220
rect 26570 56189 26815 56217
rect 26570 56177 26576 56189
rect 26803 56186 26815 56189
rect 26849 56186 26861 56220
rect 26803 56180 26861 56186
rect 27475 56220 27533 56226
rect 27475 56186 27487 56220
rect 27521 56217 27533 56220
rect 27664 56217 27670 56229
rect 27521 56189 27670 56217
rect 27521 56186 27533 56189
rect 27475 56180 27533 56186
rect 27664 56177 27670 56189
rect 27722 56177 27728 56229
rect 28144 56217 28150 56229
rect 28105 56189 28150 56217
rect 28144 56177 28150 56189
rect 28202 56217 28208 56229
rect 28531 56220 28589 56226
rect 28531 56217 28543 56220
rect 28202 56189 28543 56217
rect 28202 56177 28208 56189
rect 28531 56186 28543 56189
rect 28577 56186 28589 56220
rect 29296 56217 29302 56229
rect 29257 56189 29302 56217
rect 28531 56180 28589 56186
rect 29296 56177 29302 56189
rect 29354 56217 29360 56229
rect 29587 56220 29645 56226
rect 29587 56217 29599 56220
rect 29354 56189 29599 56217
rect 29354 56177 29360 56189
rect 29587 56186 29599 56189
rect 29633 56186 29645 56220
rect 30928 56217 30934 56229
rect 30889 56189 30934 56217
rect 29587 56180 29645 56186
rect 30928 56177 30934 56189
rect 30986 56177 30992 56229
rect 32464 56217 32470 56229
rect 32425 56189 32470 56217
rect 32464 56177 32470 56189
rect 32522 56177 32528 56229
rect 32947 56220 33005 56226
rect 32947 56186 32959 56220
rect 32993 56217 33005 56220
rect 33040 56217 33046 56229
rect 32993 56189 33046 56217
rect 32993 56186 33005 56189
rect 32947 56180 33005 56186
rect 33040 56177 33046 56189
rect 33098 56217 33104 56229
rect 33139 56220 33197 56226
rect 33139 56217 33151 56220
rect 33098 56189 33151 56217
rect 33098 56177 33104 56189
rect 33139 56186 33151 56189
rect 33185 56186 33197 56220
rect 33139 56180 33197 56186
rect 33235 56220 33293 56226
rect 33235 56186 33247 56220
rect 33281 56186 33293 56220
rect 34384 56217 34390 56229
rect 34345 56189 34390 56217
rect 33235 56180 33293 56186
rect 15434 56115 15902 56143
rect 15434 56103 15440 56115
rect 32752 56103 32758 56155
rect 32810 56143 32816 56155
rect 33250 56143 33278 56180
rect 34384 56177 34390 56189
rect 34442 56217 34448 56229
rect 34675 56220 34733 56226
rect 34675 56217 34687 56220
rect 34442 56189 34687 56217
rect 34442 56177 34448 56189
rect 34675 56186 34687 56189
rect 34721 56186 34733 56220
rect 34675 56180 34733 56186
rect 35923 56220 35981 56226
rect 35923 56186 35935 56220
rect 35969 56217 35981 56220
rect 36208 56217 36214 56229
rect 35969 56189 36214 56217
rect 35969 56186 35981 56189
rect 35923 56180 35981 56186
rect 36208 56177 36214 56189
rect 36266 56177 36272 56229
rect 36592 56217 36598 56229
rect 36553 56189 36598 56217
rect 36592 56177 36598 56189
rect 36650 56217 36656 56229
rect 36883 56220 36941 56226
rect 36883 56217 36895 56220
rect 36650 56189 36895 56217
rect 36650 56177 36656 56189
rect 36883 56186 36895 56189
rect 36929 56186 36941 56220
rect 36883 56180 36941 56186
rect 37459 56220 37517 56226
rect 37459 56186 37471 56220
rect 37505 56217 37517 56220
rect 37648 56217 37654 56229
rect 37505 56189 37654 56217
rect 37505 56186 37517 56189
rect 37459 56180 37517 56186
rect 37648 56177 37654 56189
rect 37706 56177 37712 56229
rect 38608 56177 38614 56229
rect 38666 56217 38672 56229
rect 38803 56220 38861 56226
rect 38803 56217 38815 56220
rect 38666 56189 38815 56217
rect 38666 56177 38672 56189
rect 38803 56186 38815 56189
rect 38849 56186 38861 56220
rect 39856 56217 39862 56229
rect 39817 56189 39862 56217
rect 38803 56180 38861 56186
rect 39856 56177 39862 56189
rect 39914 56217 39920 56229
rect 40243 56220 40301 56226
rect 40243 56217 40255 56220
rect 39914 56189 40255 56217
rect 39914 56177 39920 56189
rect 40243 56186 40255 56189
rect 40289 56186 40301 56220
rect 40243 56180 40301 56186
rect 41104 56177 41110 56229
rect 41162 56217 41168 56229
rect 42451 56220 42509 56226
rect 41162 56189 42398 56217
rect 41162 56177 41168 56189
rect 32810 56115 33278 56143
rect 32810 56103 32816 56115
rect 37072 56103 37078 56155
rect 37130 56143 37136 56155
rect 40816 56143 40822 56155
rect 37130 56115 40822 56143
rect 37130 56103 37136 56115
rect 40816 56103 40822 56115
rect 40874 56103 40880 56155
rect 42370 56143 42398 56189
rect 42451 56186 42463 56220
rect 42497 56217 42509 56220
rect 42640 56217 42646 56229
rect 42497 56189 42646 56217
rect 42497 56186 42509 56189
rect 42451 56180 42509 56186
rect 42640 56177 42646 56189
rect 42698 56177 42704 56229
rect 44275 56220 44333 56226
rect 44275 56217 44287 56220
rect 42754 56189 44287 56217
rect 42754 56143 42782 56189
rect 44275 56186 44287 56189
rect 44321 56186 44333 56220
rect 44275 56180 44333 56186
rect 44368 56177 44374 56229
rect 44426 56217 44432 56229
rect 46771 56220 46829 56226
rect 46771 56217 46783 56220
rect 44426 56189 46783 56217
rect 44426 56177 44432 56189
rect 46771 56186 46783 56189
rect 46817 56186 46829 56220
rect 46771 56180 46829 56186
rect 46864 56177 46870 56229
rect 46922 56217 46928 56229
rect 48211 56220 48269 56226
rect 48211 56217 48223 56220
rect 46922 56189 48223 56217
rect 46922 56177 46928 56189
rect 48211 56186 48223 56189
rect 48257 56186 48269 56220
rect 48211 56180 48269 56186
rect 48691 56220 48749 56226
rect 48691 56186 48703 56220
rect 48737 56217 48749 56220
rect 48880 56217 48886 56229
rect 48737 56189 48886 56217
rect 48737 56186 48749 56189
rect 48691 56180 48749 56186
rect 48880 56177 48886 56189
rect 48938 56177 48944 56229
rect 48979 56220 49037 56226
rect 48979 56186 48991 56220
rect 49025 56186 49037 56220
rect 48979 56180 49037 56186
rect 49555 56220 49613 56226
rect 49555 56186 49567 56220
rect 49601 56217 49613 56220
rect 49843 56220 49901 56226
rect 49843 56217 49855 56220
rect 49601 56189 49855 56217
rect 49601 56186 49613 56189
rect 49555 56180 49613 56186
rect 49843 56186 49855 56189
rect 49889 56217 49901 56220
rect 52162 56217 52190 56263
rect 52624 56217 52630 56229
rect 49889 56189 52190 56217
rect 52585 56189 52630 56217
rect 49889 56186 49901 56189
rect 49843 56180 49901 56186
rect 42370 56115 42782 56143
rect 48592 56103 48598 56155
rect 48650 56143 48656 56155
rect 48994 56143 49022 56180
rect 52624 56177 52630 56189
rect 52682 56217 52688 56229
rect 52915 56220 52973 56226
rect 52915 56217 52927 56220
rect 52682 56189 52927 56217
rect 52682 56177 52688 56189
rect 52915 56186 52927 56189
rect 52961 56217 52973 56220
rect 53203 56220 53261 56226
rect 53203 56217 53215 56220
rect 52961 56189 53215 56217
rect 52961 56186 52973 56189
rect 52915 56180 52973 56186
rect 53203 56186 53215 56189
rect 53249 56186 53261 56220
rect 53203 56180 53261 56186
rect 53491 56220 53549 56226
rect 53491 56186 53503 56220
rect 53537 56217 53549 56220
rect 53680 56217 53686 56229
rect 53537 56189 53686 56217
rect 53537 56186 53549 56189
rect 53491 56180 53549 56186
rect 53680 56177 53686 56189
rect 53738 56177 53744 56229
rect 53794 56217 53822 56263
rect 54544 56251 54550 56263
rect 54602 56251 54608 56303
rect 55024 56251 55030 56303
rect 55082 56291 55088 56303
rect 55699 56294 55757 56300
rect 55699 56291 55711 56294
rect 55082 56263 55711 56291
rect 55082 56251 55088 56263
rect 55699 56260 55711 56263
rect 55745 56291 55757 56294
rect 55987 56294 56045 56300
rect 55987 56291 55999 56294
rect 55745 56263 55999 56291
rect 55745 56260 55757 56263
rect 55699 56254 55757 56260
rect 55987 56260 55999 56263
rect 56033 56260 56045 56294
rect 55987 56254 56045 56260
rect 57811 56294 57869 56300
rect 57811 56260 57823 56294
rect 57857 56291 57869 56294
rect 58576 56291 58582 56303
rect 57857 56263 58582 56291
rect 57857 56260 57869 56263
rect 57811 56254 57869 56260
rect 58576 56251 58582 56263
rect 58634 56251 58640 56303
rect 55312 56217 55318 56229
rect 53794 56189 55166 56217
rect 55273 56189 55318 56217
rect 48650 56115 49022 56143
rect 55138 56143 55166 56189
rect 55312 56177 55318 56189
rect 55370 56177 55376 56229
rect 56944 56217 56950 56229
rect 55426 56189 56950 56217
rect 55426 56143 55454 56189
rect 56944 56177 56950 56189
rect 57002 56177 57008 56229
rect 55138 56115 55454 56143
rect 48650 56103 48656 56115
rect 1152 55970 58848 55992
rect 1152 55918 4294 55970
rect 4346 55918 4358 55970
rect 4410 55918 4422 55970
rect 4474 55918 4486 55970
rect 4538 55918 35014 55970
rect 35066 55918 35078 55970
rect 35130 55918 35142 55970
rect 35194 55918 35206 55970
rect 35258 55918 58848 55970
rect 1152 55896 58848 55918
rect 1168 55659 1174 55711
rect 1226 55699 1232 55711
rect 1651 55702 1709 55708
rect 1651 55699 1663 55702
rect 1226 55671 1663 55699
rect 1226 55659 1232 55671
rect 1651 55668 1663 55671
rect 1697 55668 1709 55702
rect 1651 55662 1709 55668
rect 4435 55702 4493 55708
rect 4435 55668 4447 55702
rect 4481 55699 4493 55702
rect 4624 55699 4630 55711
rect 4481 55671 4630 55699
rect 4481 55668 4493 55671
rect 4435 55662 4493 55668
rect 4624 55659 4630 55671
rect 4682 55659 4688 55711
rect 7504 55659 7510 55711
rect 7562 55699 7568 55711
rect 7603 55702 7661 55708
rect 7603 55699 7615 55702
rect 7562 55671 7615 55699
rect 7562 55659 7568 55671
rect 7603 55668 7615 55671
rect 7649 55668 7661 55702
rect 7603 55662 7661 55668
rect 9136 55659 9142 55711
rect 9194 55699 9200 55711
rect 9331 55702 9389 55708
rect 9331 55699 9343 55702
rect 9194 55671 9343 55699
rect 9194 55659 9200 55671
rect 9331 55668 9343 55671
rect 9377 55668 9389 55702
rect 9331 55662 9389 55668
rect 13840 55659 13846 55711
rect 13898 55699 13904 55711
rect 13939 55702 13997 55708
rect 13939 55699 13951 55702
rect 13898 55671 13951 55699
rect 13898 55659 13904 55671
rect 13939 55668 13951 55671
rect 13985 55668 13997 55702
rect 13939 55662 13997 55668
rect 20176 55659 20182 55711
rect 20234 55699 20240 55711
rect 20275 55702 20333 55708
rect 20275 55699 20287 55702
rect 20234 55671 20287 55699
rect 20234 55659 20240 55671
rect 20275 55668 20287 55671
rect 20321 55668 20333 55702
rect 20275 55662 20333 55668
rect 23344 55659 23350 55711
rect 23402 55699 23408 55711
rect 23539 55702 23597 55708
rect 23539 55699 23551 55702
rect 23402 55671 23551 55699
rect 23402 55659 23408 55671
rect 23539 55668 23551 55671
rect 23585 55668 23597 55702
rect 23539 55662 23597 55668
rect 24880 55659 24886 55711
rect 24938 55699 24944 55711
rect 24979 55702 25037 55708
rect 24979 55699 24991 55702
rect 24938 55671 24991 55699
rect 24938 55659 24944 55671
rect 24979 55668 24991 55671
rect 25025 55668 25037 55702
rect 24979 55662 25037 55668
rect 39088 55659 39094 55711
rect 39146 55699 39152 55711
rect 39283 55702 39341 55708
rect 39283 55699 39295 55702
rect 39146 55671 39295 55699
rect 39146 55659 39152 55671
rect 39283 55668 39295 55671
rect 39329 55668 39341 55702
rect 39283 55662 39341 55668
rect 40720 55659 40726 55711
rect 40778 55699 40784 55711
rect 40915 55702 40973 55708
rect 40915 55699 40927 55702
rect 40778 55671 40927 55699
rect 40778 55659 40784 55671
rect 40915 55668 40927 55671
rect 40961 55668 40973 55702
rect 40915 55662 40973 55668
rect 45424 55659 45430 55711
rect 45482 55699 45488 55711
rect 45619 55702 45677 55708
rect 45619 55699 45631 55702
rect 45482 55671 45631 55699
rect 45482 55659 45488 55671
rect 45619 55668 45631 55671
rect 45665 55668 45677 55702
rect 45619 55662 45677 55668
rect 46960 55659 46966 55711
rect 47018 55699 47024 55711
rect 47059 55702 47117 55708
rect 47059 55699 47071 55702
rect 47018 55671 47071 55699
rect 47018 55659 47024 55671
rect 47059 55668 47071 55671
rect 47105 55668 47117 55702
rect 47059 55662 47117 55668
rect 51760 55659 51766 55711
rect 51818 55699 51824 55711
rect 51859 55702 51917 55708
rect 51859 55699 51871 55702
rect 51818 55671 51871 55699
rect 51818 55659 51824 55671
rect 51859 55668 51871 55671
rect 51905 55668 51917 55702
rect 51859 55662 51917 55668
rect 56464 55659 56470 55711
rect 56522 55699 56528 55711
rect 56659 55702 56717 55708
rect 56659 55699 56671 55702
rect 56522 55671 56671 55699
rect 56522 55659 56528 55671
rect 56659 55668 56671 55671
rect 56705 55668 56717 55702
rect 56659 55662 56717 55668
rect 57520 55659 57526 55711
rect 57578 55699 57584 55711
rect 57715 55702 57773 55708
rect 57715 55699 57727 55702
rect 57578 55671 57727 55699
rect 57578 55659 57584 55671
rect 57715 55668 57727 55671
rect 57761 55668 57773 55702
rect 57715 55662 57773 55668
rect 38800 55585 38806 55637
rect 38858 55625 38864 55637
rect 51955 55628 52013 55634
rect 51955 55625 51967 55628
rect 38858 55597 51967 55625
rect 38858 55585 38864 55597
rect 51955 55594 51967 55597
rect 52001 55594 52013 55628
rect 51955 55588 52013 55594
rect 1747 55554 1805 55560
rect 1747 55520 1759 55554
rect 1793 55551 1805 55554
rect 1840 55551 1846 55563
rect 1793 55523 1846 55551
rect 1793 55520 1805 55523
rect 1747 55514 1805 55520
rect 1840 55511 1846 55523
rect 1898 55511 1904 55563
rect 4243 55554 4301 55560
rect 4243 55520 4255 55554
rect 4289 55551 4301 55554
rect 4531 55554 4589 55560
rect 4531 55551 4543 55554
rect 4289 55523 4543 55551
rect 4289 55520 4301 55523
rect 4243 55514 4301 55520
rect 4531 55520 4543 55523
rect 4577 55551 4589 55554
rect 4624 55551 4630 55563
rect 4577 55523 4630 55551
rect 4577 55520 4589 55523
rect 4531 55514 4589 55520
rect 4624 55511 4630 55523
rect 4682 55511 4688 55563
rect 7411 55554 7469 55560
rect 7411 55520 7423 55554
rect 7457 55551 7469 55554
rect 7696 55551 7702 55563
rect 7457 55523 7702 55551
rect 7457 55520 7469 55523
rect 7411 55514 7469 55520
rect 7696 55511 7702 55523
rect 7754 55511 7760 55563
rect 9235 55554 9293 55560
rect 9235 55551 9247 55554
rect 8962 55523 9247 55551
rect 8962 55415 8990 55523
rect 9235 55520 9247 55523
rect 9281 55520 9293 55554
rect 14035 55554 14093 55560
rect 14035 55551 14047 55554
rect 9235 55514 9293 55520
rect 13666 55523 14047 55551
rect 13666 55415 13694 55523
rect 14035 55520 14047 55523
rect 14081 55520 14093 55554
rect 14035 55514 14093 55520
rect 20083 55554 20141 55560
rect 20083 55520 20095 55554
rect 20129 55551 20141 55554
rect 20368 55551 20374 55563
rect 20129 55523 20374 55551
rect 20129 55520 20141 55523
rect 20083 55514 20141 55520
rect 20368 55511 20374 55523
rect 20426 55511 20432 55563
rect 23251 55554 23309 55560
rect 23251 55520 23263 55554
rect 23297 55551 23309 55554
rect 23440 55551 23446 55563
rect 23297 55523 23446 55551
rect 23297 55520 23309 55523
rect 23251 55514 23309 55520
rect 23440 55511 23446 55523
rect 23498 55511 23504 55563
rect 24787 55554 24845 55560
rect 24787 55520 24799 55554
rect 24833 55551 24845 55554
rect 25072 55551 25078 55563
rect 24833 55523 25078 55551
rect 24833 55520 24845 55523
rect 24787 55514 24845 55520
rect 25072 55511 25078 55523
rect 25130 55511 25136 55563
rect 27955 55554 28013 55560
rect 27955 55520 27967 55554
rect 28001 55551 28013 55554
rect 28240 55551 28246 55563
rect 28001 55523 28246 55551
rect 28001 55520 28013 55523
rect 27955 55514 28013 55520
rect 28240 55511 28246 55523
rect 28298 55511 28304 55563
rect 29011 55554 29069 55560
rect 29011 55520 29023 55554
rect 29057 55520 29069 55554
rect 39187 55554 39245 55560
rect 39187 55551 39199 55554
rect 29011 55514 29069 55520
rect 38914 55523 39199 55551
rect 29026 55415 29054 55514
rect 38914 55415 38942 55523
rect 39187 55520 39199 55523
rect 39233 55520 39245 55554
rect 39187 55514 39245 55520
rect 40627 55554 40685 55560
rect 40627 55520 40639 55554
rect 40673 55551 40685 55554
rect 40816 55551 40822 55563
rect 40673 55523 40822 55551
rect 40673 55520 40685 55523
rect 40627 55514 40685 55520
rect 40816 55511 40822 55523
rect 40874 55511 40880 55563
rect 45523 55554 45581 55560
rect 45523 55551 45535 55554
rect 45250 55523 45535 55551
rect 8944 55403 8950 55415
rect 8905 55375 8950 55403
rect 8944 55363 8950 55375
rect 9002 55363 9008 55415
rect 13648 55403 13654 55415
rect 13609 55375 13654 55403
rect 13648 55363 13654 55375
rect 13706 55363 13712 55415
rect 28915 55406 28973 55412
rect 28915 55372 28927 55406
rect 28961 55403 28973 55406
rect 29008 55403 29014 55415
rect 28961 55375 29014 55403
rect 28961 55372 28973 55375
rect 28915 55366 28973 55372
rect 29008 55363 29014 55375
rect 29066 55363 29072 55415
rect 38896 55403 38902 55415
rect 38857 55375 38902 55403
rect 38896 55363 38902 55375
rect 38954 55363 38960 55415
rect 45136 55363 45142 55415
rect 45194 55403 45200 55415
rect 45250 55412 45278 55523
rect 45523 55520 45535 55523
rect 45569 55520 45581 55554
rect 47152 55551 47158 55563
rect 47113 55523 47158 55551
rect 45523 55514 45581 55520
rect 47152 55511 47158 55523
rect 47210 55511 47216 55563
rect 49171 55554 49229 55560
rect 49171 55520 49183 55554
rect 49217 55520 49229 55554
rect 49171 55514 49229 55520
rect 56371 55554 56429 55560
rect 56371 55520 56383 55554
rect 56417 55551 56429 55554
rect 56560 55551 56566 55563
rect 56417 55523 56566 55551
rect 56417 55520 56429 55523
rect 56371 55514 56429 55520
rect 49186 55415 49214 55514
rect 56560 55511 56566 55523
rect 56618 55511 56624 55563
rect 57424 55551 57430 55563
rect 57337 55523 57430 55551
rect 57424 55511 57430 55523
rect 57482 55551 57488 55563
rect 57619 55554 57677 55560
rect 57619 55551 57631 55554
rect 57482 55523 57631 55551
rect 57482 55511 57488 55523
rect 57619 55520 57631 55523
rect 57665 55520 57677 55554
rect 57619 55514 57677 55520
rect 45235 55406 45293 55412
rect 45235 55403 45247 55406
rect 45194 55375 45247 55403
rect 45194 55363 45200 55375
rect 45235 55372 45247 55375
rect 45281 55372 45293 55406
rect 45235 55366 45293 55372
rect 49075 55406 49133 55412
rect 49075 55372 49087 55406
rect 49121 55403 49133 55406
rect 49168 55403 49174 55415
rect 49121 55375 49174 55403
rect 49121 55372 49133 55375
rect 49075 55366 49133 55372
rect 49168 55363 49174 55375
rect 49226 55363 49232 55415
rect 1152 55304 58848 55326
rect 1152 55252 19654 55304
rect 19706 55252 19718 55304
rect 19770 55252 19782 55304
rect 19834 55252 19846 55304
rect 19898 55252 50374 55304
rect 50426 55252 50438 55304
rect 50490 55252 50502 55304
rect 50554 55252 50566 55304
rect 50618 55252 58848 55304
rect 1152 55230 58848 55252
rect 57907 55184 57965 55190
rect 57907 55150 57919 55184
rect 57953 55181 57965 55184
rect 59152 55181 59158 55193
rect 57953 55153 59158 55181
rect 57953 55150 57965 55153
rect 57907 55144 57965 55150
rect 59152 55141 59158 55153
rect 59210 55141 59216 55193
rect 35344 55067 35350 55119
rect 35402 55107 35408 55119
rect 47152 55107 47158 55119
rect 35402 55079 47158 55107
rect 35402 55067 35408 55079
rect 47152 55067 47158 55079
rect 47210 55067 47216 55119
rect 28240 54993 28246 55045
rect 28298 55033 28304 55045
rect 55600 55033 55606 55045
rect 28298 55005 55606 55033
rect 28298 54993 28304 55005
rect 55600 54993 55606 55005
rect 55658 54993 55664 55045
rect 27571 54888 27629 54894
rect 27571 54885 27583 54888
rect 27394 54857 27583 54885
rect 27283 54814 27341 54820
rect 27283 54780 27295 54814
rect 27329 54811 27341 54814
rect 27394 54811 27422 54857
rect 27571 54854 27583 54857
rect 27617 54885 27629 54888
rect 57619 54888 57677 54894
rect 27617 54857 37454 54885
rect 27617 54854 27629 54857
rect 27571 54848 27629 54854
rect 37426 54811 37454 54857
rect 57619 54854 57631 54888
rect 57665 54885 57677 54888
rect 57811 54888 57869 54894
rect 57811 54885 57823 54888
rect 57665 54857 57823 54885
rect 57665 54854 57677 54857
rect 57619 54848 57677 54854
rect 57811 54854 57823 54857
rect 57857 54854 57869 54888
rect 57811 54848 57869 54854
rect 50224 54811 50230 54823
rect 27329 54783 27422 54811
rect 27490 54783 27710 54811
rect 37426 54783 50230 54811
rect 27329 54780 27341 54783
rect 27283 54774 27341 54780
rect 25264 54737 25270 54749
rect 25225 54709 25270 54737
rect 25264 54697 25270 54709
rect 25322 54737 25328 54749
rect 25651 54740 25709 54746
rect 25651 54737 25663 54740
rect 25322 54709 25663 54737
rect 25322 54697 25328 54709
rect 25651 54706 25663 54709
rect 25697 54706 25709 54740
rect 25651 54700 25709 54706
rect 26611 54740 26669 54746
rect 26611 54706 26623 54740
rect 26657 54737 26669 54740
rect 26899 54740 26957 54746
rect 26899 54737 26911 54740
rect 26657 54709 26911 54737
rect 26657 54706 26669 54709
rect 26611 54700 26669 54706
rect 26899 54706 26911 54709
rect 26945 54737 26957 54740
rect 27490 54737 27518 54783
rect 26945 54709 27518 54737
rect 27682 54737 27710 54783
rect 50224 54771 50230 54783
rect 50282 54771 50288 54823
rect 57634 54737 57662 54848
rect 27682 54709 57662 54737
rect 26945 54706 26957 54709
rect 26899 54700 26957 54706
rect 1152 54638 58848 54660
rect 1152 54586 4294 54638
rect 4346 54586 4358 54638
rect 4410 54586 4422 54638
rect 4474 54586 4486 54638
rect 4538 54586 35014 54638
rect 35066 54586 35078 54638
rect 35130 54586 35142 54638
rect 35194 54586 35206 54638
rect 35258 54586 58848 54638
rect 1152 54564 58848 54586
rect 57907 54370 57965 54376
rect 57907 54336 57919 54370
rect 57953 54367 57965 54370
rect 58096 54367 58102 54379
rect 57953 54339 58102 54367
rect 57953 54336 57965 54339
rect 57907 54330 57965 54336
rect 58096 54327 58102 54339
rect 58154 54327 58160 54379
rect 56563 54222 56621 54228
rect 56563 54188 56575 54222
rect 56609 54188 56621 54222
rect 56563 54182 56621 54188
rect 57619 54222 57677 54228
rect 57619 54188 57631 54222
rect 57665 54219 57677 54222
rect 57808 54219 57814 54231
rect 57665 54191 57814 54219
rect 57665 54188 57677 54191
rect 57619 54182 57677 54188
rect 56368 54071 56374 54083
rect 56329 54043 56374 54071
rect 56368 54031 56374 54043
rect 56426 54071 56432 54083
rect 56578 54071 56606 54182
rect 57808 54179 57814 54191
rect 57866 54219 57872 54231
rect 58099 54222 58157 54228
rect 58099 54219 58111 54222
rect 57866 54191 58111 54219
rect 57866 54179 57872 54191
rect 58099 54188 58111 54191
rect 58145 54188 58157 54222
rect 58099 54182 58157 54188
rect 56426 54043 56606 54071
rect 56426 54031 56432 54043
rect 1152 53972 58848 53994
rect 1152 53920 19654 53972
rect 19706 53920 19718 53972
rect 19770 53920 19782 53972
rect 19834 53920 19846 53972
rect 19898 53920 50374 53972
rect 50426 53920 50438 53972
rect 50490 53920 50502 53972
rect 50554 53920 50566 53972
rect 50618 53920 58848 53972
rect 1152 53898 58848 53920
rect 57907 53852 57965 53858
rect 57907 53818 57919 53852
rect 57953 53849 57965 53852
rect 59632 53849 59638 53861
rect 57953 53821 59638 53849
rect 57953 53818 57965 53821
rect 57907 53812 57965 53818
rect 59632 53809 59638 53821
rect 59690 53809 59696 53861
rect 3664 53513 3670 53565
rect 3722 53553 3728 53565
rect 55795 53556 55853 53562
rect 55795 53553 55807 53556
rect 3722 53525 55807 53553
rect 3722 53513 3728 53525
rect 55795 53522 55807 53525
rect 55841 53553 55853 53556
rect 55987 53556 56045 53562
rect 55987 53553 55999 53556
rect 55841 53525 55999 53553
rect 55841 53522 55853 53525
rect 55795 53516 55853 53522
rect 55987 53522 55999 53525
rect 56033 53522 56045 53556
rect 55987 53516 56045 53522
rect 57811 53556 57869 53562
rect 57811 53522 57823 53556
rect 57857 53522 57869 53556
rect 57811 53516 57869 53522
rect 32179 53482 32237 53488
rect 32179 53448 32191 53482
rect 32225 53479 32237 53482
rect 32467 53482 32525 53488
rect 32467 53479 32479 53482
rect 32225 53451 32479 53479
rect 32225 53448 32237 53451
rect 32179 53442 32237 53448
rect 32467 53448 32479 53451
rect 32513 53479 32525 53482
rect 44464 53479 44470 53491
rect 32513 53451 44470 53479
rect 32513 53448 32525 53451
rect 32467 53442 32525 53448
rect 44464 53439 44470 53451
rect 44522 53439 44528 53491
rect 2224 53405 2230 53417
rect 2185 53377 2230 53405
rect 2224 53365 2230 53377
rect 2282 53405 2288 53417
rect 2611 53408 2669 53414
rect 2611 53405 2623 53408
rect 2282 53377 2623 53405
rect 2282 53365 2288 53377
rect 2611 53374 2623 53377
rect 2657 53374 2669 53408
rect 17584 53405 17590 53417
rect 17545 53377 17590 53405
rect 2611 53368 2669 53374
rect 17584 53365 17590 53377
rect 17642 53405 17648 53417
rect 17971 53408 18029 53414
rect 17971 53405 17983 53408
rect 17642 53377 17983 53405
rect 17642 53365 17648 53377
rect 17971 53374 17983 53377
rect 18017 53374 18029 53408
rect 39376 53405 39382 53417
rect 39337 53377 39382 53405
rect 17971 53368 18029 53374
rect 39376 53365 39382 53377
rect 39434 53405 39440 53417
rect 39571 53408 39629 53414
rect 39571 53405 39583 53408
rect 39434 53377 39583 53405
rect 39434 53365 39440 53377
rect 39571 53374 39583 53377
rect 39617 53374 39629 53408
rect 39571 53368 39629 53374
rect 43027 53408 43085 53414
rect 43027 53374 43039 53408
rect 43073 53405 43085 53408
rect 43120 53405 43126 53417
rect 43073 53377 43126 53405
rect 43073 53374 43085 53377
rect 43027 53368 43085 53374
rect 43120 53365 43126 53377
rect 43178 53365 43184 53417
rect 57619 53408 57677 53414
rect 57619 53374 57631 53408
rect 57665 53405 57677 53408
rect 57712 53405 57718 53417
rect 57665 53377 57718 53405
rect 57665 53374 57677 53377
rect 57619 53368 57677 53374
rect 57712 53365 57718 53377
rect 57770 53405 57776 53417
rect 57826 53405 57854 53516
rect 57770 53377 57854 53405
rect 57770 53365 57776 53377
rect 1152 53306 58848 53328
rect 1152 53254 4294 53306
rect 4346 53254 4358 53306
rect 4410 53254 4422 53306
rect 4474 53254 4486 53306
rect 4538 53254 35014 53306
rect 35066 53254 35078 53306
rect 35130 53254 35142 53306
rect 35194 53254 35206 53306
rect 35258 53254 58848 53306
rect 1152 53232 58848 53254
rect 15568 52995 15574 53047
rect 15626 53035 15632 53047
rect 17683 53038 17741 53044
rect 17683 53035 17695 53038
rect 15626 53007 17695 53035
rect 15626 52995 15632 53007
rect 17683 53004 17695 53007
rect 17729 53004 17741 53038
rect 17683 52998 17741 53004
rect 6931 52890 6989 52896
rect 6931 52856 6943 52890
rect 6977 52887 6989 52890
rect 7219 52890 7277 52896
rect 7219 52887 7231 52890
rect 6977 52859 7231 52887
rect 6977 52856 6989 52859
rect 6931 52850 6989 52856
rect 7219 52856 7231 52859
rect 7265 52887 7277 52890
rect 51664 52887 51670 52899
rect 7265 52859 51670 52887
rect 7265 52856 7277 52859
rect 7219 52850 7277 52856
rect 51664 52847 51670 52859
rect 51722 52847 51728 52899
rect 1152 52640 58848 52662
rect 1152 52588 19654 52640
rect 19706 52588 19718 52640
rect 19770 52588 19782 52640
rect 19834 52588 19846 52640
rect 19898 52588 50374 52640
rect 50426 52588 50438 52640
rect 50490 52588 50502 52640
rect 50554 52588 50566 52640
rect 50618 52588 58848 52640
rect 1152 52566 58848 52588
rect 37747 52372 37805 52378
rect 37747 52338 37759 52372
rect 37793 52369 37805 52372
rect 38128 52369 38134 52381
rect 37793 52341 38134 52369
rect 37793 52338 37805 52341
rect 37747 52332 37805 52338
rect 38128 52329 38134 52341
rect 38186 52329 38192 52381
rect 31312 52147 31318 52159
rect 7186 52119 31318 52147
rect 3091 52076 3149 52082
rect 3091 52042 3103 52076
rect 3137 52073 3149 52076
rect 3379 52076 3437 52082
rect 3379 52073 3391 52076
rect 3137 52045 3391 52073
rect 3137 52042 3149 52045
rect 3091 52036 3149 52042
rect 3379 52042 3391 52045
rect 3425 52073 3437 52076
rect 7186 52073 7214 52119
rect 31312 52107 31318 52119
rect 31370 52107 31376 52159
rect 3425 52045 7214 52073
rect 18067 52076 18125 52082
rect 3425 52042 3437 52045
rect 3379 52036 3437 52042
rect 18067 52042 18079 52076
rect 18113 52073 18125 52076
rect 18352 52073 18358 52085
rect 18113 52045 18358 52073
rect 18113 52042 18125 52045
rect 18067 52036 18125 52042
rect 18352 52033 18358 52045
rect 18410 52033 18416 52085
rect 39763 52076 39821 52082
rect 39763 52042 39775 52076
rect 39809 52073 39821 52076
rect 40048 52073 40054 52085
rect 39809 52045 40054 52073
rect 39809 52042 39821 52045
rect 39763 52036 39821 52042
rect 40048 52033 40054 52045
rect 40106 52033 40112 52085
rect 1152 51974 58848 51996
rect 1152 51922 4294 51974
rect 4346 51922 4358 51974
rect 4410 51922 4422 51974
rect 4474 51922 4486 51974
rect 4538 51922 35014 51974
rect 35066 51922 35078 51974
rect 35130 51922 35142 51974
rect 35194 51922 35206 51974
rect 35258 51922 58848 51974
rect 1152 51900 58848 51922
rect 29491 51706 29549 51712
rect 29491 51672 29503 51706
rect 29537 51703 29549 51706
rect 30256 51703 30262 51715
rect 29537 51675 30262 51703
rect 29537 51672 29549 51675
rect 29491 51666 29549 51672
rect 30256 51663 30262 51675
rect 30314 51663 30320 51715
rect 10291 51484 10349 51490
rect 10291 51450 10303 51484
rect 10337 51481 10349 51484
rect 44080 51481 44086 51493
rect 10337 51453 44086 51481
rect 10337 51450 10349 51453
rect 10291 51444 10349 51450
rect 44080 51441 44086 51453
rect 44138 51441 44144 51493
rect 1152 51308 58848 51330
rect 1152 51256 19654 51308
rect 19706 51256 19718 51308
rect 19770 51256 19782 51308
rect 19834 51256 19846 51308
rect 19898 51256 50374 51308
rect 50426 51256 50438 51308
rect 50490 51256 50502 51308
rect 50554 51256 50566 51308
rect 50618 51256 58848 51308
rect 1152 51234 58848 51256
rect 15763 50744 15821 50750
rect 15763 50710 15775 50744
rect 15809 50741 15821 50744
rect 16051 50744 16109 50750
rect 16051 50741 16063 50744
rect 15809 50713 16063 50741
rect 15809 50710 15821 50713
rect 15763 50704 15821 50710
rect 16051 50710 16063 50713
rect 16097 50741 16109 50744
rect 45232 50741 45238 50753
rect 16097 50713 45238 50741
rect 16097 50710 16109 50713
rect 16051 50704 16109 50710
rect 45232 50701 45238 50713
rect 45290 50701 45296 50753
rect 53584 50741 53590 50753
rect 53545 50713 53590 50741
rect 53584 50701 53590 50713
rect 53642 50741 53648 50753
rect 53779 50744 53837 50750
rect 53779 50741 53791 50744
rect 53642 50713 53791 50741
rect 53642 50701 53648 50713
rect 53779 50710 53791 50713
rect 53825 50710 53837 50744
rect 53779 50704 53837 50710
rect 1152 50642 58848 50664
rect 1152 50590 4294 50642
rect 4346 50590 4358 50642
rect 4410 50590 4422 50642
rect 4474 50590 4486 50642
rect 4538 50590 35014 50642
rect 35066 50590 35078 50642
rect 35130 50590 35142 50642
rect 35194 50590 35206 50642
rect 35258 50590 58848 50642
rect 1152 50568 58848 50590
rect 39472 50223 39478 50235
rect 39433 50195 39478 50223
rect 39472 50183 39478 50195
rect 39530 50183 39536 50235
rect 57619 50226 57677 50232
rect 57619 50192 57631 50226
rect 57665 50192 57677 50226
rect 57619 50186 57677 50192
rect 51571 50152 51629 50158
rect 51571 50149 51583 50152
rect 27346 50121 51583 50149
rect 18256 50035 18262 50087
rect 18314 50075 18320 50087
rect 27346 50075 27374 50121
rect 51571 50118 51583 50121
rect 51617 50118 51629 50152
rect 51571 50112 51629 50118
rect 57634 50087 57662 50186
rect 18314 50047 27374 50075
rect 39379 50078 39437 50084
rect 18314 50035 18320 50047
rect 39379 50044 39391 50078
rect 39425 50075 39437 50078
rect 39472 50075 39478 50087
rect 39425 50047 39478 50075
rect 39425 50044 39437 50047
rect 39379 50038 39437 50044
rect 39472 50035 39478 50047
rect 39530 50035 39536 50087
rect 57523 50078 57581 50084
rect 57523 50044 57535 50078
rect 57569 50075 57581 50078
rect 57616 50075 57622 50087
rect 57569 50047 57622 50075
rect 57569 50044 57581 50047
rect 57523 50038 57581 50044
rect 57616 50035 57622 50047
rect 57674 50075 57680 50087
rect 57674 50047 57767 50075
rect 57674 50035 57680 50047
rect 1152 49976 58848 49998
rect 1152 49924 19654 49976
rect 19706 49924 19718 49976
rect 19770 49924 19782 49976
rect 19834 49924 19846 49976
rect 19898 49924 50374 49976
rect 50426 49924 50438 49976
rect 50490 49924 50502 49976
rect 50554 49924 50566 49976
rect 50618 49924 58848 49976
rect 1152 49902 58848 49924
rect 28816 49813 28822 49865
rect 28874 49853 28880 49865
rect 57616 49853 57622 49865
rect 28874 49825 57622 49853
rect 28874 49813 28880 49825
rect 57616 49813 57622 49825
rect 57674 49813 57680 49865
rect 11827 49412 11885 49418
rect 11827 49378 11839 49412
rect 11873 49409 11885 49412
rect 11920 49409 11926 49421
rect 11873 49381 11926 49409
rect 11873 49378 11885 49381
rect 11827 49372 11885 49378
rect 11920 49369 11926 49381
rect 11978 49369 11984 49421
rect 15571 49412 15629 49418
rect 15571 49378 15583 49412
rect 15617 49409 15629 49412
rect 15664 49409 15670 49421
rect 15617 49381 15670 49409
rect 15617 49378 15629 49381
rect 15571 49372 15629 49378
rect 15664 49369 15670 49381
rect 15722 49369 15728 49421
rect 52432 49409 52438 49421
rect 52393 49381 52438 49409
rect 52432 49369 52438 49381
rect 52490 49369 52496 49421
rect 1152 49310 58848 49332
rect 1152 49258 4294 49310
rect 4346 49258 4358 49310
rect 4410 49258 4422 49310
rect 4474 49258 4486 49310
rect 4538 49258 35014 49310
rect 35066 49258 35078 49310
rect 35130 49258 35142 49310
rect 35194 49258 35206 49310
rect 35258 49258 58848 49310
rect 1152 49236 58848 49258
rect 18547 49042 18605 49048
rect 18547 49008 18559 49042
rect 18593 49039 18605 49042
rect 32656 49039 32662 49051
rect 18593 49011 32662 49039
rect 18593 49008 18605 49011
rect 18547 49002 18605 49008
rect 32656 48999 32662 49011
rect 32714 48999 32720 49051
rect 32080 48965 32086 48977
rect 7186 48937 32086 48965
rect 3283 48894 3341 48900
rect 3283 48860 3295 48894
rect 3329 48891 3341 48894
rect 3571 48894 3629 48900
rect 3571 48891 3583 48894
rect 3329 48863 3583 48891
rect 3329 48860 3341 48863
rect 3283 48854 3341 48860
rect 3571 48860 3583 48863
rect 3617 48891 3629 48894
rect 7186 48891 7214 48937
rect 32080 48925 32086 48937
rect 32138 48925 32144 48977
rect 3617 48863 7214 48891
rect 49075 48894 49133 48900
rect 3617 48860 3629 48863
rect 3571 48854 3629 48860
rect 49075 48860 49087 48894
rect 49121 48891 49133 48894
rect 49363 48894 49421 48900
rect 49363 48891 49375 48894
rect 49121 48863 49375 48891
rect 49121 48860 49133 48863
rect 49075 48854 49133 48860
rect 49363 48860 49375 48863
rect 49409 48891 49421 48894
rect 51760 48891 51766 48903
rect 49409 48863 51766 48891
rect 49409 48860 49421 48863
rect 49363 48854 49421 48860
rect 51760 48851 51766 48863
rect 51818 48851 51824 48903
rect 22771 48746 22829 48752
rect 22771 48712 22783 48746
rect 22817 48743 22829 48746
rect 44368 48743 44374 48755
rect 22817 48715 44374 48743
rect 22817 48712 22829 48715
rect 22771 48706 22829 48712
rect 44368 48703 44374 48715
rect 44426 48703 44432 48755
rect 1152 48644 58848 48666
rect 1152 48592 19654 48644
rect 19706 48592 19718 48644
rect 19770 48592 19782 48644
rect 19834 48592 19846 48644
rect 19898 48592 50374 48644
rect 50426 48592 50438 48644
rect 50490 48592 50502 48644
rect 50554 48592 50566 48644
rect 50618 48592 58848 48644
rect 1152 48570 58848 48592
rect 41296 48521 41302 48533
rect 41257 48493 41302 48521
rect 41296 48481 41302 48493
rect 41354 48481 41360 48533
rect 3760 48037 3766 48089
rect 3818 48077 3824 48089
rect 4339 48080 4397 48086
rect 4339 48077 4351 48080
rect 3818 48049 4351 48077
rect 3818 48037 3824 48049
rect 4339 48046 4351 48049
rect 4385 48077 4397 48080
rect 4435 48080 4493 48086
rect 4435 48077 4447 48080
rect 4385 48049 4447 48077
rect 4385 48046 4397 48049
rect 4339 48040 4397 48046
rect 4435 48046 4447 48049
rect 4481 48046 4493 48080
rect 4435 48040 4493 48046
rect 52240 48037 52246 48089
rect 52298 48077 52304 48089
rect 52627 48080 52685 48086
rect 52627 48077 52639 48080
rect 52298 48049 52639 48077
rect 52298 48037 52304 48049
rect 52627 48046 52639 48049
rect 52673 48077 52685 48080
rect 52819 48080 52877 48086
rect 52819 48077 52831 48080
rect 52673 48049 52831 48077
rect 52673 48046 52685 48049
rect 52627 48040 52685 48046
rect 52819 48046 52831 48049
rect 52865 48046 52877 48080
rect 52819 48040 52877 48046
rect 1152 47978 58848 48000
rect 1152 47926 4294 47978
rect 4346 47926 4358 47978
rect 4410 47926 4422 47978
rect 4474 47926 4486 47978
rect 4538 47926 35014 47978
rect 35066 47926 35078 47978
rect 35130 47926 35142 47978
rect 35194 47926 35206 47978
rect 35258 47926 58848 47978
rect 1152 47904 58848 47926
rect 34576 47559 34582 47571
rect 34489 47531 34582 47559
rect 34576 47519 34582 47531
rect 34634 47559 34640 47571
rect 34675 47562 34733 47568
rect 34675 47559 34687 47562
rect 34634 47531 34687 47559
rect 34634 47519 34640 47531
rect 34675 47528 34687 47531
rect 34721 47528 34733 47562
rect 34675 47522 34733 47528
rect 1152 47312 58848 47334
rect 1152 47260 19654 47312
rect 19706 47260 19718 47312
rect 19770 47260 19782 47312
rect 19834 47260 19846 47312
rect 19898 47260 50374 47312
rect 50426 47260 50438 47312
rect 50490 47260 50502 47312
rect 50554 47260 50566 47312
rect 50618 47260 58848 47312
rect 1152 47238 58848 47260
rect 6736 47041 6742 47053
rect 6697 47013 6742 47041
rect 6736 47001 6742 47013
rect 6794 47001 6800 47053
rect 23632 46745 23638 46757
rect 23593 46717 23638 46745
rect 23632 46705 23638 46717
rect 23690 46745 23696 46757
rect 23923 46748 23981 46754
rect 23923 46745 23935 46748
rect 23690 46717 23935 46745
rect 23690 46705 23696 46717
rect 23923 46714 23935 46717
rect 23969 46714 23981 46748
rect 23923 46708 23981 46714
rect 1152 46646 58848 46668
rect 1152 46594 4294 46646
rect 4346 46594 4358 46646
rect 4410 46594 4422 46646
rect 4474 46594 4486 46646
rect 4538 46594 35014 46646
rect 35066 46594 35078 46646
rect 35130 46594 35142 46646
rect 35194 46594 35206 46646
rect 35258 46594 58848 46646
rect 1152 46572 58848 46594
rect 9619 46230 9677 46236
rect 9619 46196 9631 46230
rect 9665 46227 9677 46230
rect 9904 46227 9910 46239
rect 9665 46199 9910 46227
rect 9665 46196 9677 46199
rect 9619 46190 9677 46196
rect 9904 46187 9910 46199
rect 9962 46187 9968 46239
rect 9442 46125 9662 46153
rect 2512 46039 2518 46091
rect 2570 46079 2576 46091
rect 9442 46079 9470 46125
rect 2570 46051 9470 46079
rect 9634 46079 9662 46125
rect 12595 46082 12653 46088
rect 12595 46079 12607 46082
rect 9634 46051 12607 46079
rect 2570 46039 2576 46051
rect 12595 46048 12607 46051
rect 12641 46048 12653 46082
rect 12595 46042 12653 46048
rect 1152 45980 58848 46002
rect 1152 45928 19654 45980
rect 19706 45928 19718 45980
rect 19770 45928 19782 45980
rect 19834 45928 19846 45980
rect 19898 45928 50374 45980
rect 50426 45928 50438 45980
rect 50490 45928 50502 45980
rect 50554 45928 50566 45980
rect 50618 45928 58848 45980
rect 1152 45906 58848 45928
rect 35059 45712 35117 45718
rect 35059 45678 35071 45712
rect 35105 45709 35117 45712
rect 35344 45709 35350 45721
rect 35105 45681 35350 45709
rect 35105 45678 35117 45681
rect 35059 45672 35117 45678
rect 35344 45669 35350 45681
rect 35402 45669 35408 45721
rect 51568 45373 51574 45425
rect 51626 45413 51632 45425
rect 51667 45416 51725 45422
rect 51667 45413 51679 45416
rect 51626 45385 51679 45413
rect 51626 45373 51632 45385
rect 51667 45382 51679 45385
rect 51713 45413 51725 45416
rect 51859 45416 51917 45422
rect 51859 45413 51871 45416
rect 51713 45385 51871 45413
rect 51713 45382 51725 45385
rect 51667 45376 51725 45382
rect 51859 45382 51871 45385
rect 51905 45382 51917 45416
rect 51859 45376 51917 45382
rect 1152 45314 58848 45336
rect 1152 45262 4294 45314
rect 4346 45262 4358 45314
rect 4410 45262 4422 45314
rect 4474 45262 4486 45314
rect 4538 45262 35014 45314
rect 35066 45262 35078 45314
rect 35130 45262 35142 45314
rect 35194 45262 35206 45314
rect 35258 45262 58848 45314
rect 1152 45240 58848 45262
rect 19984 45151 19990 45203
rect 20042 45191 20048 45203
rect 38800 45191 38806 45203
rect 20042 45163 27374 45191
rect 38761 45163 38806 45191
rect 20042 45151 20048 45163
rect 27346 45117 27374 45163
rect 38800 45151 38806 45163
rect 38858 45151 38864 45203
rect 51568 45117 51574 45129
rect 27346 45089 51574 45117
rect 51568 45077 51574 45089
rect 51626 45077 51632 45129
rect 39667 45046 39725 45052
rect 39667 45012 39679 45046
rect 39713 45043 39725 45046
rect 42448 45043 42454 45055
rect 39713 45015 42454 45043
rect 39713 45012 39725 45015
rect 39667 45006 39725 45012
rect 42448 45003 42454 45015
rect 42506 45003 42512 45055
rect 11152 44929 11158 44981
rect 11210 44969 11216 44981
rect 53491 44972 53549 44978
rect 53491 44969 53503 44972
rect 11210 44941 53503 44969
rect 11210 44929 11216 44941
rect 53491 44938 53503 44941
rect 53537 44938 53549 44972
rect 53491 44932 53549 44938
rect 8179 44898 8237 44904
rect 8179 44864 8191 44898
rect 8225 44895 8237 44898
rect 8464 44895 8470 44907
rect 8225 44867 8470 44895
rect 8225 44864 8237 44867
rect 8179 44858 8237 44864
rect 8464 44855 8470 44867
rect 8522 44855 8528 44907
rect 21043 44898 21101 44904
rect 21043 44864 21055 44898
rect 21089 44895 21101 44898
rect 21328 44895 21334 44907
rect 21089 44867 21334 44895
rect 21089 44864 21101 44867
rect 21043 44858 21101 44864
rect 21328 44855 21334 44867
rect 21386 44855 21392 44907
rect 41203 44898 41261 44904
rect 41203 44864 41215 44898
rect 41249 44864 41261 44898
rect 41203 44858 41261 44864
rect 7603 44824 7661 44830
rect 7603 44790 7615 44824
rect 7649 44821 7661 44824
rect 7649 44793 27374 44821
rect 7649 44790 7661 44793
rect 7603 44784 7661 44790
rect 27346 44747 27374 44793
rect 39667 44750 39725 44756
rect 39667 44747 39679 44750
rect 27346 44719 39679 44747
rect 39667 44716 39679 44719
rect 39713 44716 39725 44750
rect 41008 44747 41014 44759
rect 40969 44719 41014 44747
rect 39667 44710 39725 44716
rect 41008 44707 41014 44719
rect 41066 44747 41072 44759
rect 41218 44747 41246 44858
rect 41066 44719 41246 44747
rect 41066 44707 41072 44719
rect 1152 44648 58848 44670
rect 1152 44596 19654 44648
rect 19706 44596 19718 44648
rect 19770 44596 19782 44648
rect 19834 44596 19846 44648
rect 19898 44596 50374 44648
rect 50426 44596 50438 44648
rect 50490 44596 50502 44648
rect 50554 44596 50566 44648
rect 50618 44596 58848 44648
rect 1152 44574 58848 44596
rect 11059 44084 11117 44090
rect 11059 44050 11071 44084
rect 11105 44081 11117 44084
rect 11347 44084 11405 44090
rect 11347 44081 11359 44084
rect 11105 44053 11359 44081
rect 11105 44050 11117 44053
rect 11059 44044 11117 44050
rect 11347 44050 11359 44053
rect 11393 44081 11405 44084
rect 44368 44081 44374 44093
rect 11393 44053 44374 44081
rect 11393 44050 11405 44053
rect 11347 44044 11405 44050
rect 44368 44041 44374 44053
rect 44426 44041 44432 44093
rect 1152 43982 58848 44004
rect 1152 43930 4294 43982
rect 4346 43930 4358 43982
rect 4410 43930 4422 43982
rect 4474 43930 4486 43982
rect 4538 43930 35014 43982
rect 35066 43930 35078 43982
rect 35130 43930 35142 43982
rect 35194 43930 35206 43982
rect 35258 43930 58848 43982
rect 1152 43908 58848 43930
rect 12403 43566 12461 43572
rect 12403 43532 12415 43566
rect 12449 43563 12461 43566
rect 12691 43566 12749 43572
rect 12691 43563 12703 43566
rect 12449 43535 12703 43563
rect 12449 43532 12461 43535
rect 12403 43526 12461 43532
rect 12691 43532 12703 43535
rect 12737 43563 12749 43566
rect 15760 43563 15766 43575
rect 12737 43535 15766 43563
rect 12737 43532 12749 43535
rect 12691 43526 12749 43532
rect 15760 43523 15766 43535
rect 15818 43523 15824 43575
rect 50035 43566 50093 43572
rect 50035 43532 50047 43566
rect 50081 43532 50093 43566
rect 50035 43526 50093 43532
rect 50050 43427 50078 43526
rect 49939 43418 49997 43424
rect 49939 43384 49951 43418
rect 49985 43415 49997 43418
rect 50032 43415 50038 43427
rect 49985 43387 50038 43415
rect 49985 43384 49997 43387
rect 49939 43378 49997 43384
rect 50032 43375 50038 43387
rect 50090 43375 50096 43427
rect 1152 43316 58848 43338
rect 1152 43264 19654 43316
rect 19706 43264 19718 43316
rect 19770 43264 19782 43316
rect 19834 43264 19846 43316
rect 19898 43264 50374 43316
rect 50426 43264 50438 43316
rect 50490 43264 50502 43316
rect 50554 43264 50566 43316
rect 50618 43264 58848 43316
rect 1152 43242 58848 43264
rect 6547 42752 6605 42758
rect 6547 42718 6559 42752
rect 6593 42749 6605 42752
rect 40816 42749 40822 42761
rect 6593 42721 40822 42749
rect 6593 42718 6605 42721
rect 6547 42712 6605 42718
rect 40816 42709 40822 42721
rect 40874 42709 40880 42761
rect 46384 42749 46390 42761
rect 46345 42721 46390 42749
rect 46384 42709 46390 42721
rect 46442 42749 46448 42761
rect 46771 42752 46829 42758
rect 46771 42749 46783 42752
rect 46442 42721 46783 42749
rect 46442 42709 46448 42721
rect 46771 42718 46783 42721
rect 46817 42718 46829 42752
rect 46771 42712 46829 42718
rect 53872 42709 53878 42761
rect 53930 42749 53936 42761
rect 53971 42752 54029 42758
rect 53971 42749 53983 42752
rect 53930 42721 53983 42749
rect 53930 42709 53936 42721
rect 53971 42718 53983 42721
rect 54017 42749 54029 42752
rect 54163 42752 54221 42758
rect 54163 42749 54175 42752
rect 54017 42721 54175 42749
rect 54017 42718 54029 42721
rect 53971 42712 54029 42718
rect 54163 42718 54175 42721
rect 54209 42718 54221 42752
rect 54163 42712 54221 42718
rect 1152 42650 58848 42672
rect 1152 42598 4294 42650
rect 4346 42598 4358 42650
rect 4410 42598 4422 42650
rect 4474 42598 4486 42650
rect 4538 42598 35014 42650
rect 35066 42598 35078 42650
rect 35130 42598 35142 42650
rect 35194 42598 35206 42650
rect 35258 42598 58848 42650
rect 1152 42576 58848 42598
rect 32656 42487 32662 42539
rect 32714 42527 32720 42539
rect 53872 42527 53878 42539
rect 32714 42499 53878 42527
rect 32714 42487 32720 42499
rect 53872 42487 53878 42499
rect 53930 42487 53936 42539
rect 7699 42234 7757 42240
rect 7699 42200 7711 42234
rect 7745 42231 7757 42234
rect 7987 42234 8045 42240
rect 7987 42231 7999 42234
rect 7745 42203 7999 42231
rect 7745 42200 7757 42203
rect 7699 42194 7757 42200
rect 7987 42200 7999 42203
rect 8033 42231 8045 42234
rect 8033 42203 17294 42231
rect 8033 42200 8045 42203
rect 7987 42194 8045 42200
rect 17266 42083 17294 42203
rect 57328 42083 57334 42095
rect 17266 42055 57334 42083
rect 57328 42043 57334 42055
rect 57386 42043 57392 42095
rect 1152 41984 58848 42006
rect 1152 41932 19654 41984
rect 19706 41932 19718 41984
rect 19770 41932 19782 41984
rect 19834 41932 19846 41984
rect 19898 41932 50374 41984
rect 50426 41932 50438 41984
rect 50490 41932 50502 41984
rect 50554 41932 50566 41984
rect 50618 41932 58848 41984
rect 1152 41910 58848 41932
rect 4723 41790 4781 41796
rect 4723 41756 4735 41790
rect 4769 41787 4781 41790
rect 43984 41787 43990 41799
rect 4769 41759 43990 41787
rect 4769 41756 4781 41759
rect 4723 41750 4781 41756
rect 43984 41747 43990 41759
rect 44042 41747 44048 41799
rect 27283 41420 27341 41426
rect 27283 41386 27295 41420
rect 27329 41417 27341 41420
rect 27571 41420 27629 41426
rect 27571 41417 27583 41420
rect 27329 41389 27583 41417
rect 27329 41386 27341 41389
rect 27283 41380 27341 41386
rect 27571 41386 27583 41389
rect 27617 41417 27629 41420
rect 52336 41417 52342 41429
rect 27617 41389 52342 41417
rect 27617 41386 27629 41389
rect 27571 41380 27629 41386
rect 52336 41377 52342 41389
rect 52394 41377 52400 41429
rect 1152 41318 58848 41340
rect 1152 41266 4294 41318
rect 4346 41266 4358 41318
rect 4410 41266 4422 41318
rect 4474 41266 4486 41318
rect 4538 41266 35014 41318
rect 35066 41266 35078 41318
rect 35130 41266 35142 41318
rect 35194 41266 35206 41318
rect 35258 41266 58848 41318
rect 1152 41244 58848 41266
rect 8275 40976 8333 40982
rect 8275 40942 8287 40976
rect 8321 40973 8333 40976
rect 8563 40976 8621 40982
rect 8563 40973 8575 40976
rect 8321 40945 8575 40973
rect 8321 40942 8333 40945
rect 8275 40936 8333 40942
rect 8563 40942 8575 40945
rect 8609 40973 8621 40976
rect 44560 40973 44566 40985
rect 8609 40945 17294 40973
rect 8609 40942 8621 40945
rect 8563 40936 8621 40942
rect 12211 40902 12269 40908
rect 12211 40868 12223 40902
rect 12257 40868 12269 40902
rect 12211 40862 12269 40868
rect 12226 40763 12254 40862
rect 17266 40825 17294 40945
rect 27346 40945 44566 40973
rect 19603 40902 19661 40908
rect 19603 40868 19615 40902
rect 19649 40899 19661 40902
rect 19891 40902 19949 40908
rect 19891 40899 19903 40902
rect 19649 40871 19903 40899
rect 19649 40868 19661 40871
rect 19603 40862 19661 40868
rect 19891 40868 19903 40871
rect 19937 40899 19949 40902
rect 26128 40899 26134 40911
rect 19937 40871 26134 40899
rect 19937 40868 19949 40871
rect 19891 40862 19949 40868
rect 26128 40859 26134 40871
rect 26186 40859 26192 40911
rect 27346 40825 27374 40945
rect 44560 40933 44566 40945
rect 44618 40933 44624 40985
rect 40531 40902 40589 40908
rect 40531 40899 40543 40902
rect 17266 40797 27374 40825
rect 40354 40871 40543 40899
rect 12115 40754 12173 40760
rect 12115 40720 12127 40754
rect 12161 40751 12173 40754
rect 12208 40751 12214 40763
rect 12161 40723 12214 40751
rect 12161 40720 12173 40723
rect 12115 40714 12173 40720
rect 12208 40711 12214 40723
rect 12266 40711 12272 40763
rect 25360 40711 25366 40763
rect 25418 40751 25424 40763
rect 40354 40760 40382 40871
rect 40531 40868 40543 40871
rect 40577 40868 40589 40902
rect 40531 40862 40589 40868
rect 40339 40754 40397 40760
rect 40339 40751 40351 40754
rect 25418 40723 40351 40751
rect 25418 40711 25424 40723
rect 40339 40720 40351 40723
rect 40385 40720 40397 40754
rect 40339 40714 40397 40720
rect 1152 40652 58848 40674
rect 1152 40600 19654 40652
rect 19706 40600 19718 40652
rect 19770 40600 19782 40652
rect 19834 40600 19846 40652
rect 19898 40600 50374 40652
rect 50426 40600 50438 40652
rect 50490 40600 50502 40652
rect 50554 40600 50566 40652
rect 50618 40600 58848 40652
rect 1152 40578 58848 40600
rect 29104 40045 29110 40097
rect 29162 40085 29168 40097
rect 45043 40088 45101 40094
rect 45043 40085 45055 40088
rect 29162 40057 45055 40085
rect 29162 40045 29168 40057
rect 45043 40054 45055 40057
rect 45089 40085 45101 40088
rect 45235 40088 45293 40094
rect 45235 40085 45247 40088
rect 45089 40057 45247 40085
rect 45089 40054 45101 40057
rect 45043 40048 45101 40054
rect 45235 40054 45247 40057
rect 45281 40054 45293 40088
rect 45235 40048 45293 40054
rect 1152 39986 58848 40008
rect 1152 39934 4294 39986
rect 4346 39934 4358 39986
rect 4410 39934 4422 39986
rect 4474 39934 4486 39986
rect 4538 39934 35014 39986
rect 35066 39934 35078 39986
rect 35130 39934 35142 39986
rect 35194 39934 35206 39986
rect 35258 39934 58848 39986
rect 1152 39912 58848 39934
rect 45811 39866 45869 39872
rect 45811 39832 45823 39866
rect 45857 39863 45869 39866
rect 46864 39863 46870 39875
rect 45857 39835 46870 39863
rect 45857 39832 45869 39835
rect 45811 39826 45869 39832
rect 46864 39823 46870 39835
rect 46922 39823 46928 39875
rect 7123 39570 7181 39576
rect 7123 39567 7135 39570
rect 6754 39539 7135 39567
rect 6754 39431 6782 39539
rect 7123 39536 7135 39539
rect 7169 39536 7181 39570
rect 7123 39530 7181 39536
rect 23635 39570 23693 39576
rect 23635 39536 23647 39570
rect 23681 39567 23693 39570
rect 32464 39567 32470 39579
rect 23681 39539 32470 39567
rect 23681 39536 23693 39539
rect 23635 39530 23693 39536
rect 32464 39527 32470 39539
rect 32522 39527 32528 39579
rect 43795 39570 43853 39576
rect 43795 39536 43807 39570
rect 43841 39567 43853 39570
rect 44080 39567 44086 39579
rect 43841 39539 44086 39567
rect 43841 39536 43853 39539
rect 43795 39530 43853 39536
rect 44080 39527 44086 39539
rect 44138 39527 44144 39579
rect 49555 39570 49613 39576
rect 49555 39567 49567 39570
rect 49378 39539 49567 39567
rect 30640 39453 30646 39505
rect 30698 39493 30704 39505
rect 49378 39502 49406 39539
rect 49555 39536 49567 39539
rect 49601 39536 49613 39570
rect 49555 39530 49613 39536
rect 49363 39496 49421 39502
rect 49363 39493 49375 39496
rect 30698 39465 49375 39493
rect 30698 39453 30704 39465
rect 49363 39462 49375 39465
rect 49409 39462 49421 39496
rect 49363 39456 49421 39462
rect 6736 39419 6742 39431
rect 6697 39391 6742 39419
rect 6736 39379 6742 39391
rect 6794 39379 6800 39431
rect 1152 39320 58848 39342
rect 1152 39268 19654 39320
rect 19706 39268 19718 39320
rect 19770 39268 19782 39320
rect 19834 39268 19846 39320
rect 19898 39268 50374 39320
rect 50426 39268 50438 39320
rect 50490 39268 50502 39320
rect 50554 39268 50566 39320
rect 50618 39268 58848 39320
rect 1152 39246 58848 39268
rect 44080 39157 44086 39209
rect 44138 39197 44144 39209
rect 53200 39197 53206 39209
rect 44138 39169 53206 39197
rect 44138 39157 44144 39169
rect 53200 39157 53206 39169
rect 53258 39157 53264 39209
rect 15280 38827 15286 38839
rect 15241 38799 15286 38827
rect 15280 38787 15286 38799
rect 15338 38787 15344 38839
rect 21904 38713 21910 38765
rect 21962 38753 21968 38765
rect 47923 38756 47981 38762
rect 47923 38753 47935 38756
rect 21962 38725 47935 38753
rect 21962 38713 21968 38725
rect 47923 38722 47935 38725
rect 47969 38753 47981 38756
rect 48019 38756 48077 38762
rect 48019 38753 48031 38756
rect 47969 38725 48031 38753
rect 47969 38722 47981 38725
rect 47923 38716 47981 38722
rect 48019 38722 48031 38725
rect 48065 38722 48077 38756
rect 48019 38716 48077 38722
rect 56464 38713 56470 38765
rect 56522 38753 56528 38765
rect 56947 38756 57005 38762
rect 56947 38753 56959 38756
rect 56522 38725 56959 38753
rect 56522 38713 56528 38725
rect 56947 38722 56959 38725
rect 56993 38753 57005 38756
rect 57139 38756 57197 38762
rect 57139 38753 57151 38756
rect 56993 38725 57151 38753
rect 56993 38722 57005 38725
rect 56947 38716 57005 38722
rect 57139 38722 57151 38725
rect 57185 38722 57197 38756
rect 57139 38716 57197 38722
rect 1152 38654 58848 38676
rect 1152 38602 4294 38654
rect 4346 38602 4358 38654
rect 4410 38602 4422 38654
rect 4474 38602 4486 38654
rect 4538 38602 35014 38654
rect 35066 38602 35078 38654
rect 35130 38602 35142 38654
rect 35194 38602 35206 38654
rect 35258 38602 58848 38654
rect 1152 38580 58848 38602
rect 30739 38534 30797 38540
rect 30739 38500 30751 38534
rect 30785 38531 30797 38534
rect 39568 38531 39574 38543
rect 30785 38503 39574 38531
rect 30785 38500 30797 38503
rect 30739 38494 30797 38500
rect 39568 38491 39574 38503
rect 39626 38491 39632 38543
rect 13552 38269 13558 38321
rect 13610 38309 13616 38321
rect 38608 38309 38614 38321
rect 13610 38281 22334 38309
rect 13610 38269 13616 38281
rect 14419 38238 14477 38244
rect 14419 38235 14431 38238
rect 14242 38207 14431 38235
rect 14242 38099 14270 38207
rect 14419 38204 14431 38207
rect 14465 38204 14477 38238
rect 18259 38238 18317 38244
rect 18259 38235 18271 38238
rect 14419 38198 14477 38204
rect 18082 38207 18271 38235
rect 18082 38099 18110 38207
rect 18259 38204 18271 38207
rect 18305 38204 18317 38238
rect 18259 38198 18317 38204
rect 22306 38161 22334 38281
rect 27346 38281 38614 38309
rect 23923 38238 23981 38244
rect 23923 38204 23935 38238
rect 23969 38235 23981 38238
rect 27346 38235 27374 38281
rect 38608 38269 38614 38281
rect 38666 38269 38672 38321
rect 23969 38207 27374 38235
rect 38707 38238 38765 38244
rect 23969 38204 23981 38207
rect 23923 38198 23981 38204
rect 38707 38204 38719 38238
rect 38753 38204 38765 38238
rect 38707 38198 38765 38204
rect 29875 38164 29933 38170
rect 29875 38161 29887 38164
rect 22306 38133 29887 38161
rect 29875 38130 29887 38133
rect 29921 38130 29933 38164
rect 29875 38124 29933 38130
rect 14224 38087 14230 38099
rect 14185 38059 14230 38087
rect 14224 38047 14230 38059
rect 14282 38047 14288 38099
rect 18064 38087 18070 38099
rect 18025 38059 18070 38087
rect 18064 38047 18070 38059
rect 18122 38047 18128 38099
rect 38320 38047 38326 38099
rect 38378 38087 38384 38099
rect 38515 38090 38573 38096
rect 38515 38087 38527 38090
rect 38378 38059 38527 38087
rect 38378 38047 38384 38059
rect 38515 38056 38527 38059
rect 38561 38087 38573 38090
rect 38722 38087 38750 38198
rect 38561 38059 38750 38087
rect 38561 38056 38573 38059
rect 38515 38050 38573 38056
rect 1152 37988 58848 38010
rect 1152 37936 19654 37988
rect 19706 37936 19718 37988
rect 19770 37936 19782 37988
rect 19834 37936 19846 37988
rect 19898 37936 50374 37988
rect 50426 37936 50438 37988
rect 50490 37936 50502 37988
rect 50554 37936 50566 37988
rect 50618 37936 58848 37988
rect 1152 37914 58848 37936
rect 6832 37825 6838 37877
rect 6890 37865 6896 37877
rect 18064 37865 18070 37877
rect 6890 37837 18070 37865
rect 6890 37825 6896 37837
rect 18064 37825 18070 37837
rect 18122 37825 18128 37877
rect 32947 37498 33005 37504
rect 32947 37464 32959 37498
rect 32993 37495 33005 37498
rect 32993 37467 33278 37495
rect 32993 37464 33005 37467
rect 32947 37458 33005 37464
rect 10963 37424 11021 37430
rect 10963 37390 10975 37424
rect 11009 37421 11021 37424
rect 11251 37424 11309 37430
rect 11251 37421 11263 37424
rect 11009 37393 11263 37421
rect 11009 37390 11021 37393
rect 10963 37384 11021 37390
rect 11251 37390 11263 37393
rect 11297 37421 11309 37424
rect 11344 37421 11350 37433
rect 11297 37393 11350 37421
rect 11297 37390 11309 37393
rect 11251 37384 11309 37390
rect 11344 37381 11350 37393
rect 11402 37381 11408 37433
rect 33250 37430 33278 37467
rect 33235 37424 33293 37430
rect 33235 37421 33247 37424
rect 33145 37393 33247 37421
rect 33235 37390 33247 37393
rect 33281 37421 33293 37424
rect 51280 37421 51286 37433
rect 33281 37393 51286 37421
rect 33281 37390 33293 37393
rect 33235 37384 33293 37390
rect 51280 37381 51286 37393
rect 51338 37381 51344 37433
rect 55888 37381 55894 37433
rect 55946 37421 55952 37433
rect 57331 37424 57389 37430
rect 57331 37421 57343 37424
rect 55946 37393 57343 37421
rect 55946 37381 55952 37393
rect 57331 37390 57343 37393
rect 57377 37390 57389 37424
rect 57331 37384 57389 37390
rect 1152 37322 58848 37344
rect 1152 37270 4294 37322
rect 4346 37270 4358 37322
rect 4410 37270 4422 37322
rect 4474 37270 4486 37322
rect 4538 37270 35014 37322
rect 35066 37270 35078 37322
rect 35130 37270 35142 37322
rect 35194 37270 35206 37322
rect 35258 37270 58848 37322
rect 1152 37248 58848 37270
rect 15088 36863 15094 36915
rect 15146 36903 15152 36915
rect 43987 36906 44045 36912
rect 43987 36903 43999 36906
rect 15146 36875 43999 36903
rect 15146 36863 15152 36875
rect 43987 36872 43999 36875
rect 44033 36903 44045 36906
rect 44179 36906 44237 36912
rect 44179 36903 44191 36906
rect 44033 36875 44191 36903
rect 44033 36872 44045 36875
rect 43987 36866 44045 36872
rect 44179 36872 44191 36875
rect 44225 36872 44237 36906
rect 44179 36866 44237 36872
rect 1152 36656 58848 36678
rect 1152 36604 19654 36656
rect 19706 36604 19718 36656
rect 19770 36604 19782 36656
rect 19834 36604 19846 36656
rect 19898 36604 50374 36656
rect 50426 36604 50438 36656
rect 50490 36604 50502 36656
rect 50554 36604 50566 36656
rect 50618 36604 58848 36656
rect 1152 36582 58848 36604
rect 14992 36089 14998 36101
rect 14953 36061 14998 36089
rect 14992 36049 14998 36061
rect 15050 36089 15056 36101
rect 15187 36092 15245 36098
rect 15187 36089 15199 36092
rect 15050 36061 15199 36089
rect 15050 36049 15056 36061
rect 15187 36058 15199 36061
rect 15233 36058 15245 36092
rect 15187 36052 15245 36058
rect 40051 36092 40109 36098
rect 40051 36058 40063 36092
rect 40097 36089 40109 36092
rect 40339 36092 40397 36098
rect 40339 36089 40351 36092
rect 40097 36061 40351 36089
rect 40097 36058 40109 36061
rect 40051 36052 40109 36058
rect 40339 36058 40351 36061
rect 40385 36089 40397 36092
rect 46192 36089 46198 36101
rect 40385 36061 46198 36089
rect 40385 36058 40397 36061
rect 40339 36052 40397 36058
rect 46192 36049 46198 36061
rect 46250 36049 46256 36101
rect 46288 36049 46294 36101
rect 46346 36089 46352 36101
rect 46387 36092 46445 36098
rect 46387 36089 46399 36092
rect 46346 36061 46399 36089
rect 46346 36049 46352 36061
rect 46387 36058 46399 36061
rect 46433 36089 46445 36092
rect 46579 36092 46637 36098
rect 46579 36089 46591 36092
rect 46433 36061 46591 36089
rect 46433 36058 46445 36061
rect 46387 36052 46445 36058
rect 46579 36058 46591 36061
rect 46625 36058 46637 36092
rect 46579 36052 46637 36058
rect 1152 35990 58848 36012
rect 1152 35938 4294 35990
rect 4346 35938 4358 35990
rect 4410 35938 4422 35990
rect 4474 35938 4486 35990
rect 4538 35938 35014 35990
rect 35066 35938 35078 35990
rect 35130 35938 35142 35990
rect 35194 35938 35206 35990
rect 35258 35938 58848 35990
rect 1152 35916 58848 35938
rect 31024 35679 31030 35731
rect 31082 35719 31088 35731
rect 36019 35722 36077 35728
rect 36019 35719 36031 35722
rect 31082 35691 36031 35719
rect 31082 35679 31088 35691
rect 36019 35688 36031 35691
rect 36065 35688 36077 35722
rect 36019 35682 36077 35688
rect 8560 35605 8566 35657
rect 8618 35645 8624 35657
rect 52051 35648 52109 35654
rect 52051 35645 52063 35648
rect 8618 35617 52063 35645
rect 8618 35605 8624 35617
rect 52051 35614 52063 35617
rect 52097 35614 52109 35648
rect 52051 35608 52109 35614
rect 33235 35574 33293 35580
rect 33235 35540 33247 35574
rect 33281 35571 33293 35574
rect 33520 35571 33526 35583
rect 33281 35543 33526 35571
rect 33281 35540 33293 35543
rect 33235 35534 33293 35540
rect 33520 35531 33526 35543
rect 33578 35531 33584 35583
rect 1152 35324 58848 35346
rect 1152 35272 19654 35324
rect 19706 35272 19718 35324
rect 19770 35272 19782 35324
rect 19834 35272 19846 35324
rect 19898 35272 50374 35324
rect 50426 35272 50438 35324
rect 50490 35272 50502 35324
rect 50554 35272 50566 35324
rect 50618 35272 58848 35324
rect 1152 35250 58848 35272
rect 27346 34803 37454 34831
rect 14800 34757 14806 34769
rect 14761 34729 14806 34757
rect 14800 34717 14806 34729
rect 14858 34757 14864 34769
rect 15091 34760 15149 34766
rect 15091 34757 15103 34760
rect 14858 34729 15103 34757
rect 14858 34717 14864 34729
rect 15091 34726 15103 34729
rect 15137 34726 15149 34760
rect 15091 34720 15149 34726
rect 19024 34717 19030 34769
rect 19082 34757 19088 34769
rect 27346 34757 27374 34803
rect 19082 34729 27374 34757
rect 32659 34760 32717 34766
rect 19082 34717 19088 34729
rect 32659 34726 32671 34760
rect 32705 34757 32717 34760
rect 32752 34757 32758 34769
rect 32705 34729 32758 34757
rect 32705 34726 32717 34729
rect 32659 34720 32717 34726
rect 32752 34717 32758 34729
rect 32810 34717 32816 34769
rect 37426 34757 37454 34803
rect 41491 34760 41549 34766
rect 41491 34757 41503 34760
rect 37426 34729 41503 34757
rect 41491 34726 41503 34729
rect 41537 34726 41549 34760
rect 41491 34720 41549 34726
rect 1152 34658 58848 34680
rect 1152 34606 4294 34658
rect 4346 34606 4358 34658
rect 4410 34606 4422 34658
rect 4474 34606 4486 34658
rect 4538 34606 35014 34658
rect 35066 34606 35078 34658
rect 35130 34606 35142 34658
rect 35194 34606 35206 34658
rect 35258 34606 58848 34658
rect 1152 34584 58848 34606
rect 24016 34199 24022 34251
rect 24074 34239 24080 34251
rect 47251 34242 47309 34248
rect 47251 34239 47263 34242
rect 24074 34211 47263 34239
rect 24074 34199 24080 34211
rect 47251 34208 47263 34211
rect 47297 34208 47309 34242
rect 47251 34202 47309 34208
rect 1152 33992 58848 34014
rect 1152 33940 19654 33992
rect 19706 33940 19718 33992
rect 19770 33940 19782 33992
rect 19834 33940 19846 33992
rect 19898 33940 50374 33992
rect 50426 33940 50438 33992
rect 50490 33940 50502 33992
rect 50554 33940 50566 33992
rect 50618 33940 58848 33992
rect 1152 33918 58848 33940
rect 1840 33607 1846 33659
rect 1898 33647 1904 33659
rect 28240 33647 28246 33659
rect 1898 33619 28246 33647
rect 1898 33607 1904 33619
rect 28240 33607 28246 33619
rect 28298 33607 28304 33659
rect 28336 33459 28342 33511
rect 28394 33499 28400 33511
rect 57139 33502 57197 33508
rect 57139 33499 57151 33502
rect 28394 33471 57151 33499
rect 28394 33459 28400 33471
rect 57139 33468 57151 33471
rect 57185 33499 57197 33502
rect 57331 33502 57389 33508
rect 57331 33499 57343 33502
rect 57185 33471 57343 33499
rect 57185 33468 57197 33471
rect 57139 33462 57197 33468
rect 57331 33468 57343 33471
rect 57377 33468 57389 33502
rect 57331 33462 57389 33468
rect 12688 33385 12694 33437
rect 12746 33425 12752 33437
rect 47728 33425 47734 33437
rect 12746 33397 47734 33425
rect 12746 33385 12752 33397
rect 47728 33385 47734 33397
rect 47786 33385 47792 33437
rect 1152 33326 58848 33348
rect 1152 33274 4294 33326
rect 4346 33274 4358 33326
rect 4410 33274 4422 33326
rect 4474 33274 4486 33326
rect 4538 33274 35014 33326
rect 35066 33274 35078 33326
rect 35130 33274 35142 33326
rect 35194 33274 35206 33326
rect 35258 33274 58848 33326
rect 1152 33252 58848 33274
rect 19027 33206 19085 33212
rect 19027 33172 19039 33206
rect 19073 33203 19085 33206
rect 47728 33203 47734 33215
rect 19073 33175 47582 33203
rect 47689 33175 47734 33203
rect 19073 33172 19085 33175
rect 19027 33166 19085 33172
rect 28240 33129 28246 33141
rect 28201 33101 28246 33129
rect 28240 33089 28246 33101
rect 28298 33089 28304 33141
rect 47554 33129 47582 33175
rect 47728 33163 47734 33175
rect 47786 33163 47792 33215
rect 56560 33203 56566 33215
rect 47842 33175 56566 33203
rect 47842 33129 47870 33175
rect 56560 33163 56566 33175
rect 56618 33163 56624 33215
rect 47554 33101 47870 33129
rect 42352 32907 42358 32919
rect 42313 32879 42358 32907
rect 42352 32867 42358 32879
rect 42410 32867 42416 32919
rect 1152 32660 58848 32682
rect 1152 32608 19654 32660
rect 19706 32608 19718 32660
rect 19770 32608 19782 32660
rect 19834 32608 19846 32660
rect 19898 32608 50374 32660
rect 50426 32608 50438 32660
rect 50490 32608 50502 32660
rect 50554 32608 50566 32660
rect 50618 32608 58848 32660
rect 1152 32586 58848 32608
rect 19027 32540 19085 32546
rect 19027 32506 19039 32540
rect 19073 32537 19085 32540
rect 20560 32537 20566 32549
rect 19073 32509 20566 32537
rect 19073 32506 19085 32509
rect 19027 32500 19085 32506
rect 20560 32497 20566 32509
rect 20618 32497 20624 32549
rect 13936 32093 13942 32105
rect 13897 32065 13942 32093
rect 13936 32053 13942 32065
rect 13994 32053 14000 32105
rect 30931 32096 30989 32102
rect 30931 32062 30943 32096
rect 30977 32093 30989 32096
rect 31216 32093 31222 32105
rect 30977 32065 31222 32093
rect 30977 32062 30989 32065
rect 30931 32056 30989 32062
rect 31216 32053 31222 32065
rect 31274 32053 31280 32105
rect 34099 32096 34157 32102
rect 34099 32062 34111 32096
rect 34145 32093 34157 32096
rect 34768 32093 34774 32105
rect 34145 32065 34774 32093
rect 34145 32062 34157 32065
rect 34099 32056 34157 32062
rect 34768 32053 34774 32065
rect 34826 32053 34832 32105
rect 1152 31994 58848 32016
rect 1152 31942 4294 31994
rect 4346 31942 4358 31994
rect 4410 31942 4422 31994
rect 4474 31942 4486 31994
rect 4538 31942 35014 31994
rect 35066 31942 35078 31994
rect 35130 31942 35142 31994
rect 35194 31942 35206 31994
rect 35258 31942 58848 31994
rect 1152 31920 58848 31942
rect 39859 31874 39917 31880
rect 39859 31840 39871 31874
rect 39905 31871 39917 31874
rect 41104 31871 41110 31883
rect 39905 31843 41110 31871
rect 39905 31840 39917 31843
rect 39859 31834 39917 31840
rect 41104 31831 41110 31843
rect 41162 31831 41168 31883
rect 48304 31683 48310 31735
rect 48362 31723 48368 31735
rect 58003 31726 58061 31732
rect 58003 31723 58015 31726
rect 48362 31695 58015 31723
rect 48362 31683 48368 31695
rect 58003 31692 58015 31695
rect 58049 31692 58061 31726
rect 58003 31686 58061 31692
rect 1152 31328 58848 31350
rect 1152 31276 19654 31328
rect 19706 31276 19718 31328
rect 19770 31276 19782 31328
rect 19834 31276 19846 31328
rect 19898 31276 50374 31328
rect 50426 31276 50438 31328
rect 50490 31276 50502 31328
rect 50554 31276 50566 31328
rect 50618 31276 58848 31328
rect 1152 31254 58848 31276
rect 16915 30838 16973 30844
rect 16915 30804 16927 30838
rect 16961 30835 16973 30838
rect 45136 30835 45142 30847
rect 16961 30807 45142 30835
rect 16961 30804 16973 30807
rect 16915 30798 16973 30804
rect 45136 30795 45142 30807
rect 45194 30795 45200 30847
rect 17587 30764 17645 30770
rect 17587 30730 17599 30764
rect 17633 30761 17645 30764
rect 17680 30761 17686 30773
rect 17633 30733 17686 30761
rect 17633 30730 17645 30733
rect 17587 30724 17645 30730
rect 17680 30721 17686 30733
rect 17738 30721 17744 30773
rect 1152 30662 58848 30684
rect 1152 30610 4294 30662
rect 4346 30610 4358 30662
rect 4410 30610 4422 30662
rect 4474 30610 4486 30662
rect 4538 30610 35014 30662
rect 35066 30610 35078 30662
rect 35130 30610 35142 30662
rect 35194 30610 35206 30662
rect 35258 30610 58848 30662
rect 1152 30588 58848 30610
rect 25456 30351 25462 30403
rect 25514 30391 25520 30403
rect 31795 30394 31853 30400
rect 31795 30391 31807 30394
rect 25514 30363 31807 30391
rect 25514 30351 25520 30363
rect 31795 30360 31807 30363
rect 31841 30360 31853 30394
rect 31795 30354 31853 30360
rect 29968 30317 29974 30329
rect 29929 30289 29974 30317
rect 29968 30277 29974 30289
rect 30026 30277 30032 30329
rect 1152 29996 58848 30018
rect 1152 29944 19654 29996
rect 19706 29944 19718 29996
rect 19770 29944 19782 29996
rect 19834 29944 19846 29996
rect 19898 29944 50374 29996
rect 50426 29944 50438 29996
rect 50490 29944 50502 29996
rect 50554 29944 50566 29996
rect 50618 29944 58848 29996
rect 1152 29922 58848 29944
rect 6352 29611 6358 29663
rect 6410 29651 6416 29663
rect 55504 29651 55510 29663
rect 6410 29623 55510 29651
rect 6410 29611 6416 29623
rect 55504 29611 55510 29623
rect 55562 29611 55568 29663
rect 1936 29537 1942 29589
rect 1994 29577 2000 29589
rect 14128 29577 14134 29589
rect 1994 29549 14134 29577
rect 1994 29537 2000 29549
rect 14128 29537 14134 29549
rect 14186 29537 14192 29589
rect 52435 29580 52493 29586
rect 52435 29546 52447 29580
rect 52481 29546 52493 29580
rect 52435 29540 52493 29546
rect 11536 29463 11542 29515
rect 11594 29503 11600 29515
rect 52243 29506 52301 29512
rect 52243 29503 52255 29506
rect 11594 29475 52255 29503
rect 11594 29463 11600 29475
rect 52243 29472 52255 29475
rect 52289 29503 52301 29506
rect 52450 29503 52478 29540
rect 52289 29475 52478 29503
rect 52289 29472 52301 29475
rect 52243 29466 52301 29472
rect 17776 29429 17782 29441
rect 17737 29401 17782 29429
rect 17776 29389 17782 29401
rect 17834 29389 17840 29441
rect 19216 29429 19222 29441
rect 19177 29401 19222 29429
rect 19216 29389 19222 29401
rect 19274 29389 19280 29441
rect 40336 29429 40342 29441
rect 40297 29401 40342 29429
rect 40336 29389 40342 29401
rect 40394 29389 40400 29441
rect 49936 29389 49942 29441
rect 49994 29429 50000 29441
rect 50035 29432 50093 29438
rect 50035 29429 50047 29432
rect 49994 29401 50047 29429
rect 49994 29389 50000 29401
rect 50035 29398 50047 29401
rect 50081 29398 50093 29432
rect 50035 29392 50093 29398
rect 50608 29389 50614 29441
rect 50666 29429 50672 29441
rect 53683 29432 53741 29438
rect 53683 29429 53695 29432
rect 50666 29401 53695 29429
rect 50666 29389 50672 29401
rect 53683 29398 53695 29401
rect 53729 29398 53741 29432
rect 53683 29392 53741 29398
rect 54547 29432 54605 29438
rect 54547 29398 54559 29432
rect 54593 29429 54605 29432
rect 54640 29429 54646 29441
rect 54593 29401 54646 29429
rect 54593 29398 54605 29401
rect 54547 29392 54605 29398
rect 54640 29389 54646 29401
rect 54698 29389 54704 29441
rect 55696 29429 55702 29441
rect 55657 29401 55702 29429
rect 55696 29389 55702 29401
rect 55754 29389 55760 29441
rect 1152 29330 58848 29352
rect 1152 29278 4294 29330
rect 4346 29278 4358 29330
rect 4410 29278 4422 29330
rect 4474 29278 4486 29330
rect 4538 29278 35014 29330
rect 35066 29278 35078 29330
rect 35130 29278 35142 29330
rect 35194 29278 35206 29330
rect 35258 29278 58848 29330
rect 1152 29256 58848 29278
rect 9040 29167 9046 29219
rect 9098 29167 9104 29219
rect 14128 29167 14134 29219
rect 14186 29207 14192 29219
rect 14227 29210 14285 29216
rect 14227 29207 14239 29210
rect 14186 29179 14239 29207
rect 14186 29167 14192 29179
rect 14227 29176 14239 29179
rect 14273 29207 14285 29210
rect 14273 29179 14462 29207
rect 14273 29176 14285 29179
rect 14227 29170 14285 29176
rect 8368 29093 8374 29145
rect 8426 29133 8432 29145
rect 8426 29105 8558 29133
rect 8426 29093 8432 29105
rect 8530 28837 8558 29105
rect 14434 29068 14462 29179
rect 22672 29167 22678 29219
rect 22730 29207 22736 29219
rect 50608 29207 50614 29219
rect 22730 29179 50614 29207
rect 22730 29167 22736 29179
rect 50608 29167 50614 29179
rect 50666 29167 50672 29219
rect 55504 29167 55510 29219
rect 55562 29207 55568 29219
rect 55699 29210 55757 29216
rect 55699 29207 55711 29210
rect 55562 29179 55711 29207
rect 55562 29167 55568 29179
rect 55699 29176 55711 29179
rect 55745 29207 55757 29210
rect 55891 29210 55949 29216
rect 55891 29207 55903 29210
rect 55745 29179 55903 29207
rect 55745 29176 55757 29179
rect 55699 29170 55757 29176
rect 55891 29176 55903 29179
rect 55937 29176 55949 29210
rect 55891 29170 55949 29176
rect 14419 29062 14477 29068
rect 14419 29028 14431 29062
rect 14465 29028 14477 29062
rect 14419 29022 14477 29028
rect 41296 28945 41302 28997
rect 41354 28985 41360 28997
rect 46867 28988 46925 28994
rect 46867 28985 46879 28988
rect 41354 28957 46879 28985
rect 41354 28945 41360 28957
rect 46867 28954 46879 28957
rect 46913 28954 46925 28988
rect 46867 28948 46925 28954
rect 15280 28911 15286 28923
rect 15241 28883 15286 28911
rect 15280 28871 15286 28883
rect 15338 28871 15344 28923
rect 44755 28914 44813 28920
rect 44755 28880 44767 28914
rect 44801 28911 44813 28914
rect 44848 28911 44854 28923
rect 44801 28883 44854 28911
rect 44801 28880 44813 28883
rect 44755 28874 44813 28880
rect 44848 28871 44854 28883
rect 44906 28871 44912 28923
rect 8400 28809 8558 28837
rect 8752 28723 8758 28775
rect 8810 28723 8816 28775
rect 1152 28664 58848 28686
rect 1152 28612 19654 28664
rect 19706 28612 19718 28664
rect 19770 28612 19782 28664
rect 19834 28612 19846 28664
rect 19898 28612 50374 28664
rect 50426 28612 50438 28664
rect 50490 28612 50502 28664
rect 50554 28612 50566 28664
rect 50618 28612 58848 28664
rect 1152 28590 58848 28612
rect 2896 28131 2902 28183
rect 2954 28171 2960 28183
rect 38131 28174 38189 28180
rect 38131 28171 38143 28174
rect 2954 28143 38143 28171
rect 2954 28131 2960 28143
rect 38131 28140 38143 28143
rect 38177 28171 38189 28174
rect 38323 28174 38381 28180
rect 38323 28171 38335 28174
rect 38177 28143 38335 28171
rect 38177 28140 38189 28143
rect 38131 28134 38189 28140
rect 38323 28140 38335 28143
rect 38369 28140 38381 28174
rect 38323 28134 38381 28140
rect 20371 28100 20429 28106
rect 20371 28066 20383 28100
rect 20417 28097 20429 28100
rect 20464 28097 20470 28109
rect 20417 28069 20470 28097
rect 20417 28066 20429 28069
rect 20371 28060 20429 28066
rect 20464 28057 20470 28069
rect 20522 28057 20528 28109
rect 41776 28097 41782 28109
rect 41737 28069 41782 28097
rect 41776 28057 41782 28069
rect 41834 28057 41840 28109
rect 1152 27998 58848 28020
rect 1152 27946 4294 27998
rect 4346 27946 4358 27998
rect 4410 27946 4422 27998
rect 4474 27946 4486 27998
rect 4538 27946 35014 27998
rect 35066 27946 35078 27998
rect 35130 27946 35142 27998
rect 35194 27946 35206 27998
rect 35258 27946 58848 27998
rect 1152 27924 58848 27946
rect 7120 27835 7126 27887
rect 7178 27875 7184 27887
rect 7178 27847 7982 27875
rect 7178 27835 7184 27847
rect 7954 27713 7982 27847
rect 26416 27835 26422 27887
rect 26474 27875 26480 27887
rect 41776 27875 41782 27887
rect 26474 27847 41782 27875
rect 26474 27835 26480 27847
rect 41776 27835 41782 27847
rect 41834 27835 41840 27887
rect 8368 27727 8374 27739
rect 8256 27699 8374 27727
rect 8368 27687 8374 27699
rect 8426 27687 8432 27739
rect 14320 27579 14326 27591
rect 14281 27551 14326 27579
rect 14320 27539 14326 27551
rect 14378 27539 14384 27591
rect 25072 27539 25078 27591
rect 25130 27579 25136 27591
rect 55219 27582 55277 27588
rect 55219 27579 55231 27582
rect 25130 27551 55231 27579
rect 25130 27539 25136 27551
rect 55219 27548 55231 27551
rect 55265 27579 55277 27582
rect 55411 27582 55469 27588
rect 55411 27579 55423 27582
rect 55265 27551 55423 27579
rect 55265 27548 55277 27551
rect 55219 27542 55277 27548
rect 55411 27548 55423 27551
rect 55457 27548 55469 27582
rect 55411 27542 55469 27548
rect 8848 27431 8854 27443
rect 8640 27403 8854 27431
rect 8848 27391 8854 27403
rect 8906 27391 8912 27443
rect 1152 27332 58848 27354
rect 1152 27280 19654 27332
rect 19706 27280 19718 27332
rect 19770 27280 19782 27332
rect 19834 27280 19846 27332
rect 19898 27280 50374 27332
rect 50426 27280 50438 27332
rect 50490 27280 50502 27332
rect 50554 27280 50566 27332
rect 50618 27280 58848 27332
rect 1152 27258 58848 27280
rect 14803 26916 14861 26922
rect 14803 26882 14815 26916
rect 14849 26913 14861 26916
rect 15091 26916 15149 26922
rect 15091 26913 15103 26916
rect 14849 26885 15103 26913
rect 14849 26882 14861 26885
rect 14803 26876 14861 26882
rect 15091 26882 15103 26885
rect 15137 26913 15149 26916
rect 15137 26885 15854 26913
rect 15137 26882 15149 26885
rect 15091 26876 15149 26882
rect 15826 26839 15854 26885
rect 24304 26839 24310 26851
rect 15826 26811 24310 26839
rect 24304 26799 24310 26811
rect 24362 26799 24368 26851
rect 27346 26811 37454 26839
rect 7696 26725 7702 26777
rect 7754 26765 7760 26777
rect 27346 26765 27374 26811
rect 28624 26765 28630 26777
rect 7754 26737 27374 26765
rect 28585 26737 28630 26765
rect 7754 26725 7760 26737
rect 28624 26725 28630 26737
rect 28682 26725 28688 26777
rect 37426 26765 37454 26811
rect 47251 26768 47309 26774
rect 47251 26765 47263 26768
rect 37426 26737 47263 26765
rect 47251 26734 47263 26737
rect 47297 26765 47309 26768
rect 47443 26768 47501 26774
rect 47443 26765 47455 26768
rect 47297 26737 47455 26765
rect 47297 26734 47309 26737
rect 47251 26728 47309 26734
rect 47443 26734 47455 26737
rect 47489 26734 47501 26768
rect 47443 26728 47501 26734
rect 1152 26666 58848 26688
rect 1152 26614 4294 26666
rect 4346 26614 4358 26666
rect 4410 26614 4422 26666
rect 4474 26614 4486 26666
rect 4538 26614 35014 26666
rect 35066 26614 35078 26666
rect 35130 26614 35142 26666
rect 35194 26614 35206 26666
rect 35258 26614 58848 26666
rect 1152 26592 58848 26614
rect 8080 26355 8086 26407
rect 8138 26395 8144 26407
rect 8138 26367 8256 26395
rect 8138 26355 8144 26367
rect 7942 26333 7994 26339
rect 7942 26275 7994 26281
rect 24208 26247 24214 26259
rect 24169 26219 24214 26247
rect 24208 26207 24214 26219
rect 24266 26207 24272 26259
rect 36112 26207 36118 26259
rect 36170 26247 36176 26259
rect 38995 26250 39053 26256
rect 38995 26247 39007 26250
rect 36170 26219 39007 26247
rect 36170 26207 36176 26219
rect 38995 26216 39007 26219
rect 39041 26216 39053 26250
rect 57331 26250 57389 26256
rect 57331 26247 57343 26250
rect 38995 26210 39053 26216
rect 47506 26219 57343 26247
rect 16240 26133 16246 26185
rect 16298 26173 16304 26185
rect 47506 26173 47534 26219
rect 57331 26216 57343 26219
rect 57377 26216 57389 26250
rect 57331 26210 57389 26216
rect 16298 26145 47534 26173
rect 16298 26133 16304 26145
rect 9232 26099 9238 26111
rect 8640 26071 9238 26099
rect 9232 26059 9238 26071
rect 9290 26059 9296 26111
rect 1152 26000 58848 26022
rect 1152 25948 19654 26000
rect 19706 25948 19718 26000
rect 19770 25948 19782 26000
rect 19834 25948 19846 26000
rect 19898 25948 50374 26000
rect 50426 25948 50438 26000
rect 50490 25948 50502 26000
rect 50554 25948 50566 26000
rect 50618 25948 58848 26000
rect 1152 25926 58848 25948
rect 55120 25837 55126 25889
rect 55178 25877 55184 25889
rect 55315 25880 55373 25886
rect 55315 25877 55327 25880
rect 55178 25849 55327 25877
rect 55178 25837 55184 25849
rect 55315 25846 55327 25849
rect 55361 25846 55373 25880
rect 55315 25840 55373 25846
rect 7027 25732 7085 25738
rect 7027 25698 7039 25732
rect 7073 25729 7085 25732
rect 7315 25732 7373 25738
rect 7315 25729 7327 25732
rect 7073 25701 7327 25729
rect 7073 25698 7085 25701
rect 7027 25692 7085 25698
rect 7315 25698 7327 25701
rect 7361 25729 7373 25732
rect 14704 25729 14710 25741
rect 7361 25701 14710 25729
rect 7361 25698 7373 25701
rect 7315 25692 7373 25698
rect 14704 25689 14710 25701
rect 14762 25689 14768 25741
rect 55330 25729 55358 25840
rect 55507 25732 55565 25738
rect 55507 25729 55519 25732
rect 55330 25701 55519 25729
rect 55507 25698 55519 25701
rect 55553 25698 55565 25732
rect 55507 25692 55565 25698
rect 4531 25436 4589 25442
rect 4531 25402 4543 25436
rect 4577 25433 4589 25436
rect 5680 25433 5686 25445
rect 4577 25405 5686 25433
rect 4577 25402 4589 25405
rect 4531 25396 4589 25402
rect 5680 25393 5686 25405
rect 5738 25393 5744 25445
rect 21139 25436 21197 25442
rect 21139 25402 21151 25436
rect 21185 25433 21197 25436
rect 21427 25436 21485 25442
rect 21427 25433 21439 25436
rect 21185 25405 21439 25433
rect 21185 25402 21197 25405
rect 21139 25396 21197 25402
rect 21427 25402 21439 25405
rect 21473 25433 21485 25436
rect 37648 25433 37654 25445
rect 21473 25405 37654 25433
rect 21473 25402 21485 25405
rect 21427 25396 21485 25402
rect 37648 25393 37654 25405
rect 37706 25393 37712 25445
rect 1152 25334 58848 25356
rect 1152 25282 4294 25334
rect 4346 25282 4358 25334
rect 4410 25282 4422 25334
rect 4474 25282 4486 25334
rect 4538 25282 35014 25334
rect 35066 25282 35078 25334
rect 35130 25282 35142 25334
rect 35194 25282 35206 25334
rect 35258 25282 58848 25334
rect 1152 25260 58848 25282
rect 9616 25211 9622 25223
rect 8770 25183 9622 25211
rect 8770 25123 8798 25183
rect 9616 25171 9622 25183
rect 9674 25171 9680 25223
rect 8386 25035 8544 25063
rect 8386 25001 8414 25035
rect 8368 24949 8374 25001
rect 8426 24949 8432 25001
rect 8832 24998 8990 25026
rect 8962 24989 8990 24998
rect 9136 24989 9142 25001
rect 8962 24961 9142 24989
rect 9136 24949 9142 24961
rect 9194 24949 9200 25001
rect 7942 24927 7994 24933
rect 7942 24869 7994 24875
rect 8230 24927 8282 24933
rect 14608 24915 14614 24927
rect 14569 24887 14614 24915
rect 14608 24875 14614 24887
rect 14666 24875 14672 24927
rect 49840 24915 49846 24927
rect 49801 24887 49846 24915
rect 49840 24875 49846 24887
rect 49898 24875 49904 24927
rect 52528 24915 52534 24927
rect 52489 24887 52534 24915
rect 52528 24875 52534 24887
rect 52586 24875 52592 24927
rect 8230 24869 8282 24875
rect 1152 24668 58848 24690
rect 1152 24616 19654 24668
rect 19706 24616 19718 24668
rect 19770 24616 19782 24668
rect 19834 24616 19846 24668
rect 19898 24616 50374 24668
rect 50426 24616 50438 24668
rect 50490 24616 50502 24668
rect 50554 24616 50566 24668
rect 50618 24616 58848 24668
rect 1152 24594 58848 24616
rect 8176 24505 8182 24557
rect 8234 24545 8240 24557
rect 8560 24545 8566 24557
rect 8234 24517 8566 24545
rect 8234 24505 8240 24517
rect 8560 24505 8566 24517
rect 8618 24505 8624 24557
rect 5200 24135 5206 24187
rect 5258 24175 5264 24187
rect 34864 24175 34870 24187
rect 5258 24147 34870 24175
rect 5258 24135 5264 24147
rect 34864 24135 34870 24147
rect 34922 24135 34928 24187
rect 8368 24061 8374 24113
rect 8426 24101 8432 24113
rect 8560 24101 8566 24113
rect 8426 24073 8566 24101
rect 8426 24061 8432 24073
rect 8560 24061 8566 24073
rect 8618 24061 8624 24113
rect 11632 24101 11638 24113
rect 11593 24073 11638 24101
rect 11632 24061 11638 24073
rect 11690 24061 11696 24113
rect 22867 24104 22925 24110
rect 22867 24070 22879 24104
rect 22913 24101 22925 24104
rect 30160 24101 30166 24113
rect 22913 24073 30166 24101
rect 22913 24070 22925 24073
rect 22867 24064 22925 24070
rect 30160 24061 30166 24073
rect 30218 24061 30224 24113
rect 1152 24002 58848 24024
rect 1152 23950 4294 24002
rect 4346 23950 4358 24002
rect 4410 23950 4422 24002
rect 4474 23950 4486 24002
rect 4538 23950 35014 24002
rect 35066 23950 35078 24002
rect 35130 23950 35142 24002
rect 35194 23950 35206 24002
rect 35258 23950 58848 24002
rect 1152 23928 58848 23950
rect 7408 23839 7414 23891
rect 7466 23879 7472 23891
rect 7792 23879 7798 23891
rect 7466 23851 7798 23879
rect 7466 23839 7472 23851
rect 7792 23839 7798 23851
rect 7850 23839 7856 23891
rect 15856 23879 15862 23891
rect 8482 23851 15862 23879
rect 8482 23791 8510 23851
rect 15856 23839 15862 23851
rect 15914 23839 15920 23891
rect 34864 23839 34870 23891
rect 34922 23879 34928 23891
rect 35059 23882 35117 23888
rect 35059 23879 35071 23882
rect 34922 23851 35071 23879
rect 34922 23839 34928 23851
rect 35059 23848 35071 23851
rect 35105 23879 35117 23882
rect 35105 23851 35294 23879
rect 35105 23848 35117 23851
rect 35059 23842 35117 23848
rect 35266 23740 35294 23851
rect 35251 23734 35309 23740
rect 8098 23703 8256 23731
rect 8098 23669 8126 23703
rect 35251 23700 35263 23734
rect 35297 23700 35309 23734
rect 35251 23694 35309 23700
rect 8080 23617 8086 23669
rect 8138 23617 8144 23669
rect 8368 23543 8374 23595
rect 8426 23543 8432 23595
rect 12400 23583 12406 23595
rect 12361 23555 12406 23583
rect 12400 23543 12406 23555
rect 12458 23543 12464 23595
rect 21715 23586 21773 23592
rect 21715 23552 21727 23586
rect 21761 23583 21773 23586
rect 36880 23583 36886 23595
rect 21761 23555 36886 23583
rect 21761 23552 21773 23555
rect 21715 23546 21773 23552
rect 36880 23543 36886 23555
rect 36938 23543 36944 23595
rect 42736 23543 42742 23595
rect 42794 23583 42800 23595
rect 42931 23586 42989 23592
rect 42931 23583 42943 23586
rect 42794 23555 42943 23583
rect 42794 23543 42800 23555
rect 42931 23552 42943 23555
rect 42977 23552 42989 23586
rect 42931 23546 42989 23552
rect 7936 23469 7942 23521
rect 7994 23469 8000 23521
rect 8386 23509 8414 23543
rect 8386 23481 8544 23509
rect 1152 23336 58848 23358
rect 1152 23284 19654 23336
rect 19706 23284 19718 23336
rect 19770 23284 19782 23336
rect 19834 23284 19846 23336
rect 19898 23284 50374 23336
rect 50426 23284 50438 23336
rect 50490 23284 50502 23336
rect 50554 23284 50566 23336
rect 50618 23284 58848 23336
rect 1152 23262 58848 23284
rect 7312 23173 7318 23225
rect 7370 23213 7376 23225
rect 8368 23213 8374 23225
rect 7370 23185 8374 23213
rect 7370 23173 7376 23185
rect 8368 23173 8374 23185
rect 8426 23173 8432 23225
rect 7888 22729 7894 22781
rect 7946 22769 7952 22781
rect 8080 22769 8086 22781
rect 7946 22741 8086 22769
rect 7946 22729 7952 22741
rect 8080 22729 8086 22741
rect 8138 22729 8144 22781
rect 12304 22729 12310 22781
rect 12362 22769 12368 22781
rect 13267 22772 13325 22778
rect 13267 22769 13279 22772
rect 12362 22741 13279 22769
rect 12362 22729 12368 22741
rect 13267 22738 13279 22741
rect 13313 22738 13325 22772
rect 42832 22769 42838 22781
rect 42793 22741 42838 22769
rect 13267 22732 13325 22738
rect 42832 22729 42838 22741
rect 42890 22729 42896 22781
rect 1152 22670 58848 22692
rect 1152 22618 4294 22670
rect 4346 22618 4358 22670
rect 4410 22618 4422 22670
rect 4474 22618 4486 22670
rect 4538 22618 35014 22670
rect 35066 22618 35078 22670
rect 35130 22618 35142 22670
rect 35194 22618 35206 22670
rect 35258 22618 58848 22670
rect 1152 22596 58848 22618
rect 7504 22507 7510 22559
rect 7562 22547 7568 22559
rect 7696 22547 7702 22559
rect 7562 22519 7702 22547
rect 7562 22507 7568 22519
rect 7696 22507 7702 22519
rect 7754 22507 7760 22559
rect 8272 22507 8278 22559
rect 8330 22547 8336 22559
rect 8464 22547 8470 22559
rect 8330 22519 8470 22547
rect 8330 22507 8336 22519
rect 8464 22507 8470 22519
rect 8522 22507 8528 22559
rect 7120 22433 7126 22485
rect 7178 22473 7184 22485
rect 7600 22473 7606 22485
rect 7178 22445 7606 22473
rect 7178 22433 7184 22445
rect 7600 22433 7606 22445
rect 7658 22433 7664 22485
rect 7888 22433 7894 22485
rect 7946 22473 7952 22485
rect 7946 22445 8270 22473
rect 7946 22433 7952 22445
rect 7696 22359 7702 22411
rect 7754 22399 7760 22411
rect 7754 22371 7968 22399
rect 8242 22385 8270 22445
rect 7754 22359 7760 22371
rect 9139 22254 9197 22260
rect 9139 22220 9151 22254
rect 9185 22251 9197 22254
rect 28720 22251 28726 22263
rect 9185 22223 28726 22251
rect 9185 22220 9197 22223
rect 9139 22214 9197 22220
rect 28720 22211 28726 22223
rect 28778 22211 28784 22263
rect 34864 22211 34870 22263
rect 34922 22251 34928 22263
rect 34963 22254 35021 22260
rect 34963 22251 34975 22254
rect 34922 22223 34975 22251
rect 34922 22211 34928 22223
rect 34963 22220 34975 22223
rect 35009 22220 35021 22254
rect 34963 22214 35021 22220
rect 36499 22254 36557 22260
rect 36499 22220 36511 22254
rect 36545 22251 36557 22254
rect 36976 22251 36982 22263
rect 36545 22223 36982 22251
rect 36545 22220 36557 22223
rect 36499 22214 36557 22220
rect 36976 22211 36982 22223
rect 37034 22211 37040 22263
rect 8272 22063 8278 22115
rect 8330 22063 8336 22115
rect 1152 22004 58848 22026
rect 1152 21952 19654 22004
rect 19706 21952 19718 22004
rect 19770 21952 19782 22004
rect 19834 21952 19846 22004
rect 19898 21952 50374 22004
rect 50426 21952 50438 22004
rect 50490 21952 50502 22004
rect 50554 21952 50566 22004
rect 50618 21952 58848 22004
rect 1152 21930 58848 21952
rect 8272 21841 8278 21893
rect 8330 21881 8336 21893
rect 14704 21881 14710 21893
rect 8330 21853 14710 21881
rect 8330 21841 8336 21853
rect 14704 21841 14710 21853
rect 14762 21841 14768 21893
rect 20563 21736 20621 21742
rect 20563 21702 20575 21736
rect 20609 21733 20621 21736
rect 20851 21736 20909 21742
rect 20851 21733 20863 21736
rect 20609 21705 20863 21733
rect 20609 21702 20621 21705
rect 20563 21696 20621 21702
rect 20851 21702 20863 21705
rect 20897 21733 20909 21736
rect 22864 21733 22870 21745
rect 20897 21705 22870 21733
rect 20897 21702 20909 21705
rect 20851 21696 20909 21702
rect 22864 21693 22870 21705
rect 22922 21693 22928 21745
rect 8272 21545 8278 21597
rect 8330 21585 8336 21597
rect 43888 21585 43894 21597
rect 8330 21557 43894 21585
rect 8330 21545 8336 21557
rect 43888 21545 43894 21557
rect 43946 21545 43952 21597
rect 9811 21440 9869 21446
rect 9811 21406 9823 21440
rect 9857 21437 9869 21440
rect 10000 21437 10006 21449
rect 9857 21409 10006 21437
rect 9857 21406 9869 21409
rect 9811 21400 9869 21406
rect 10000 21397 10006 21409
rect 10058 21397 10064 21449
rect 1152 21338 58848 21360
rect 1152 21286 4294 21338
rect 4346 21286 4358 21338
rect 4410 21286 4422 21338
rect 4474 21286 4486 21338
rect 4538 21286 35014 21338
rect 35066 21286 35078 21338
rect 35130 21286 35142 21338
rect 35194 21286 35206 21338
rect 35258 21286 58848 21338
rect 1152 21264 58848 21286
rect 7603 21218 7661 21224
rect 7603 21184 7615 21218
rect 7649 21215 7661 21218
rect 7891 21218 7949 21224
rect 7891 21215 7903 21218
rect 7649 21187 7903 21215
rect 7649 21184 7661 21187
rect 7603 21178 7661 21184
rect 7891 21184 7903 21187
rect 7937 21184 7949 21218
rect 7891 21178 7949 21184
rect 8179 21218 8237 21224
rect 8179 21184 8191 21218
rect 8225 21215 8237 21218
rect 8225 21187 8558 21215
rect 8225 21184 8237 21187
rect 8179 21178 8237 21184
rect 8194 21127 8222 21178
rect 8530 21141 8558 21187
rect 57712 21141 57718 21153
rect 8530 21113 57718 21141
rect 57712 21101 57718 21113
rect 57770 21101 57776 21153
rect 8230 21005 8282 21011
rect 8230 20947 8282 20953
rect 15568 20879 15574 20931
rect 15626 20919 15632 20931
rect 15763 20922 15821 20928
rect 15763 20919 15775 20922
rect 15626 20891 15775 20919
rect 15626 20879 15632 20891
rect 15763 20888 15775 20891
rect 15809 20888 15821 20922
rect 15763 20882 15821 20888
rect 28243 20922 28301 20928
rect 28243 20888 28255 20922
rect 28289 20919 28301 20922
rect 28336 20919 28342 20931
rect 28289 20891 28342 20919
rect 28289 20888 28301 20891
rect 28243 20882 28301 20888
rect 28336 20879 28342 20891
rect 28394 20879 28400 20931
rect 10768 20845 10774 20857
rect 7954 20771 7982 20831
rect 8544 20817 10774 20845
rect 10768 20805 10774 20817
rect 10826 20805 10832 20857
rect 8272 20771 8278 20783
rect 7954 20743 8278 20771
rect 8272 20731 8278 20743
rect 8330 20731 8336 20783
rect 9328 20731 9334 20783
rect 9386 20771 9392 20783
rect 16624 20771 16630 20783
rect 9386 20743 16630 20771
rect 9386 20731 9392 20743
rect 16624 20731 16630 20743
rect 16682 20731 16688 20783
rect 1152 20672 58848 20694
rect 1152 20620 19654 20672
rect 19706 20620 19718 20672
rect 19770 20620 19782 20672
rect 19834 20620 19846 20672
rect 19898 20620 50374 20672
rect 50426 20620 50438 20672
rect 50490 20620 50502 20672
rect 50554 20620 50566 20672
rect 50618 20620 58848 20672
rect 1152 20598 58848 20620
rect 8272 20509 8278 20561
rect 8330 20549 8336 20561
rect 9328 20549 9334 20561
rect 8330 20521 9334 20549
rect 8330 20509 8336 20521
rect 9328 20509 9334 20521
rect 9386 20509 9392 20561
rect 10768 20509 10774 20561
rect 10826 20549 10832 20561
rect 53968 20549 53974 20561
rect 10826 20521 53974 20549
rect 10826 20509 10832 20521
rect 53968 20509 53974 20521
rect 54026 20509 54032 20561
rect 30928 20435 30934 20487
rect 30986 20475 30992 20487
rect 37939 20478 37997 20484
rect 37939 20475 37951 20478
rect 30986 20447 37951 20475
rect 30986 20435 30992 20447
rect 37939 20444 37951 20447
rect 37985 20444 37997 20478
rect 37939 20438 37997 20444
rect 27088 20105 27094 20117
rect 27049 20077 27094 20105
rect 27088 20065 27094 20077
rect 27146 20065 27152 20117
rect 53008 20105 53014 20117
rect 52969 20077 53014 20105
rect 53008 20065 53014 20077
rect 53066 20065 53072 20117
rect 1152 20006 58848 20028
rect 1152 19954 4294 20006
rect 4346 19954 4358 20006
rect 4410 19954 4422 20006
rect 4474 19954 4486 20006
rect 4538 19954 35014 20006
rect 35066 19954 35078 20006
rect 35130 19954 35142 20006
rect 35194 19954 35206 20006
rect 35258 19954 58848 20006
rect 1152 19932 58848 19954
rect 7603 19886 7661 19892
rect 7603 19852 7615 19886
rect 7649 19883 7661 19886
rect 7891 19886 7949 19892
rect 7891 19883 7903 19886
rect 7649 19855 7903 19883
rect 7649 19852 7661 19855
rect 7603 19846 7661 19852
rect 7891 19852 7903 19855
rect 7937 19852 7949 19886
rect 7891 19846 7949 19852
rect 8179 19886 8237 19892
rect 8179 19852 8191 19886
rect 8225 19883 8237 19886
rect 8225 19855 17294 19883
rect 8225 19852 8237 19855
rect 8179 19846 8237 19852
rect 8194 19795 8222 19846
rect 17266 19809 17294 19855
rect 53680 19809 53686 19821
rect 17266 19781 53686 19809
rect 53680 19769 53686 19781
rect 53738 19769 53744 19821
rect 27184 19547 27190 19599
rect 27242 19587 27248 19599
rect 44083 19590 44141 19596
rect 44083 19587 44095 19590
rect 27242 19559 44095 19587
rect 27242 19547 27248 19559
rect 44083 19556 44095 19559
rect 44129 19556 44141 19590
rect 44083 19550 44141 19556
rect 8080 19513 8086 19525
rect 7968 19485 8086 19513
rect 8080 19473 8086 19485
rect 8138 19473 8144 19525
rect 16528 19513 16534 19525
rect 8256 19485 16534 19513
rect 16528 19473 16534 19485
rect 16586 19473 16592 19525
rect 1152 19340 58848 19362
rect 1152 19288 19654 19340
rect 19706 19288 19718 19340
rect 19770 19288 19782 19340
rect 19834 19288 19846 19340
rect 19898 19288 50374 19340
rect 50426 19288 50438 19340
rect 50490 19288 50502 19340
rect 50554 19288 50566 19340
rect 50618 19288 58848 19340
rect 1152 19266 58848 19288
rect 8080 19177 8086 19229
rect 8138 19217 8144 19229
rect 50800 19217 50806 19229
rect 8138 19189 50806 19217
rect 8138 19177 8144 19189
rect 50800 19177 50806 19189
rect 50858 19177 50864 19229
rect 7024 18881 7030 18933
rect 7082 18921 7088 18933
rect 7792 18921 7798 18933
rect 7082 18893 7798 18921
rect 7082 18881 7088 18893
rect 7792 18881 7798 18893
rect 7850 18881 7856 18933
rect 7504 18733 7510 18785
rect 7562 18773 7568 18785
rect 7792 18773 7798 18785
rect 7562 18745 7798 18773
rect 7562 18733 7568 18745
rect 7792 18733 7798 18745
rect 7850 18733 7856 18785
rect 8371 18776 8429 18782
rect 8371 18742 8383 18776
rect 8417 18773 8429 18776
rect 22960 18773 22966 18785
rect 8417 18745 22966 18773
rect 8417 18742 8429 18745
rect 8371 18736 8429 18742
rect 22960 18733 22966 18745
rect 23018 18733 23024 18785
rect 1152 18674 58848 18696
rect 1152 18622 4294 18674
rect 4346 18622 4358 18674
rect 4410 18622 4422 18674
rect 4474 18622 4486 18674
rect 4538 18622 35014 18674
rect 35066 18622 35078 18674
rect 35130 18622 35142 18674
rect 35194 18622 35206 18674
rect 35258 18622 58848 18674
rect 1152 18600 58848 18622
rect 7603 18554 7661 18560
rect 7603 18520 7615 18554
rect 7649 18551 7661 18554
rect 7649 18523 7982 18551
rect 7649 18520 7661 18523
rect 7603 18514 7661 18520
rect 7954 18477 7982 18523
rect 8656 18511 8662 18563
rect 8714 18551 8720 18563
rect 9331 18554 9389 18560
rect 8714 18523 9134 18551
rect 8714 18511 8720 18523
rect 8275 18480 8333 18486
rect 8275 18477 8287 18480
rect 7954 18449 8287 18477
rect 8275 18446 8287 18449
rect 8321 18446 8333 18480
rect 8275 18440 8333 18446
rect 8467 18480 8525 18486
rect 8467 18446 8479 18480
rect 8513 18477 8525 18480
rect 8947 18480 9005 18486
rect 8947 18477 8959 18480
rect 8513 18449 8959 18477
rect 8513 18446 8525 18449
rect 8467 18440 8525 18446
rect 8947 18446 8959 18449
rect 8993 18446 9005 18480
rect 9106 18477 9134 18523
rect 9331 18520 9343 18554
rect 9377 18551 9389 18554
rect 9377 18523 17294 18551
rect 9377 18520 9389 18523
rect 9331 18514 9389 18520
rect 9106 18449 12974 18477
rect 8947 18440 9005 18446
rect 8230 18287 8282 18293
rect 8230 18229 8282 18235
rect 12946 18255 12974 18449
rect 17266 18403 17294 18523
rect 24403 18480 24461 18486
rect 24403 18446 24415 18480
rect 24449 18477 24461 18480
rect 24691 18480 24749 18486
rect 24691 18477 24703 18480
rect 24449 18449 24703 18477
rect 24449 18446 24461 18449
rect 24403 18440 24461 18446
rect 24691 18446 24703 18449
rect 24737 18477 24749 18480
rect 34384 18477 34390 18489
rect 24737 18449 34390 18477
rect 24737 18446 24749 18449
rect 24691 18440 24749 18446
rect 34384 18437 34390 18449
rect 34442 18437 34448 18489
rect 17266 18375 24926 18403
rect 20656 18329 20662 18341
rect 20617 18301 20662 18329
rect 20656 18289 20662 18301
rect 20714 18289 20720 18341
rect 24898 18329 24926 18375
rect 48880 18329 48886 18341
rect 24898 18301 48886 18329
rect 48880 18289 48886 18301
rect 48938 18289 48944 18341
rect 46096 18255 46102 18267
rect 12946 18227 46102 18255
rect 46096 18215 46102 18227
rect 46154 18215 46160 18267
rect 50128 18215 50134 18267
rect 50186 18255 50192 18267
rect 51667 18258 51725 18264
rect 51667 18255 51679 18258
rect 50186 18227 51679 18255
rect 50186 18215 50192 18227
rect 51667 18224 51679 18227
rect 51713 18224 51725 18258
rect 51667 18218 51725 18224
rect 44752 18181 44758 18193
rect 9120 18153 44758 18181
rect 44752 18141 44758 18153
rect 44810 18141 44816 18193
rect 7120 18067 7126 18119
rect 7178 18107 7184 18119
rect 7312 18107 7318 18119
rect 7178 18079 7318 18107
rect 7178 18067 7184 18079
rect 7312 18067 7318 18079
rect 7370 18067 7376 18119
rect 8656 18067 8662 18119
rect 8714 18067 8720 18119
rect 1152 18008 58848 18030
rect 1152 17956 19654 18008
rect 19706 17956 19718 18008
rect 19770 17956 19782 18008
rect 19834 17956 19846 18008
rect 19898 17956 50374 18008
rect 50426 17956 50438 18008
rect 50490 17956 50502 18008
rect 50554 17956 50566 18008
rect 50618 17956 58848 18008
rect 1152 17934 58848 17956
rect 8656 17845 8662 17897
rect 8714 17885 8720 17897
rect 9040 17885 9046 17897
rect 8714 17857 9046 17885
rect 8714 17845 8720 17857
rect 9040 17845 9046 17857
rect 9098 17845 9104 17897
rect 8176 17771 8182 17823
rect 8234 17811 8240 17823
rect 42928 17811 42934 17823
rect 8234 17783 42934 17811
rect 8234 17771 8240 17783
rect 42928 17771 42934 17783
rect 42986 17771 42992 17823
rect 1747 17444 1805 17450
rect 1747 17410 1759 17444
rect 1793 17441 1805 17444
rect 48880 17441 48886 17453
rect 1793 17413 48886 17441
rect 1793 17410 1805 17413
rect 1747 17404 1805 17410
rect 48880 17401 48886 17413
rect 48938 17401 48944 17453
rect 1152 17342 58848 17364
rect 1152 17290 4294 17342
rect 4346 17290 4358 17342
rect 4410 17290 4422 17342
rect 4474 17290 4486 17342
rect 4538 17290 35014 17342
rect 35066 17290 35078 17342
rect 35130 17290 35142 17342
rect 35194 17290 35206 17342
rect 35258 17290 58848 17342
rect 1152 17268 58848 17290
rect 7408 17179 7414 17231
rect 7466 17219 7472 17231
rect 7507 17222 7565 17228
rect 7507 17219 7519 17222
rect 7466 17191 7519 17219
rect 7466 17179 7472 17191
rect 7507 17188 7519 17191
rect 7553 17188 7565 17222
rect 9040 17219 9046 17231
rect 7507 17182 7565 17188
rect 8770 17191 9046 17219
rect 8770 17131 8798 17191
rect 9040 17179 9046 17191
rect 9098 17219 9104 17231
rect 42640 17219 42646 17231
rect 9098 17191 42646 17219
rect 9098 17179 9104 17191
rect 42640 17179 42646 17191
rect 42698 17179 42704 17231
rect 9043 17074 9101 17080
rect 9043 17040 9055 17074
rect 9089 17071 9101 17074
rect 39760 17071 39766 17083
rect 9089 17043 39766 17071
rect 9089 17040 9101 17043
rect 8674 16932 8702 17036
rect 9043 17034 9101 17040
rect 39760 17031 39766 17043
rect 39818 17031 39824 17083
rect 8659 16926 8717 16932
rect 8659 16892 8671 16926
rect 8705 16892 8717 16926
rect 8659 16886 8717 16892
rect 24496 16883 24502 16935
rect 24554 16923 24560 16935
rect 30451 16926 30509 16932
rect 30451 16923 30463 16926
rect 24554 16895 30463 16923
rect 24554 16883 24560 16895
rect 30451 16892 30463 16895
rect 30497 16892 30509 16926
rect 30451 16886 30509 16892
rect 1152 16676 58848 16698
rect 1152 16624 19654 16676
rect 19706 16624 19718 16676
rect 19770 16624 19782 16676
rect 19834 16624 19846 16676
rect 19898 16624 50374 16676
rect 50426 16624 50438 16676
rect 50490 16624 50502 16676
rect 50554 16624 50566 16676
rect 50618 16624 58848 16676
rect 1152 16602 58848 16624
rect 7408 16069 7414 16121
rect 7466 16109 7472 16121
rect 8176 16109 8182 16121
rect 7466 16081 8182 16109
rect 7466 16069 7472 16081
rect 8176 16069 8182 16081
rect 8234 16069 8240 16121
rect 1152 16010 58848 16032
rect 1152 15958 4294 16010
rect 4346 15958 4358 16010
rect 4410 15958 4422 16010
rect 4474 15958 4486 16010
rect 4538 15958 35014 16010
rect 35066 15958 35078 16010
rect 35130 15958 35142 16010
rect 35194 15958 35206 16010
rect 35258 15958 58848 16010
rect 1152 15936 58848 15958
rect 7408 15847 7414 15899
rect 7466 15887 7472 15899
rect 7507 15890 7565 15896
rect 7507 15887 7519 15890
rect 7466 15859 7519 15887
rect 7466 15847 7472 15859
rect 7507 15856 7519 15859
rect 7553 15856 7565 15890
rect 7507 15850 7565 15856
rect 8176 15847 8182 15899
rect 8234 15887 8240 15899
rect 8234 15859 10094 15887
rect 8234 15847 8240 15859
rect 8194 15799 8222 15847
rect 10066 15813 10094 15859
rect 20368 15847 20374 15899
rect 20426 15887 20432 15899
rect 55315 15890 55373 15896
rect 55315 15887 55327 15890
rect 20426 15859 55327 15887
rect 20426 15847 20432 15859
rect 55315 15856 55327 15859
rect 55361 15887 55373 15890
rect 55507 15890 55565 15896
rect 55507 15887 55519 15890
rect 55361 15859 55519 15887
rect 55361 15856 55373 15859
rect 55315 15850 55373 15856
rect 55507 15856 55519 15859
rect 55553 15856 55565 15890
rect 55507 15850 55565 15856
rect 38896 15813 38902 15825
rect 10066 15785 38902 15813
rect 38896 15773 38902 15785
rect 38954 15773 38960 15825
rect 19219 15594 19277 15600
rect 19219 15560 19231 15594
rect 19265 15591 19277 15594
rect 19507 15594 19565 15600
rect 19507 15591 19519 15594
rect 19265 15563 19519 15591
rect 19265 15560 19277 15563
rect 19219 15554 19277 15560
rect 19507 15560 19519 15563
rect 19553 15591 19565 15594
rect 27664 15591 27670 15603
rect 19553 15563 27670 15591
rect 19553 15560 19565 15563
rect 19507 15554 19565 15560
rect 27664 15551 27670 15563
rect 27722 15551 27728 15603
rect 8176 15477 8182 15529
rect 8234 15477 8240 15529
rect 1152 15344 58848 15366
rect 1152 15292 19654 15344
rect 19706 15292 19718 15344
rect 19770 15292 19782 15344
rect 19834 15292 19846 15344
rect 19898 15292 50374 15344
rect 50426 15292 50438 15344
rect 50490 15292 50502 15344
rect 50554 15292 50566 15344
rect 50618 15292 58848 15344
rect 1152 15270 58848 15292
rect 8176 15181 8182 15233
rect 8234 15221 8240 15233
rect 36688 15221 36694 15233
rect 8234 15193 36694 15221
rect 8234 15181 8240 15193
rect 36688 15181 36694 15193
rect 36746 15181 36752 15233
rect 7888 15107 7894 15159
rect 7946 15147 7952 15159
rect 8272 15147 8278 15159
rect 7946 15119 8278 15147
rect 7946 15107 7952 15119
rect 8272 15107 8278 15119
rect 8330 15107 8336 15159
rect 15091 14854 15149 14860
rect 15091 14820 15103 14854
rect 15137 14851 15149 14854
rect 18448 14851 18454 14863
rect 15137 14823 18454 14851
rect 15137 14820 15149 14823
rect 15091 14814 15149 14820
rect 18448 14811 18454 14823
rect 18506 14811 18512 14863
rect 18259 14780 18317 14786
rect 18259 14746 18271 14780
rect 18305 14777 18317 14780
rect 24688 14777 24694 14789
rect 18305 14749 24694 14777
rect 18305 14746 18317 14749
rect 18259 14740 18317 14746
rect 24688 14737 24694 14749
rect 24746 14737 24752 14789
rect 1152 14678 58848 14700
rect 1152 14626 4294 14678
rect 4346 14626 4358 14678
rect 4410 14626 4422 14678
rect 4474 14626 4486 14678
rect 4538 14626 35014 14678
rect 35066 14626 35078 14678
rect 35130 14626 35142 14678
rect 35194 14626 35206 14678
rect 35258 14626 58848 14678
rect 1152 14604 58848 14626
rect 44371 14484 44429 14490
rect 44371 14450 44383 14484
rect 44417 14481 44429 14484
rect 53392 14481 53398 14493
rect 44417 14453 53398 14481
rect 44417 14450 44429 14453
rect 44371 14444 44429 14450
rect 53392 14441 53398 14453
rect 53450 14441 53456 14493
rect 51184 14259 51190 14271
rect 51145 14231 51190 14259
rect 51184 14219 51190 14231
rect 51242 14219 51248 14271
rect 25552 14185 25558 14197
rect 7968 14157 25558 14185
rect 25552 14145 25558 14157
rect 25610 14145 25616 14197
rect 7603 14114 7661 14120
rect 7603 14080 7615 14114
rect 7649 14111 7661 14114
rect 36592 14111 36598 14123
rect 7649 14083 36598 14111
rect 7649 14080 7661 14083
rect 7603 14074 7661 14080
rect 36592 14071 36598 14083
rect 36650 14071 36656 14123
rect 1152 14012 58848 14034
rect 1152 13960 19654 14012
rect 19706 13960 19718 14012
rect 19770 13960 19782 14012
rect 19834 13960 19846 14012
rect 19898 13960 50374 14012
rect 50426 13960 50438 14012
rect 50490 13960 50502 14012
rect 50554 13960 50566 14012
rect 50618 13960 58848 14012
rect 1152 13938 58848 13960
rect 15952 13889 15958 13901
rect 15913 13861 15958 13889
rect 15952 13849 15958 13861
rect 16010 13889 16016 13901
rect 16010 13861 16286 13889
rect 16010 13849 16016 13861
rect 16258 13750 16286 13861
rect 16243 13744 16301 13750
rect 16243 13710 16255 13744
rect 16289 13710 16301 13744
rect 16243 13704 16301 13710
rect 3280 13405 3286 13457
rect 3338 13445 3344 13457
rect 8176 13445 8182 13457
rect 3338 13417 8182 13445
rect 3338 13405 3344 13417
rect 8176 13405 8182 13417
rect 8234 13405 8240 13457
rect 11440 13445 11446 13457
rect 11401 13417 11446 13445
rect 11440 13405 11446 13417
rect 11498 13405 11504 13457
rect 45136 13445 45142 13457
rect 45097 13417 45142 13445
rect 45136 13405 45142 13417
rect 45194 13405 45200 13457
rect 1152 13346 58848 13368
rect 1152 13294 4294 13346
rect 4346 13294 4358 13346
rect 4410 13294 4422 13346
rect 4474 13294 4486 13346
rect 4538 13294 35014 13346
rect 35066 13294 35078 13346
rect 35130 13294 35142 13346
rect 35194 13294 35206 13346
rect 35258 13294 58848 13346
rect 1152 13272 58848 13294
rect 7504 13183 7510 13235
rect 7562 13183 7568 13235
rect 8176 13183 8182 13235
rect 8234 13223 8240 13235
rect 45136 13223 45142 13235
rect 8234 13195 45142 13223
rect 8234 13183 8240 13195
rect 45136 13183 45142 13195
rect 45194 13183 45200 13235
rect 56851 13226 56909 13232
rect 56851 13192 56863 13226
rect 56897 13223 56909 13226
rect 56944 13223 56950 13235
rect 56897 13195 56950 13223
rect 56897 13192 56909 13195
rect 56851 13186 56909 13192
rect 56944 13183 56950 13195
rect 57002 13183 57008 13235
rect 7216 12961 7222 13013
rect 7274 13001 7280 13013
rect 7522 13001 7550 13183
rect 7603 13152 7661 13158
rect 7603 13118 7615 13152
rect 7649 13149 7661 13152
rect 33040 13149 33046 13161
rect 7649 13121 33046 13149
rect 7649 13118 7661 13121
rect 7603 13112 7661 13118
rect 33040 13109 33046 13121
rect 33098 13109 33104 13161
rect 56962 13084 56990 13183
rect 56947 13078 57005 13084
rect 56947 13044 56959 13078
rect 56993 13044 57005 13078
rect 56947 13038 57005 13044
rect 7274 12973 7550 13001
rect 7274 12961 7280 12973
rect 56272 12961 56278 13013
rect 56330 13001 56336 13013
rect 57811 13004 57869 13010
rect 57811 13001 57823 13004
rect 56330 12973 57823 13001
rect 56330 12961 56336 12973
rect 57811 12970 57823 12973
rect 57857 12970 57869 13004
rect 57811 12964 57869 12970
rect 30064 12853 30070 12865
rect 7968 12825 30070 12853
rect 30064 12813 30070 12825
rect 30122 12813 30128 12865
rect 1152 12680 58848 12702
rect 1152 12628 19654 12680
rect 19706 12628 19718 12680
rect 19770 12628 19782 12680
rect 19834 12628 19846 12680
rect 19898 12628 50374 12680
rect 50426 12628 50438 12680
rect 50490 12628 50502 12680
rect 50554 12628 50566 12680
rect 50618 12628 58848 12680
rect 1152 12606 58848 12628
rect 7600 12517 7606 12569
rect 7658 12557 7664 12569
rect 7792 12557 7798 12569
rect 7658 12529 7798 12557
rect 7658 12517 7664 12529
rect 7792 12517 7798 12529
rect 7850 12517 7856 12569
rect 57328 12557 57334 12569
rect 57289 12529 57334 12557
rect 57328 12517 57334 12529
rect 57386 12517 57392 12569
rect 57346 12409 57374 12517
rect 57619 12412 57677 12418
rect 57619 12409 57631 12412
rect 57346 12381 57631 12409
rect 57619 12378 57631 12381
rect 57665 12409 57677 12412
rect 57907 12412 57965 12418
rect 57907 12409 57919 12412
rect 57665 12381 57919 12409
rect 57665 12378 57677 12381
rect 57619 12372 57677 12378
rect 57907 12378 57919 12381
rect 57953 12378 57965 12412
rect 57907 12372 57965 12378
rect 10000 12295 10006 12347
rect 10058 12335 10064 12347
rect 17968 12335 17974 12347
rect 10058 12307 17974 12335
rect 10058 12295 10064 12307
rect 17968 12295 17974 12307
rect 18026 12295 18032 12347
rect 37459 12264 37517 12270
rect 37459 12230 37471 12264
rect 37505 12261 37517 12264
rect 37747 12264 37805 12270
rect 37747 12261 37759 12264
rect 37505 12233 37759 12261
rect 37505 12230 37517 12233
rect 37459 12224 37517 12230
rect 37747 12230 37759 12233
rect 37793 12261 37805 12264
rect 57424 12261 57430 12273
rect 37793 12233 57430 12261
rect 37793 12230 37805 12233
rect 37747 12224 37805 12230
rect 57424 12221 57430 12233
rect 57482 12221 57488 12273
rect 57715 12264 57773 12270
rect 57715 12230 57727 12264
rect 57761 12230 57773 12264
rect 57715 12224 57773 12230
rect 2131 12190 2189 12196
rect 2131 12156 2143 12190
rect 2177 12187 2189 12190
rect 10000 12187 10006 12199
rect 2177 12159 10006 12187
rect 2177 12156 2189 12159
rect 2131 12150 2189 12156
rect 10000 12147 10006 12159
rect 10058 12147 10064 12199
rect 48979 12190 49037 12196
rect 48979 12187 48991 12190
rect 23026 12159 48991 12187
rect 6544 12113 6550 12125
rect 6505 12085 6550 12113
rect 6544 12073 6550 12085
rect 6602 12073 6608 12125
rect 13648 12073 13654 12125
rect 13706 12113 13712 12125
rect 23026 12113 23054 12159
rect 48979 12156 48991 12159
rect 49025 12187 49037 12190
rect 49171 12190 49229 12196
rect 49171 12187 49183 12190
rect 49025 12159 49183 12187
rect 49025 12156 49037 12159
rect 48979 12150 49037 12156
rect 49171 12156 49183 12159
rect 49217 12156 49229 12190
rect 49171 12150 49229 12156
rect 57520 12147 57526 12199
rect 57578 12187 57584 12199
rect 57730 12187 57758 12224
rect 57578 12159 57758 12187
rect 57578 12147 57584 12159
rect 13706 12085 23054 12113
rect 13706 12073 13712 12085
rect 1152 12014 58848 12036
rect 1152 11962 4294 12014
rect 4346 11962 4358 12014
rect 4410 11962 4422 12014
rect 4474 11962 4486 12014
rect 4538 11962 35014 12014
rect 35066 11962 35078 12014
rect 35130 11962 35142 12014
rect 35194 11962 35206 12014
rect 35258 11962 58848 12014
rect 1152 11940 58848 11962
rect 7024 11851 7030 11903
rect 7082 11891 7088 11903
rect 7312 11891 7318 11903
rect 7082 11863 7318 11891
rect 7082 11851 7088 11863
rect 7312 11851 7318 11863
rect 7370 11851 7376 11903
rect 7603 11820 7661 11826
rect 7603 11786 7615 11820
rect 7649 11817 7661 11820
rect 29296 11817 29302 11829
rect 7649 11789 29302 11817
rect 7649 11786 7661 11789
rect 7603 11780 7661 11786
rect 29296 11777 29302 11789
rect 29354 11777 29360 11829
rect 56851 11820 56909 11826
rect 56851 11817 56863 11820
rect 43186 11789 56863 11817
rect 7968 11715 12974 11743
rect 12946 11669 12974 11715
rect 17968 11703 17974 11755
rect 18026 11743 18032 11755
rect 43186 11743 43214 11789
rect 56851 11786 56863 11789
rect 56897 11817 56909 11820
rect 56947 11820 57005 11826
rect 56947 11817 56959 11820
rect 56897 11789 56959 11817
rect 56897 11786 56909 11789
rect 56851 11780 56909 11786
rect 56947 11786 56959 11789
rect 56993 11786 57005 11820
rect 56947 11780 57005 11786
rect 18026 11715 43214 11743
rect 56563 11746 56621 11752
rect 18026 11703 18032 11715
rect 56563 11712 56575 11746
rect 56609 11743 56621 11746
rect 56609 11715 57614 11743
rect 56609 11712 56621 11715
rect 56563 11706 56621 11712
rect 25168 11669 25174 11681
rect 12946 11641 25174 11669
rect 25168 11629 25174 11641
rect 25226 11629 25232 11681
rect 27088 11629 27094 11681
rect 27146 11669 27152 11681
rect 56179 11672 56237 11678
rect 56179 11669 56191 11672
rect 27146 11641 56191 11669
rect 27146 11629 27152 11641
rect 56179 11638 56191 11641
rect 56225 11669 56237 11672
rect 56467 11672 56525 11678
rect 56467 11669 56479 11672
rect 56225 11641 56479 11669
rect 56225 11638 56237 11641
rect 56179 11632 56237 11638
rect 56467 11638 56479 11641
rect 56513 11638 56525 11672
rect 56467 11632 56525 11638
rect 56851 11672 56909 11678
rect 56851 11638 56863 11672
rect 56897 11669 56909 11672
rect 57235 11672 57293 11678
rect 57235 11669 57247 11672
rect 56897 11641 57247 11669
rect 56897 11638 56909 11641
rect 56851 11632 56909 11638
rect 57235 11638 57247 11641
rect 57281 11638 57293 11672
rect 57235 11632 57293 11638
rect 23923 11598 23981 11604
rect 23923 11564 23935 11598
rect 23969 11595 23981 11598
rect 24400 11595 24406 11607
rect 23969 11567 24406 11595
rect 23969 11564 23981 11567
rect 23923 11558 23981 11564
rect 24400 11555 24406 11567
rect 24458 11555 24464 11607
rect 54736 11555 54742 11607
rect 54794 11595 54800 11607
rect 55891 11598 55949 11604
rect 55891 11595 55903 11598
rect 54794 11567 55903 11595
rect 54794 11555 54800 11567
rect 55891 11564 55903 11567
rect 55937 11564 55949 11598
rect 57586 11595 57614 11715
rect 58192 11595 58198 11607
rect 57586 11567 58198 11595
rect 55891 11558 55949 11564
rect 58192 11555 58198 11567
rect 58250 11555 58256 11607
rect 57136 11407 57142 11459
rect 57194 11447 57200 11459
rect 57331 11450 57389 11456
rect 57331 11447 57343 11450
rect 57194 11419 57343 11447
rect 57194 11407 57200 11419
rect 57331 11416 57343 11419
rect 57377 11416 57389 11450
rect 57331 11410 57389 11416
rect 1152 11348 58848 11370
rect 1152 11296 19654 11348
rect 19706 11296 19718 11348
rect 19770 11296 19782 11348
rect 19834 11296 19846 11348
rect 19898 11296 50374 11348
rect 50426 11296 50438 11348
rect 50490 11296 50502 11348
rect 50554 11296 50566 11348
rect 50618 11296 58848 11348
rect 1152 11274 58848 11296
rect 7792 11185 7798 11237
rect 7850 11225 7856 11237
rect 8080 11225 8086 11237
rect 7850 11197 8086 11225
rect 7850 11185 7856 11197
rect 8080 11185 8086 11197
rect 8138 11185 8144 11237
rect 8080 11037 8086 11089
rect 8138 11077 8144 11089
rect 22288 11077 22294 11089
rect 8138 11049 22294 11077
rect 8138 11037 8144 11049
rect 22288 11037 22294 11049
rect 22346 11037 22352 11089
rect 28144 11037 28150 11089
rect 28202 11077 28208 11089
rect 37939 11080 37997 11086
rect 37939 11077 37951 11080
rect 28202 11049 37951 11077
rect 28202 11037 28208 11049
rect 37939 11046 37951 11049
rect 37985 11046 37997 11080
rect 56947 11080 57005 11086
rect 56947 11077 56959 11080
rect 37939 11040 37997 11046
rect 43186 11049 56959 11077
rect 17776 10963 17782 11015
rect 17834 11003 17840 11015
rect 43186 11003 43214 11049
rect 56947 11046 56959 11049
rect 56993 11077 57005 11080
rect 57235 11080 57293 11086
rect 57235 11077 57247 11080
rect 56993 11049 57247 11077
rect 56993 11046 57005 11049
rect 56947 11040 57005 11046
rect 57235 11046 57247 11049
rect 57281 11046 57293 11080
rect 57235 11040 57293 11046
rect 56083 11006 56141 11012
rect 56083 11003 56095 11006
rect 17834 10975 43214 11003
rect 53266 10975 56095 11003
rect 17834 10963 17840 10975
rect 9616 10889 9622 10941
rect 9674 10929 9680 10941
rect 26512 10929 26518 10941
rect 9674 10901 26518 10929
rect 9674 10889 9680 10901
rect 26512 10889 26518 10901
rect 26570 10889 26576 10941
rect 29776 10889 29782 10941
rect 29834 10929 29840 10941
rect 53266 10929 53294 10975
rect 56083 10972 56095 10975
rect 56129 10972 56141 11006
rect 56083 10966 56141 10972
rect 29834 10901 53294 10929
rect 55987 10932 56045 10938
rect 29834 10889 29840 10901
rect 55987 10898 55999 10932
rect 56033 10929 56045 10932
rect 56752 10929 56758 10941
rect 56033 10901 56758 10929
rect 56033 10898 56045 10901
rect 55987 10892 56045 10898
rect 56752 10889 56758 10901
rect 56810 10889 56816 10941
rect 57331 10932 57389 10938
rect 57331 10898 57343 10932
rect 57377 10898 57389 10932
rect 57331 10892 57389 10898
rect 4720 10815 4726 10867
rect 4778 10855 4784 10867
rect 18835 10858 18893 10864
rect 18835 10855 18847 10858
rect 4778 10827 18847 10855
rect 4778 10815 4784 10827
rect 18835 10824 18847 10827
rect 18881 10855 18893 10858
rect 19027 10858 19085 10864
rect 19027 10855 19039 10858
rect 18881 10827 19039 10855
rect 18881 10824 18893 10827
rect 18835 10818 18893 10824
rect 19027 10824 19039 10827
rect 19073 10824 19085 10858
rect 19027 10818 19085 10824
rect 29395 10858 29453 10864
rect 29395 10824 29407 10858
rect 29441 10855 29453 10858
rect 34288 10855 34294 10867
rect 29441 10827 34294 10855
rect 29441 10824 29453 10827
rect 29395 10818 29453 10824
rect 34288 10815 34294 10827
rect 34346 10815 34352 10867
rect 37939 10858 37997 10864
rect 37939 10824 37951 10858
rect 37985 10855 37997 10858
rect 48595 10858 48653 10864
rect 48595 10855 48607 10858
rect 37985 10827 48607 10855
rect 37985 10824 37997 10827
rect 37939 10818 37997 10824
rect 48595 10824 48607 10827
rect 48641 10855 48653 10858
rect 48787 10858 48845 10864
rect 48787 10855 48799 10858
rect 48641 10827 48799 10855
rect 48641 10824 48653 10827
rect 48595 10818 48653 10824
rect 48787 10824 48799 10827
rect 48833 10824 48845 10858
rect 48787 10818 48845 10824
rect 56560 10815 56566 10867
rect 56618 10855 56624 10867
rect 57346 10855 57374 10892
rect 56618 10827 57374 10855
rect 56618 10815 56624 10827
rect 7984 10741 7990 10793
rect 8042 10781 8048 10793
rect 8083 10784 8141 10790
rect 8083 10781 8095 10784
rect 8042 10753 8095 10781
rect 8042 10741 8048 10753
rect 8083 10750 8095 10753
rect 8129 10750 8141 10784
rect 8083 10744 8141 10750
rect 9907 10784 9965 10790
rect 9907 10750 9919 10784
rect 9953 10781 9965 10784
rect 11152 10781 11158 10793
rect 9953 10753 11158 10781
rect 9953 10750 9965 10753
rect 9907 10744 9965 10750
rect 11152 10741 11158 10753
rect 11210 10741 11216 10793
rect 31696 10741 31702 10793
rect 31754 10781 31760 10793
rect 32467 10784 32525 10790
rect 32467 10781 32479 10784
rect 31754 10753 32479 10781
rect 31754 10741 31760 10753
rect 32467 10750 32479 10753
rect 32513 10750 32525 10784
rect 32467 10744 32525 10750
rect 48208 10741 48214 10793
rect 48266 10781 48272 10793
rect 54643 10784 54701 10790
rect 54643 10781 54655 10784
rect 48266 10753 54655 10781
rect 48266 10741 48272 10753
rect 54643 10750 54655 10753
rect 54689 10750 54701 10784
rect 54643 10744 54701 10750
rect 1152 10682 58848 10704
rect 1152 10630 4294 10682
rect 4346 10630 4358 10682
rect 4410 10630 4422 10682
rect 4474 10630 4486 10682
rect 4538 10630 35014 10682
rect 35066 10630 35078 10682
rect 35130 10630 35142 10682
rect 35194 10630 35206 10682
rect 35258 10630 58848 10682
rect 1152 10608 58848 10630
rect 7603 10562 7661 10568
rect 7603 10528 7615 10562
rect 7649 10559 7661 10562
rect 7649 10531 7982 10559
rect 7649 10528 7661 10531
rect 7603 10522 7661 10528
rect 7954 10485 7982 10531
rect 8176 10519 8182 10571
rect 8234 10559 8240 10571
rect 8464 10559 8470 10571
rect 8234 10531 8470 10559
rect 8234 10519 8240 10531
rect 8464 10519 8470 10531
rect 8522 10519 8528 10571
rect 33808 10519 33814 10571
rect 33866 10559 33872 10571
rect 48208 10559 48214 10571
rect 33866 10531 48214 10559
rect 33866 10519 33872 10531
rect 48208 10519 48214 10531
rect 48266 10519 48272 10571
rect 56371 10562 56429 10568
rect 56371 10528 56383 10562
rect 56417 10559 56429 10562
rect 56464 10559 56470 10571
rect 56417 10531 56470 10559
rect 56417 10528 56429 10531
rect 56371 10522 56429 10528
rect 56464 10519 56470 10531
rect 56522 10559 56528 10571
rect 56522 10531 56702 10559
rect 56522 10519 56528 10531
rect 9616 10485 9622 10497
rect 7954 10457 9622 10485
rect 9616 10445 9622 10457
rect 9674 10445 9680 10497
rect 8080 10411 8086 10423
rect 7968 10383 8086 10411
rect 8080 10371 8086 10383
rect 8138 10371 8144 10423
rect 55888 10411 55894 10423
rect 55849 10383 55894 10411
rect 55888 10371 55894 10383
rect 55946 10371 55952 10423
rect 56674 10420 56702 10531
rect 56659 10414 56717 10420
rect 56659 10380 56671 10414
rect 56705 10380 56717 10414
rect 56659 10374 56717 10380
rect 11632 10297 11638 10349
rect 11690 10337 11696 10349
rect 54739 10340 54797 10346
rect 54739 10337 54751 10340
rect 11690 10309 54751 10337
rect 11690 10297 11696 10309
rect 54739 10306 54751 10309
rect 54785 10337 54797 10340
rect 55027 10340 55085 10346
rect 55027 10337 55039 10340
rect 54785 10309 55039 10337
rect 54785 10306 54797 10309
rect 54739 10300 54797 10306
rect 55027 10306 55039 10309
rect 55073 10306 55085 10340
rect 55027 10300 55085 10306
rect 55696 10297 55702 10349
rect 55754 10337 55760 10349
rect 57427 10340 57485 10346
rect 57427 10337 57439 10340
rect 55754 10309 57439 10337
rect 55754 10297 55760 10309
rect 57427 10306 57439 10309
rect 57473 10306 57485 10340
rect 57427 10300 57485 10306
rect 9136 10223 9142 10275
rect 9194 10263 9200 10275
rect 9328 10263 9334 10275
rect 9194 10235 9334 10263
rect 9194 10223 9200 10235
rect 9328 10223 9334 10235
rect 9386 10223 9392 10275
rect 39571 10266 39629 10272
rect 39571 10232 39583 10266
rect 39617 10263 39629 10266
rect 41488 10263 41494 10275
rect 39617 10235 41494 10263
rect 39617 10232 39629 10235
rect 39571 10226 39629 10232
rect 41488 10223 41494 10235
rect 41546 10223 41552 10275
rect 56464 10223 56470 10275
rect 56522 10263 56528 10275
rect 57347 10266 57405 10272
rect 57347 10263 57359 10266
rect 56522 10235 57359 10263
rect 56522 10223 56528 10235
rect 57347 10232 57359 10235
rect 57393 10232 57405 10266
rect 57347 10226 57405 10232
rect 58576 10189 58582 10201
rect 55138 10161 58582 10189
rect 8752 10075 8758 10127
rect 8810 10115 8816 10127
rect 9136 10115 9142 10127
rect 8810 10087 9142 10115
rect 8810 10075 8816 10087
rect 9136 10075 9142 10087
rect 9194 10075 9200 10127
rect 55138 10124 55166 10161
rect 58576 10149 58582 10161
rect 58634 10149 58640 10201
rect 55123 10118 55181 10124
rect 55123 10084 55135 10118
rect 55169 10084 55181 10118
rect 55123 10078 55181 10084
rect 55696 10075 55702 10127
rect 55754 10115 55760 10127
rect 55795 10118 55853 10124
rect 55795 10115 55807 10118
rect 55754 10087 55807 10115
rect 55754 10075 55760 10087
rect 55795 10084 55807 10087
rect 55841 10084 55853 10118
rect 55795 10078 55853 10084
rect 56080 10075 56086 10127
rect 56138 10115 56144 10127
rect 56563 10118 56621 10124
rect 56563 10115 56575 10118
rect 56138 10087 56575 10115
rect 56138 10075 56144 10087
rect 56563 10084 56575 10087
rect 56609 10084 56621 10118
rect 56563 10078 56621 10084
rect 1152 10016 58848 10038
rect 1152 9964 19654 10016
rect 19706 9964 19718 10016
rect 19770 9964 19782 10016
rect 19834 9964 19846 10016
rect 19898 9964 50374 10016
rect 50426 9964 50438 10016
rect 50490 9964 50502 10016
rect 50554 9964 50566 10016
rect 50618 9964 58848 10016
rect 1152 9942 58848 9964
rect 7024 9853 7030 9905
rect 7082 9893 7088 9905
rect 8752 9893 8758 9905
rect 7082 9865 8758 9893
rect 7082 9853 7088 9865
rect 8752 9853 8758 9865
rect 8810 9893 8816 9905
rect 23440 9893 23446 9905
rect 8810 9865 23446 9893
rect 8810 9853 8816 9865
rect 23440 9853 23446 9865
rect 23498 9853 23504 9905
rect 54928 9853 54934 9905
rect 54986 9893 54992 9905
rect 55219 9896 55277 9902
rect 55219 9893 55231 9896
rect 54986 9865 55231 9893
rect 54986 9853 54992 9865
rect 55219 9862 55231 9865
rect 55265 9862 55277 9896
rect 55219 9856 55277 9862
rect 55312 9853 55318 9905
rect 55370 9893 55376 9905
rect 55987 9896 56045 9902
rect 55987 9893 55999 9896
rect 55370 9865 55999 9893
rect 55370 9853 55376 9865
rect 55987 9862 55999 9865
rect 56033 9862 56045 9896
rect 55987 9856 56045 9862
rect 7984 9779 7990 9831
rect 8042 9819 8048 9831
rect 9616 9819 9622 9831
rect 8042 9791 9622 9819
rect 8042 9779 8048 9791
rect 9616 9779 9622 9791
rect 9674 9779 9680 9831
rect 41584 9779 41590 9831
rect 41642 9819 41648 9831
rect 49072 9819 49078 9831
rect 41642 9791 49078 9819
rect 41642 9779 41648 9791
rect 49072 9779 49078 9791
rect 49130 9779 49136 9831
rect 55600 9819 55606 9831
rect 55561 9791 55606 9819
rect 55600 9779 55606 9791
rect 55658 9819 55664 9831
rect 56179 9822 56237 9828
rect 56179 9819 56191 9822
rect 55658 9791 56191 9819
rect 55658 9779 55664 9791
rect 8272 9705 8278 9757
rect 8330 9745 8336 9757
rect 16144 9745 16150 9757
rect 8330 9717 16150 9745
rect 8330 9705 8336 9717
rect 16144 9705 16150 9717
rect 16202 9705 16208 9757
rect 41776 9705 41782 9757
rect 41834 9745 41840 9757
rect 49936 9745 49942 9757
rect 41834 9717 49942 9745
rect 41834 9705 41840 9717
rect 49936 9705 49942 9717
rect 49994 9705 50000 9757
rect 55906 9754 55934 9791
rect 56179 9788 56191 9791
rect 56225 9788 56237 9822
rect 56179 9782 56237 9788
rect 55891 9748 55949 9754
rect 55891 9714 55903 9748
rect 55937 9714 55949 9748
rect 55891 9708 55949 9714
rect 3376 9631 3382 9683
rect 3434 9671 3440 9683
rect 39568 9671 39574 9683
rect 3434 9643 39574 9671
rect 3434 9631 3440 9643
rect 39568 9631 39574 9643
rect 39626 9631 39632 9683
rect 54835 9674 54893 9680
rect 54835 9671 54847 9674
rect 43186 9643 54847 9671
rect 8368 9557 8374 9609
rect 8426 9597 8432 9609
rect 8560 9597 8566 9609
rect 8426 9569 8566 9597
rect 8426 9557 8432 9569
rect 8560 9557 8566 9569
rect 8618 9557 8624 9609
rect 28624 9557 28630 9609
rect 28682 9597 28688 9609
rect 43186 9597 43214 9643
rect 54835 9640 54847 9643
rect 54881 9671 54893 9674
rect 55123 9674 55181 9680
rect 55123 9671 55135 9674
rect 54881 9643 55135 9671
rect 54881 9640 54893 9643
rect 54835 9634 54893 9640
rect 55123 9640 55135 9643
rect 55169 9640 55181 9674
rect 55123 9634 55181 9640
rect 57616 9631 57622 9683
rect 57674 9671 57680 9683
rect 57674 9643 57719 9671
rect 57674 9631 57680 9643
rect 28682 9569 43214 9597
rect 28682 9557 28688 9569
rect 54256 9557 54262 9609
rect 54314 9597 54320 9609
rect 54355 9600 54413 9606
rect 54355 9597 54367 9600
rect 54314 9569 54367 9597
rect 54314 9557 54320 9569
rect 54355 9566 54367 9569
rect 54401 9566 54413 9600
rect 54355 9560 54413 9566
rect 54448 9557 54454 9609
rect 54506 9597 54512 9609
rect 54506 9569 54551 9597
rect 54506 9557 54512 9569
rect 8080 9483 8086 9535
rect 8138 9523 8144 9535
rect 17872 9523 17878 9535
rect 8138 9495 17878 9523
rect 8138 9483 8144 9495
rect 17872 9483 17878 9495
rect 17930 9483 17936 9535
rect 24211 9526 24269 9532
rect 24211 9492 24223 9526
rect 24257 9523 24269 9526
rect 24499 9526 24557 9532
rect 24499 9523 24511 9526
rect 24257 9495 24511 9523
rect 24257 9492 24269 9495
rect 24211 9486 24269 9492
rect 24499 9492 24511 9495
rect 24545 9523 24557 9526
rect 57808 9523 57814 9535
rect 24545 9495 57814 9523
rect 24545 9492 24557 9495
rect 24499 9486 24557 9492
rect 57808 9483 57814 9495
rect 57866 9483 57872 9535
rect 8560 9409 8566 9461
rect 8618 9449 8624 9461
rect 19312 9449 19318 9461
rect 8618 9421 19318 9449
rect 8618 9409 8624 9421
rect 19312 9409 19318 9421
rect 19370 9409 19376 9461
rect 47536 9409 47542 9461
rect 47594 9449 47600 9461
rect 50323 9452 50381 9458
rect 50323 9449 50335 9452
rect 47594 9421 50335 9449
rect 47594 9409 47600 9421
rect 50323 9418 50335 9421
rect 50369 9418 50381 9452
rect 52624 9449 52630 9461
rect 52585 9421 52630 9449
rect 50323 9412 50381 9418
rect 52624 9409 52630 9421
rect 52682 9409 52688 9461
rect 1152 9350 58848 9372
rect 1152 9298 4294 9350
rect 4346 9298 4358 9350
rect 4410 9298 4422 9350
rect 4474 9298 4486 9350
rect 4538 9298 35014 9350
rect 35066 9298 35078 9350
rect 35130 9298 35142 9350
rect 35194 9298 35206 9350
rect 35258 9298 58848 9350
rect 1152 9276 58848 9298
rect 7024 9187 7030 9239
rect 7082 9227 7088 9239
rect 7507 9230 7565 9236
rect 7507 9227 7519 9230
rect 7082 9199 7519 9227
rect 7082 9187 7088 9199
rect 7507 9196 7519 9199
rect 7553 9196 7565 9230
rect 7507 9190 7565 9196
rect 8179 9230 8237 9236
rect 8179 9196 8191 9230
rect 8225 9227 8237 9230
rect 8272 9227 8278 9239
rect 8225 9199 8278 9227
rect 8225 9196 8237 9199
rect 8179 9190 8237 9196
rect 8272 9187 8278 9199
rect 8330 9187 8336 9239
rect 20944 9187 20950 9239
rect 21002 9227 21008 9239
rect 52624 9227 52630 9239
rect 21002 9199 52630 9227
rect 21002 9187 21008 9199
rect 52624 9187 52630 9199
rect 52682 9187 52688 9239
rect 8560 9113 8566 9165
rect 8618 9113 8624 9165
rect 8752 9113 8758 9165
rect 8810 9113 8816 9165
rect 39568 9153 39574 9165
rect 39529 9125 39574 9153
rect 39568 9113 39574 9125
rect 39626 9113 39632 9165
rect 40624 9113 40630 9165
rect 40682 9153 40688 9165
rect 49840 9153 49846 9165
rect 40682 9125 49846 9153
rect 40682 9113 40688 9125
rect 49840 9113 49846 9125
rect 49898 9113 49904 9165
rect 49939 9156 49997 9162
rect 49939 9122 49951 9156
rect 49985 9153 49997 9156
rect 54448 9153 54454 9165
rect 49985 9125 54454 9153
rect 49985 9122 49997 9125
rect 49939 9116 49997 9122
rect 54448 9113 54454 9125
rect 54506 9113 54512 9165
rect 8578 9079 8606 9113
rect 7968 9051 8126 9079
rect 8544 9051 8606 9079
rect 8098 9017 8126 9051
rect 12592 9039 12598 9091
rect 12650 9079 12656 9091
rect 15664 9079 15670 9091
rect 12650 9051 15670 9079
rect 12650 9039 12656 9051
rect 15664 9039 15670 9051
rect 15722 9039 15728 9091
rect 54640 9079 54646 9091
rect 43186 9051 54494 9079
rect 54601 9051 54646 9079
rect 8080 8965 8086 9017
rect 8138 8965 8144 9017
rect 9040 8965 9046 9017
rect 9098 9005 9104 9017
rect 20848 9005 20854 9017
rect 9098 8977 20854 9005
rect 9098 8965 9104 8977
rect 20848 8965 20854 8977
rect 20906 8965 20912 9017
rect 40048 8965 40054 9017
rect 40106 9005 40112 9017
rect 43186 9005 43214 9051
rect 53392 9005 53398 9017
rect 40106 8977 43214 9005
rect 53353 8977 53398 9005
rect 40106 8965 40112 8977
rect 53392 8965 53398 8977
rect 53450 8965 53456 9017
rect 4723 8934 4781 8940
rect 4723 8900 4735 8934
rect 4769 8931 4781 8934
rect 5200 8931 5206 8943
rect 4769 8903 5206 8931
rect 4769 8900 4781 8903
rect 4723 8894 4781 8900
rect 5200 8891 5206 8903
rect 5258 8891 5264 8943
rect 8656 8891 8662 8943
rect 8714 8891 8720 8943
rect 11248 8931 11254 8943
rect 9058 8903 11254 8931
rect 8083 8860 8141 8866
rect 8083 8826 8095 8860
rect 8129 8857 8141 8860
rect 8674 8857 8702 8891
rect 9058 8869 9086 8903
rect 11248 8891 11254 8903
rect 11306 8891 11312 8943
rect 11440 8891 11446 8943
rect 11498 8931 11504 8943
rect 13168 8931 13174 8943
rect 11498 8903 13174 8931
rect 11498 8891 11504 8903
rect 13168 8891 13174 8903
rect 13226 8891 13232 8943
rect 32272 8891 32278 8943
rect 32330 8931 32336 8943
rect 42928 8931 42934 8943
rect 32330 8903 42934 8931
rect 32330 8891 32336 8903
rect 42928 8891 42934 8903
rect 42986 8891 42992 8943
rect 44656 8891 44662 8943
rect 44714 8931 44720 8943
rect 50707 8934 50765 8940
rect 50707 8931 50719 8934
rect 44714 8903 50719 8931
rect 44714 8891 44720 8903
rect 50707 8900 50719 8903
rect 50753 8900 50765 8934
rect 50707 8894 50765 8900
rect 52147 8934 52205 8940
rect 52147 8900 52159 8934
rect 52193 8900 52205 8934
rect 54466 8931 54494 9051
rect 54640 9039 54646 9051
rect 54698 9039 54704 9091
rect 55411 9082 55469 9088
rect 55411 9048 55423 9082
rect 55457 9048 55469 9082
rect 55411 9042 55469 9048
rect 54544 8965 54550 9017
rect 54602 9005 54608 9017
rect 55426 9005 55454 9042
rect 54602 8977 55454 9005
rect 56563 9008 56621 9014
rect 54602 8965 54608 8977
rect 56563 8974 56575 9008
rect 56609 8974 56621 9008
rect 57232 9005 57238 9017
rect 57193 8977 57238 9005
rect 56563 8968 56621 8974
rect 55027 8934 55085 8940
rect 55027 8931 55039 8934
rect 54466 8903 55039 8931
rect 52147 8894 52205 8900
rect 55027 8900 55039 8903
rect 55073 8931 55085 8934
rect 55315 8934 55373 8940
rect 55315 8931 55327 8934
rect 55073 8903 55327 8931
rect 55073 8900 55085 8903
rect 55027 8894 55085 8900
rect 55315 8900 55327 8903
rect 55361 8900 55373 8934
rect 56578 8931 56606 8968
rect 57232 8965 57238 8977
rect 57290 8965 57296 9017
rect 57328 8931 57334 8943
rect 56578 8903 57334 8931
rect 55315 8894 55373 8900
rect 8129 8829 8256 8857
rect 8674 8829 8832 8857
rect 8129 8826 8141 8829
rect 8083 8820 8141 8826
rect 9040 8817 9046 8869
rect 9098 8817 9104 8869
rect 10960 8817 10966 8869
rect 11018 8857 11024 8869
rect 11344 8857 11350 8869
rect 11018 8829 11350 8857
rect 11018 8817 11024 8829
rect 11344 8817 11350 8829
rect 11402 8817 11408 8869
rect 13936 8817 13942 8869
rect 13994 8857 14000 8869
rect 16144 8857 16150 8869
rect 13994 8829 16150 8857
rect 13994 8817 14000 8829
rect 16144 8817 16150 8829
rect 16202 8817 16208 8869
rect 17008 8817 17014 8869
rect 17066 8857 17072 8869
rect 52162 8857 52190 8894
rect 57328 8891 57334 8903
rect 57386 8891 57392 8943
rect 55984 8857 55990 8869
rect 17066 8829 52190 8857
rect 53314 8829 55990 8857
rect 17066 8817 17072 8829
rect 9424 8743 9430 8795
rect 9482 8783 9488 8795
rect 14992 8783 14998 8795
rect 9482 8755 14998 8783
rect 9482 8743 9488 8755
rect 14992 8743 14998 8755
rect 15050 8743 15056 8795
rect 23056 8743 23062 8795
rect 23114 8783 23120 8795
rect 29008 8783 29014 8795
rect 23114 8755 29014 8783
rect 23114 8743 23120 8755
rect 29008 8743 29014 8755
rect 29066 8743 29072 8795
rect 36208 8743 36214 8795
rect 36266 8783 36272 8795
rect 46384 8783 46390 8795
rect 36266 8755 46390 8783
rect 36266 8743 36272 8755
rect 46384 8743 46390 8755
rect 46442 8743 46448 8795
rect 53314 8792 53342 8829
rect 55984 8817 55990 8829
rect 56042 8817 56048 8869
rect 53299 8786 53357 8792
rect 53299 8752 53311 8786
rect 53345 8752 53357 8786
rect 53299 8746 53357 8752
rect 53872 8743 53878 8795
rect 53930 8783 53936 8795
rect 54547 8786 54605 8792
rect 54547 8783 54559 8786
rect 53930 8755 54559 8783
rect 53930 8743 53936 8755
rect 54547 8752 54559 8755
rect 54593 8752 54605 8786
rect 54547 8746 54605 8752
rect 1152 8684 58848 8706
rect 1152 8632 19654 8684
rect 19706 8632 19718 8684
rect 19770 8632 19782 8684
rect 19834 8632 19846 8684
rect 19898 8632 50374 8684
rect 50426 8632 50438 8684
rect 50490 8632 50502 8684
rect 50554 8632 50566 8684
rect 50618 8632 58848 8684
rect 1152 8610 58848 8632
rect 2035 8564 2093 8570
rect 2035 8561 2047 8564
rect 1762 8533 2047 8561
rect 1762 8422 1790 8533
rect 2035 8530 2047 8533
rect 2081 8561 2093 8564
rect 3760 8561 3766 8573
rect 2081 8533 3766 8561
rect 2081 8530 2093 8533
rect 2035 8524 2093 8530
rect 3760 8521 3766 8533
rect 3818 8521 3824 8573
rect 9616 8521 9622 8573
rect 9674 8561 9680 8573
rect 10864 8561 10870 8573
rect 9674 8533 10870 8561
rect 9674 8521 9680 8533
rect 10864 8521 10870 8533
rect 10922 8521 10928 8573
rect 11536 8521 11542 8573
rect 11594 8561 11600 8573
rect 12019 8564 12077 8570
rect 12019 8561 12031 8564
rect 11594 8533 12031 8561
rect 11594 8521 11600 8533
rect 12019 8530 12031 8533
rect 12065 8530 12077 8564
rect 12019 8524 12077 8530
rect 12496 8521 12502 8573
rect 12554 8561 12560 8573
rect 29200 8561 29206 8573
rect 12554 8533 29206 8561
rect 12554 8521 12560 8533
rect 29200 8521 29206 8533
rect 29258 8521 29264 8573
rect 31216 8521 31222 8573
rect 31274 8561 31280 8573
rect 42640 8561 42646 8573
rect 31274 8533 42646 8561
rect 31274 8521 31280 8533
rect 42640 8521 42646 8533
rect 42698 8521 42704 8573
rect 46480 8521 46486 8573
rect 46538 8561 46544 8573
rect 47731 8564 47789 8570
rect 47731 8561 47743 8564
rect 46538 8533 47743 8561
rect 46538 8521 46544 8533
rect 47731 8530 47743 8533
rect 47777 8561 47789 8564
rect 47827 8564 47885 8570
rect 47827 8561 47839 8564
rect 47777 8533 47839 8561
rect 47777 8530 47789 8533
rect 47731 8524 47789 8530
rect 47827 8530 47839 8533
rect 47873 8530 47885 8564
rect 47827 8524 47885 8530
rect 47920 8521 47926 8573
rect 47978 8561 47984 8573
rect 52336 8561 52342 8573
rect 47978 8533 52342 8561
rect 47978 8521 47984 8533
rect 52336 8521 52342 8533
rect 52394 8521 52400 8573
rect 52531 8564 52589 8570
rect 52531 8530 52543 8564
rect 52577 8561 52589 8564
rect 58960 8561 58966 8573
rect 52577 8533 58966 8561
rect 52577 8530 52589 8533
rect 52531 8524 52589 8530
rect 58960 8521 58966 8533
rect 59018 8521 59024 8573
rect 7600 8447 7606 8499
rect 7658 8487 7664 8499
rect 9331 8490 9389 8496
rect 9331 8487 9343 8490
rect 7658 8459 9343 8487
rect 7658 8447 7664 8459
rect 9331 8456 9343 8459
rect 9377 8487 9389 8490
rect 9427 8490 9485 8496
rect 9427 8487 9439 8490
rect 9377 8459 9439 8487
rect 9377 8456 9389 8459
rect 9331 8450 9389 8456
rect 9427 8456 9439 8459
rect 9473 8456 9485 8490
rect 9427 8450 9485 8456
rect 10594 8459 13118 8487
rect 1747 8416 1805 8422
rect 1747 8382 1759 8416
rect 1793 8382 1805 8416
rect 3280 8413 3286 8425
rect 3241 8385 3286 8413
rect 1747 8376 1805 8382
rect 3280 8373 3286 8385
rect 3338 8373 3344 8425
rect 10594 8422 10622 8459
rect 4531 8416 4589 8422
rect 4531 8382 4543 8416
rect 4577 8413 4589 8416
rect 10579 8416 10637 8422
rect 4577 8385 10046 8413
rect 4577 8382 4589 8385
rect 4531 8376 4589 8382
rect 2227 8342 2285 8348
rect 2227 8308 2239 8342
rect 2273 8339 2285 8342
rect 2515 8342 2573 8348
rect 2515 8339 2527 8342
rect 2273 8311 2527 8339
rect 2273 8308 2285 8311
rect 2227 8302 2285 8308
rect 2515 8308 2527 8311
rect 2561 8339 2573 8342
rect 5491 8342 5549 8348
rect 2561 8311 5438 8339
rect 2561 8308 2573 8311
rect 2515 8302 2573 8308
rect 1648 8265 1654 8277
rect 1609 8237 1654 8265
rect 1648 8225 1654 8237
rect 1706 8225 1712 8277
rect 2128 8225 2134 8277
rect 2186 8265 2192 8277
rect 2419 8268 2477 8274
rect 2419 8265 2431 8268
rect 2186 8237 2431 8265
rect 2186 8225 2192 8237
rect 2419 8234 2431 8237
rect 2465 8234 2477 8268
rect 2419 8228 2477 8234
rect 3187 8268 3245 8274
rect 3187 8234 3199 8268
rect 3233 8265 3245 8268
rect 3280 8265 3286 8277
rect 3233 8237 3286 8265
rect 3233 8234 3245 8237
rect 3187 8228 3245 8234
rect 3280 8225 3286 8237
rect 3338 8225 3344 8277
rect 4435 8268 4493 8274
rect 4435 8234 4447 8268
rect 4481 8234 4493 8268
rect 5410 8265 5438 8311
rect 5491 8308 5503 8342
rect 5537 8339 5549 8342
rect 5779 8342 5837 8348
rect 5779 8339 5791 8342
rect 5537 8311 5791 8339
rect 5537 8308 5549 8311
rect 5491 8302 5549 8308
rect 5779 8308 5791 8311
rect 5825 8339 5837 8342
rect 10018 8339 10046 8385
rect 10579 8382 10591 8416
rect 10625 8382 10637 8416
rect 10579 8376 10637 8382
rect 12208 8373 12214 8425
rect 12266 8413 12272 8425
rect 12803 8416 12861 8422
rect 12803 8413 12815 8416
rect 12266 8385 12815 8413
rect 12266 8373 12272 8385
rect 12803 8382 12815 8385
rect 12849 8382 12861 8416
rect 12803 8376 12861 8382
rect 12496 8339 12502 8351
rect 5825 8311 9950 8339
rect 10018 8311 12502 8339
rect 5825 8308 5837 8311
rect 5779 8302 5837 8308
rect 7600 8265 7606 8277
rect 5410 8237 7606 8265
rect 4435 8228 4493 8234
rect 4450 8191 4478 8228
rect 7600 8225 7606 8237
rect 7658 8225 7664 8277
rect 7696 8225 7702 8277
rect 7754 8265 7760 8277
rect 7795 8268 7853 8274
rect 7795 8265 7807 8268
rect 7754 8237 7807 8265
rect 7754 8225 7760 8237
rect 7795 8234 7807 8237
rect 7841 8234 7853 8268
rect 7795 8228 7853 8234
rect 7891 8268 7949 8274
rect 7891 8234 7903 8268
rect 7937 8265 7949 8268
rect 8560 8265 8566 8277
rect 7937 8237 8566 8265
rect 7937 8234 7949 8237
rect 7891 8228 7949 8234
rect 8560 8225 8566 8237
rect 8618 8225 8624 8277
rect 9331 8268 9389 8274
rect 9331 8234 9343 8268
rect 9377 8265 9389 8268
rect 9715 8268 9773 8274
rect 9715 8265 9727 8268
rect 9377 8237 9727 8265
rect 9377 8234 9389 8237
rect 9331 8228 9389 8234
rect 9715 8234 9727 8237
rect 9761 8234 9773 8268
rect 9715 8228 9773 8234
rect 9811 8268 9869 8274
rect 9811 8234 9823 8268
rect 9857 8234 9869 8268
rect 9811 8228 9869 8234
rect 4816 8191 4822 8203
rect 4450 8163 4822 8191
rect 4816 8151 4822 8163
rect 4874 8151 4880 8203
rect 5584 8151 5590 8203
rect 5642 8191 5648 8203
rect 9424 8191 9430 8203
rect 5642 8163 9430 8191
rect 5642 8151 5648 8163
rect 9424 8151 9430 8163
rect 9482 8151 9488 8203
rect 9520 8151 9526 8203
rect 9578 8191 9584 8203
rect 9826 8191 9854 8228
rect 9578 8163 9854 8191
rect 9922 8191 9950 8311
rect 12496 8299 12502 8311
rect 12554 8299 12560 8351
rect 12592 8299 12598 8351
rect 12650 8339 12656 8351
rect 12650 8311 12830 8339
rect 12650 8299 12656 8311
rect 10288 8225 10294 8277
rect 10346 8265 10352 8277
rect 10483 8268 10541 8274
rect 10483 8265 10495 8268
rect 10346 8237 10495 8265
rect 10346 8225 10352 8237
rect 10483 8234 10495 8237
rect 10529 8234 10541 8268
rect 10483 8228 10541 8234
rect 10672 8225 10678 8277
rect 10730 8265 10736 8277
rect 11251 8268 11309 8274
rect 11251 8265 11263 8268
rect 10730 8237 11263 8265
rect 10730 8225 10736 8237
rect 11251 8234 11263 8237
rect 11297 8234 11309 8268
rect 11251 8228 11309 8234
rect 11347 8268 11405 8274
rect 11347 8234 11359 8268
rect 11393 8265 11405 8268
rect 11440 8265 11446 8277
rect 11393 8237 11446 8265
rect 11393 8234 11405 8237
rect 11347 8228 11405 8234
rect 11440 8225 11446 8237
rect 11498 8225 11504 8277
rect 12112 8265 12118 8277
rect 12073 8237 12118 8265
rect 12112 8225 12118 8237
rect 12170 8225 12176 8277
rect 12802 8265 12830 8311
rect 12883 8268 12941 8274
rect 12883 8265 12895 8268
rect 12802 8237 12895 8265
rect 12883 8234 12895 8237
rect 12929 8234 12941 8268
rect 12883 8228 12941 8234
rect 12976 8191 12982 8203
rect 9922 8163 12982 8191
rect 9578 8151 9584 8163
rect 12976 8151 12982 8163
rect 13034 8151 13040 8203
rect 13090 8191 13118 8459
rect 13168 8447 13174 8499
rect 13226 8487 13232 8499
rect 46003 8490 46061 8496
rect 46003 8487 46015 8490
rect 13226 8459 46015 8487
rect 13226 8447 13232 8459
rect 46003 8456 46015 8459
rect 46049 8456 46061 8490
rect 46003 8450 46061 8456
rect 46210 8459 52574 8487
rect 13648 8373 13654 8425
rect 13706 8413 13712 8425
rect 13706 8385 13751 8413
rect 13706 8373 13712 8385
rect 16336 8373 16342 8425
rect 16394 8413 16400 8425
rect 20560 8413 20566 8425
rect 16394 8385 20566 8413
rect 16394 8373 16400 8385
rect 20560 8373 20566 8385
rect 20618 8373 20624 8425
rect 37939 8416 37997 8422
rect 37939 8413 37951 8416
rect 23026 8385 37951 8413
rect 16048 8299 16054 8351
rect 16106 8339 16112 8351
rect 16163 8342 16221 8348
rect 16163 8339 16175 8342
rect 16106 8311 16175 8339
rect 16106 8299 16112 8311
rect 16163 8308 16175 8311
rect 16209 8308 16221 8342
rect 16163 8302 16221 8308
rect 16432 8299 16438 8351
rect 16490 8339 16496 8351
rect 23026 8339 23054 8385
rect 37939 8382 37951 8385
rect 37985 8382 37997 8416
rect 46096 8413 46102 8425
rect 37939 8376 37997 8382
rect 38146 8385 46102 8413
rect 16490 8311 23054 8339
rect 25075 8342 25133 8348
rect 16490 8299 16496 8311
rect 25075 8308 25087 8342
rect 25121 8339 25133 8342
rect 38032 8339 38038 8351
rect 25121 8311 38038 8339
rect 25121 8308 25133 8311
rect 25075 8302 25133 8308
rect 38032 8299 38038 8311
rect 38090 8299 38096 8351
rect 13168 8225 13174 8277
rect 13226 8265 13232 8277
rect 13555 8268 13613 8274
rect 13555 8265 13567 8268
rect 13226 8237 13567 8265
rect 13226 8225 13232 8237
rect 13555 8234 13567 8237
rect 13601 8234 13613 8268
rect 13555 8228 13613 8234
rect 14800 8225 14806 8277
rect 14858 8265 14864 8277
rect 15952 8265 15958 8277
rect 14858 8237 15958 8265
rect 14858 8225 14864 8237
rect 15952 8225 15958 8237
rect 16010 8225 16016 8277
rect 16240 8265 16246 8277
rect 16201 8237 16246 8265
rect 16240 8225 16246 8237
rect 16298 8225 16304 8277
rect 16336 8225 16342 8277
rect 16394 8265 16400 8277
rect 16915 8268 16973 8274
rect 16915 8265 16927 8268
rect 16394 8237 16927 8265
rect 16394 8225 16400 8237
rect 16915 8234 16927 8237
rect 16961 8234 16973 8268
rect 16915 8228 16973 8234
rect 17008 8225 17014 8277
rect 17066 8265 17072 8277
rect 17066 8237 17111 8265
rect 17066 8225 17072 8237
rect 18832 8225 18838 8277
rect 18890 8265 18896 8277
rect 38146 8265 38174 8385
rect 46096 8373 46102 8385
rect 46154 8373 46160 8425
rect 38224 8299 38230 8351
rect 38282 8339 38288 8351
rect 46210 8339 46238 8459
rect 47731 8416 47789 8422
rect 47731 8382 47743 8416
rect 47777 8413 47789 8416
rect 48115 8416 48173 8422
rect 48115 8413 48127 8416
rect 47777 8385 48127 8413
rect 47777 8382 47789 8385
rect 47731 8376 47789 8382
rect 48115 8382 48127 8385
rect 48161 8382 48173 8416
rect 48115 8376 48173 8382
rect 48691 8416 48749 8422
rect 48691 8382 48703 8416
rect 48737 8413 48749 8416
rect 48880 8413 48886 8425
rect 48737 8385 48886 8413
rect 48737 8382 48749 8385
rect 48691 8376 48749 8382
rect 48880 8373 48886 8385
rect 48938 8373 48944 8425
rect 38282 8311 46238 8339
rect 38282 8299 38288 8311
rect 46384 8299 46390 8351
rect 46442 8339 46448 8351
rect 50515 8342 50573 8348
rect 50515 8339 50527 8342
rect 46442 8311 50527 8339
rect 46442 8299 46448 8311
rect 50515 8308 50527 8311
rect 50561 8339 50573 8342
rect 50707 8342 50765 8348
rect 50707 8339 50719 8342
rect 50561 8311 50719 8339
rect 50561 8308 50573 8311
rect 50515 8302 50573 8308
rect 50707 8308 50719 8311
rect 50753 8308 50765 8342
rect 50707 8302 50765 8308
rect 18890 8237 38174 8265
rect 18890 8225 18896 8237
rect 38800 8225 38806 8277
rect 38858 8265 38864 8277
rect 47536 8265 47542 8277
rect 38858 8237 47542 8265
rect 38858 8225 38864 8237
rect 47536 8225 47542 8237
rect 47594 8225 47600 8277
rect 48016 8225 48022 8277
rect 48074 8265 48080 8277
rect 48211 8268 48269 8274
rect 48211 8265 48223 8268
rect 48074 8237 48223 8265
rect 48074 8225 48080 8237
rect 48211 8234 48223 8237
rect 48257 8234 48269 8268
rect 48211 8228 48269 8234
rect 48688 8225 48694 8277
rect 48746 8265 48752 8277
rect 48979 8268 49037 8274
rect 48979 8265 48991 8268
rect 48746 8237 48991 8265
rect 48746 8225 48752 8237
rect 48979 8234 48991 8237
rect 49025 8234 49037 8268
rect 48979 8228 49037 8234
rect 49456 8225 49462 8277
rect 49514 8265 49520 8277
rect 49651 8268 49709 8274
rect 49651 8265 49663 8268
rect 49514 8237 49663 8265
rect 49514 8225 49520 8237
rect 49651 8234 49663 8237
rect 49697 8234 49709 8268
rect 49651 8228 49709 8234
rect 49747 8268 49805 8274
rect 49747 8234 49759 8268
rect 49793 8234 49805 8268
rect 52435 8268 52493 8274
rect 52435 8265 52447 8268
rect 49747 8228 49805 8234
rect 52162 8237 52447 8265
rect 25075 8194 25133 8200
rect 25075 8191 25087 8194
rect 13090 8163 25087 8191
rect 25075 8160 25087 8163
rect 25121 8160 25133 8194
rect 25075 8154 25133 8160
rect 25648 8151 25654 8203
rect 25706 8191 25712 8203
rect 29776 8191 29782 8203
rect 25706 8163 29438 8191
rect 29737 8163 29782 8191
rect 25706 8151 25712 8163
rect 4912 8077 4918 8129
rect 4970 8117 4976 8129
rect 24208 8117 24214 8129
rect 4970 8089 24214 8117
rect 4970 8077 4976 8089
rect 24208 8077 24214 8089
rect 24266 8077 24272 8129
rect 24400 8077 24406 8129
rect 24458 8117 24464 8129
rect 29296 8117 29302 8129
rect 24458 8089 29302 8117
rect 24458 8077 24464 8089
rect 29296 8077 29302 8089
rect 29354 8077 29360 8129
rect 29410 8117 29438 8163
rect 29776 8151 29782 8163
rect 29834 8151 29840 8203
rect 37939 8194 37997 8200
rect 37939 8160 37951 8194
rect 37985 8191 37997 8194
rect 49762 8191 49790 8228
rect 37985 8163 49790 8191
rect 37985 8160 37997 8163
rect 37939 8154 37997 8160
rect 29968 8117 29974 8129
rect 29410 8089 29974 8117
rect 29968 8077 29974 8089
rect 30026 8077 30032 8129
rect 30931 8120 30989 8126
rect 30931 8086 30943 8120
rect 30977 8117 30989 8120
rect 32944 8117 32950 8129
rect 30977 8089 32950 8117
rect 30977 8086 30989 8089
rect 30931 8080 30989 8086
rect 32944 8077 32950 8089
rect 33002 8077 33008 8129
rect 33232 8077 33238 8129
rect 33290 8117 33296 8129
rect 34387 8120 34445 8126
rect 34387 8117 34399 8120
rect 33290 8089 34399 8117
rect 33290 8077 33296 8089
rect 34387 8086 34399 8089
rect 34433 8086 34445 8120
rect 34387 8080 34445 8086
rect 35059 8120 35117 8126
rect 35059 8086 35071 8120
rect 35105 8117 35117 8120
rect 39568 8117 39574 8129
rect 35105 8089 39574 8117
rect 35105 8086 35117 8089
rect 35059 8080 35117 8086
rect 39568 8077 39574 8089
rect 39626 8077 39632 8129
rect 41104 8077 41110 8129
rect 41162 8117 41168 8129
rect 46000 8117 46006 8129
rect 41162 8089 46006 8117
rect 41162 8077 41168 8089
rect 46000 8077 46006 8089
rect 46058 8077 46064 8129
rect 52162 8126 52190 8237
rect 52435 8234 52447 8237
rect 52481 8234 52493 8268
rect 52435 8228 52493 8234
rect 46195 8120 46253 8126
rect 46195 8086 46207 8120
rect 46241 8117 46253 8120
rect 52147 8120 52205 8126
rect 52147 8117 52159 8120
rect 46241 8089 52159 8117
rect 46241 8086 46253 8089
rect 46195 8080 46253 8086
rect 52147 8086 52159 8089
rect 52193 8086 52205 8120
rect 52546 8117 52574 8459
rect 52912 8339 52918 8351
rect 52873 8311 52918 8339
rect 52912 8299 52918 8311
rect 52970 8339 52976 8351
rect 53203 8342 53261 8348
rect 53203 8339 53215 8342
rect 52970 8311 53215 8339
rect 52970 8299 52976 8311
rect 53203 8308 53215 8311
rect 53249 8308 53261 8342
rect 53203 8302 53261 8308
rect 55219 8342 55277 8348
rect 55219 8308 55231 8342
rect 55265 8339 55277 8342
rect 55987 8342 56045 8348
rect 55265 8311 55934 8339
rect 55265 8308 55277 8311
rect 55219 8302 55277 8308
rect 53299 8268 53357 8274
rect 53299 8234 53311 8268
rect 53345 8234 53357 8268
rect 53299 8228 53357 8234
rect 53104 8151 53110 8203
rect 53162 8191 53168 8203
rect 53314 8191 53342 8228
rect 53488 8225 53494 8277
rect 53546 8265 53552 8277
rect 53971 8268 54029 8274
rect 53971 8265 53983 8268
rect 53546 8237 53983 8265
rect 53546 8225 53552 8237
rect 53971 8234 53983 8237
rect 54017 8234 54029 8268
rect 53971 8228 54029 8234
rect 54064 8225 54070 8277
rect 54122 8265 54128 8277
rect 54122 8237 54167 8265
rect 54122 8225 54128 8237
rect 53162 8163 53342 8191
rect 55906 8191 55934 8311
rect 55987 8308 55999 8342
rect 56033 8308 56045 8342
rect 55987 8302 56045 8308
rect 56002 8265 56030 8302
rect 56944 8299 56950 8351
rect 57002 8339 57008 8351
rect 57139 8342 57197 8348
rect 57139 8339 57151 8342
rect 57002 8311 57151 8339
rect 57002 8299 57008 8311
rect 57139 8308 57151 8311
rect 57185 8308 57197 8342
rect 57139 8302 57197 8308
rect 58384 8265 58390 8277
rect 56002 8237 58390 8265
rect 58384 8225 58390 8237
rect 58442 8225 58448 8277
rect 59824 8191 59830 8203
rect 55906 8163 59830 8191
rect 53162 8151 53168 8163
rect 59824 8151 59830 8163
rect 59882 8151 59888 8203
rect 54736 8117 54742 8129
rect 52546 8089 54742 8117
rect 52147 8080 52205 8086
rect 54736 8077 54742 8089
rect 54794 8077 54800 8129
rect 1152 8018 58848 8040
rect 1152 7966 4294 8018
rect 4346 7966 4358 8018
rect 4410 7966 4422 8018
rect 4474 7966 4486 8018
rect 4538 7966 35014 8018
rect 35066 7966 35078 8018
rect 35130 7966 35142 8018
rect 35194 7966 35206 8018
rect 35258 7966 58848 8018
rect 1152 7944 58848 7966
rect 3664 7895 3670 7907
rect 3625 7867 3670 7895
rect 3664 7855 3670 7867
rect 3722 7895 3728 7907
rect 3722 7867 4094 7895
rect 3722 7855 3728 7867
rect 3283 7750 3341 7756
rect 3283 7716 3295 7750
rect 3329 7747 3341 7750
rect 3376 7747 3382 7759
rect 3329 7719 3382 7747
rect 3329 7716 3341 7719
rect 3283 7710 3341 7716
rect 3376 7707 3382 7719
rect 3434 7707 3440 7759
rect 4066 7756 4094 7867
rect 7888 7855 7894 7907
rect 7946 7895 7952 7907
rect 8467 7898 8525 7904
rect 7946 7867 8030 7895
rect 7946 7855 7952 7867
rect 5299 7824 5357 7830
rect 5299 7790 5311 7824
rect 5345 7821 5357 7824
rect 5345 7793 5630 7821
rect 5345 7790 5357 7793
rect 5299 7784 5357 7790
rect 5602 7759 5630 7793
rect 4051 7750 4109 7756
rect 4051 7716 4063 7750
rect 4097 7716 4109 7750
rect 4051 7710 4109 7716
rect 4819 7750 4877 7756
rect 4819 7716 4831 7750
rect 4865 7747 4877 7750
rect 4912 7747 4918 7759
rect 4865 7719 4918 7747
rect 4865 7716 4877 7719
rect 4819 7710 4877 7716
rect 4912 7707 4918 7719
rect 4970 7707 4976 7759
rect 5584 7747 5590 7759
rect 5545 7719 5590 7747
rect 5584 7707 5590 7719
rect 5642 7707 5648 7759
rect 8002 7747 8030 7867
rect 8467 7864 8479 7898
rect 8513 7895 8525 7898
rect 9712 7895 9718 7907
rect 8513 7867 9718 7895
rect 8513 7864 8525 7867
rect 8467 7858 8525 7864
rect 9712 7855 9718 7867
rect 9770 7855 9776 7907
rect 9904 7855 9910 7907
rect 9962 7895 9968 7907
rect 12019 7898 12077 7904
rect 12019 7895 12031 7898
rect 9962 7867 12031 7895
rect 9962 7855 9968 7867
rect 12019 7864 12031 7867
rect 12065 7864 12077 7898
rect 12019 7858 12077 7864
rect 10000 7781 10006 7833
rect 10058 7821 10064 7833
rect 11440 7821 11446 7833
rect 10058 7793 11446 7821
rect 10058 7781 10064 7793
rect 11440 7781 11446 7793
rect 11498 7781 11504 7833
rect 7968 7719 8030 7747
rect 9139 7750 9197 7756
rect 9139 7716 9151 7750
rect 9185 7747 9197 7750
rect 9424 7747 9430 7759
rect 9185 7719 9430 7747
rect 9185 7716 9197 7719
rect 9139 7710 9197 7716
rect 9424 7707 9430 7719
rect 9482 7707 9488 7759
rect 9907 7750 9965 7756
rect 9907 7716 9919 7750
rect 9953 7747 9965 7750
rect 10192 7747 10198 7759
rect 9953 7719 10198 7747
rect 9953 7716 9965 7719
rect 9907 7710 9965 7716
rect 10192 7707 10198 7719
rect 10250 7707 10256 7759
rect 11920 7747 11926 7759
rect 10306 7719 11926 7747
rect 8518 7685 8570 7691
rect 1456 7633 1462 7685
rect 1514 7673 1520 7685
rect 1555 7676 1613 7682
rect 1555 7673 1567 7676
rect 1514 7645 1567 7673
rect 1514 7633 1520 7645
rect 1555 7642 1567 7645
rect 1601 7642 1613 7676
rect 1555 7636 1613 7642
rect 8752 7633 8758 7685
rect 8810 7673 8816 7685
rect 10306 7673 10334 7719
rect 11920 7707 11926 7719
rect 11978 7707 11984 7759
rect 12034 7747 12062 7858
rect 12112 7855 12118 7907
rect 12170 7895 12176 7907
rect 12170 7867 13118 7895
rect 12170 7855 12176 7867
rect 12307 7750 12365 7756
rect 12307 7747 12319 7750
rect 12034 7719 12319 7747
rect 12307 7716 12319 7719
rect 12353 7716 12365 7750
rect 12307 7710 12365 7716
rect 8810 7645 10334 7673
rect 10963 7676 11021 7682
rect 8810 7633 8816 7645
rect 10963 7642 10975 7676
rect 11009 7673 11021 7676
rect 11056 7673 11062 7685
rect 11009 7645 11062 7673
rect 11009 7642 11021 7645
rect 10963 7636 11021 7642
rect 11056 7633 11062 7645
rect 11114 7633 11120 7685
rect 13090 7673 13118 7867
rect 15952 7855 15958 7907
rect 16010 7895 16016 7907
rect 25936 7895 25942 7907
rect 16010 7867 25790 7895
rect 25897 7867 25942 7895
rect 16010 7855 16016 7867
rect 25648 7821 25654 7833
rect 13186 7793 25654 7821
rect 13186 7756 13214 7793
rect 25648 7781 25654 7793
rect 25706 7781 25712 7833
rect 13171 7750 13229 7756
rect 13171 7716 13183 7750
rect 13217 7716 13229 7750
rect 13171 7710 13229 7716
rect 13264 7707 13270 7759
rect 13322 7747 13328 7759
rect 15376 7747 15382 7759
rect 13322 7719 15382 7747
rect 13322 7707 13328 7719
rect 15376 7707 15382 7719
rect 15434 7707 15440 7759
rect 15571 7750 15629 7756
rect 15571 7716 15583 7750
rect 15617 7747 15629 7750
rect 15760 7747 15766 7759
rect 15617 7719 15766 7747
rect 15617 7716 15629 7719
rect 15571 7710 15629 7716
rect 15760 7707 15766 7719
rect 15818 7707 15824 7759
rect 16144 7707 16150 7759
rect 16202 7747 16208 7759
rect 19315 7750 19373 7756
rect 19315 7747 19327 7750
rect 16202 7719 19327 7747
rect 16202 7707 16208 7719
rect 19315 7716 19327 7719
rect 19361 7716 19373 7750
rect 20944 7747 20950 7759
rect 20905 7719 20950 7747
rect 19315 7710 19373 7716
rect 20944 7707 20950 7719
rect 21002 7707 21008 7759
rect 23923 7750 23981 7756
rect 23923 7716 23935 7750
rect 23969 7747 23981 7750
rect 24016 7747 24022 7759
rect 23969 7719 24022 7747
rect 23969 7716 23981 7719
rect 23923 7710 23981 7716
rect 24016 7707 24022 7719
rect 24074 7707 24080 7759
rect 24688 7747 24694 7759
rect 24649 7719 24694 7747
rect 24688 7707 24694 7719
rect 24746 7707 24752 7759
rect 25456 7747 25462 7759
rect 25417 7719 25462 7747
rect 25456 7707 25462 7719
rect 25514 7707 25520 7759
rect 15472 7673 15478 7685
rect 13090 7645 15478 7673
rect 15472 7633 15478 7645
rect 15530 7633 15536 7685
rect 15664 7633 15670 7685
rect 15722 7673 15728 7685
rect 21040 7673 21046 7685
rect 15722 7645 21046 7673
rect 15722 7633 15728 7645
rect 21040 7633 21046 7645
rect 21098 7633 21104 7685
rect 25264 7633 25270 7685
rect 25322 7673 25328 7685
rect 25648 7673 25654 7685
rect 25322 7645 25654 7673
rect 25322 7633 25328 7645
rect 25648 7633 25654 7645
rect 25706 7633 25712 7685
rect 25762 7673 25790 7867
rect 25936 7855 25942 7867
rect 25994 7895 26000 7907
rect 29104 7895 29110 7907
rect 25994 7867 26174 7895
rect 29065 7867 29110 7895
rect 25994 7855 26000 7867
rect 26146 7756 26174 7867
rect 29104 7855 29110 7867
rect 29162 7855 29168 7907
rect 29200 7855 29206 7907
rect 29258 7895 29264 7907
rect 34864 7895 34870 7907
rect 29258 7867 34870 7895
rect 29258 7855 29264 7867
rect 34864 7855 34870 7867
rect 34922 7855 34928 7907
rect 37075 7898 37133 7904
rect 37075 7864 37087 7898
rect 37121 7895 37133 7898
rect 37121 7867 44318 7895
rect 37121 7864 37133 7867
rect 37075 7858 37133 7864
rect 26224 7781 26230 7833
rect 26282 7821 26288 7833
rect 28915 7824 28973 7830
rect 28915 7821 28927 7824
rect 26282 7793 28927 7821
rect 26282 7781 26288 7793
rect 28915 7790 28927 7793
rect 28961 7790 28973 7824
rect 28915 7784 28973 7790
rect 26131 7750 26189 7756
rect 26131 7716 26143 7750
rect 26177 7716 26189 7750
rect 28243 7750 28301 7756
rect 28243 7747 28255 7750
rect 26131 7710 26189 7716
rect 27970 7719 28255 7747
rect 27970 7682 27998 7719
rect 28243 7716 28255 7719
rect 28289 7716 28301 7750
rect 29122 7747 29150 7855
rect 29296 7781 29302 7833
rect 29354 7821 29360 7833
rect 44176 7821 44182 7833
rect 29354 7793 40382 7821
rect 29354 7781 29360 7793
rect 29395 7750 29453 7756
rect 29395 7747 29407 7750
rect 29122 7719 29407 7747
rect 28243 7710 28301 7716
rect 29395 7716 29407 7719
rect 29441 7716 29453 7750
rect 30160 7747 30166 7759
rect 30121 7719 30166 7747
rect 29395 7710 29453 7716
rect 30160 7707 30166 7719
rect 30218 7707 30224 7759
rect 30832 7747 30838 7759
rect 30793 7719 30838 7747
rect 30832 7707 30838 7719
rect 30890 7747 30896 7759
rect 31123 7750 31181 7756
rect 31123 7747 31135 7750
rect 30890 7719 31135 7747
rect 30890 7707 30896 7719
rect 31123 7716 31135 7719
rect 31169 7747 31181 7750
rect 31411 7750 31469 7756
rect 31411 7747 31423 7750
rect 31169 7719 31423 7747
rect 31169 7716 31181 7719
rect 31123 7710 31181 7716
rect 31411 7716 31423 7719
rect 31457 7716 31469 7750
rect 31411 7710 31469 7716
rect 34003 7750 34061 7756
rect 34003 7716 34015 7750
rect 34049 7747 34061 7750
rect 34291 7750 34349 7756
rect 34049 7719 34238 7747
rect 34049 7716 34061 7719
rect 34003 7710 34061 7716
rect 27955 7676 28013 7682
rect 27955 7673 27967 7676
rect 25762 7645 27967 7673
rect 27955 7642 27967 7645
rect 28001 7642 28013 7676
rect 27955 7636 28013 7642
rect 28528 7633 28534 7685
rect 28586 7673 28592 7685
rect 34210 7673 34238 7719
rect 34291 7716 34303 7750
rect 34337 7747 34349 7750
rect 34576 7747 34582 7759
rect 34337 7719 34582 7747
rect 34337 7716 34349 7719
rect 34291 7710 34349 7716
rect 34576 7707 34582 7719
rect 34634 7707 34640 7759
rect 36112 7747 36118 7759
rect 36073 7719 36118 7747
rect 36112 7707 36118 7719
rect 36170 7707 36176 7759
rect 36880 7747 36886 7759
rect 36841 7719 36886 7747
rect 36880 7707 36886 7719
rect 36938 7707 36944 7759
rect 38800 7747 38806 7759
rect 38761 7719 38806 7747
rect 38800 7707 38806 7719
rect 38858 7707 38864 7759
rect 39568 7747 39574 7759
rect 39529 7719 39574 7747
rect 39568 7707 39574 7719
rect 39626 7707 39632 7759
rect 40354 7756 40382 7793
rect 41890 7793 44182 7821
rect 40339 7750 40397 7756
rect 40339 7716 40351 7750
rect 40385 7716 40397 7750
rect 41104 7747 41110 7759
rect 41065 7719 41110 7747
rect 40339 7710 40397 7716
rect 41104 7707 41110 7719
rect 41162 7707 41168 7759
rect 41890 7756 41918 7793
rect 44176 7781 44182 7793
rect 44234 7781 44240 7833
rect 44290 7821 44318 7867
rect 44368 7855 44374 7907
rect 44426 7895 44432 7907
rect 44467 7898 44525 7904
rect 44467 7895 44479 7898
rect 44426 7867 44479 7895
rect 44426 7855 44432 7867
rect 44467 7864 44479 7867
rect 44513 7895 44525 7898
rect 45232 7895 45238 7907
rect 44513 7867 44798 7895
rect 45193 7867 45238 7895
rect 44513 7864 44525 7867
rect 44467 7858 44525 7864
rect 44656 7821 44662 7833
rect 44290 7793 44662 7821
rect 44656 7781 44662 7793
rect 44714 7781 44720 7833
rect 41875 7750 41933 7756
rect 41875 7716 41887 7750
rect 41921 7716 41933 7750
rect 42640 7747 42646 7759
rect 42601 7719 42646 7747
rect 41875 7710 41933 7716
rect 42640 7707 42646 7719
rect 42698 7707 42704 7759
rect 44770 7756 44798 7867
rect 45232 7855 45238 7867
rect 45290 7895 45296 7907
rect 51184 7895 51190 7907
rect 45290 7867 45566 7895
rect 45290 7855 45296 7867
rect 45538 7756 45566 7867
rect 46402 7867 51190 7895
rect 46000 7781 46006 7833
rect 46058 7821 46064 7833
rect 46402 7821 46430 7867
rect 51184 7855 51190 7867
rect 51242 7855 51248 7907
rect 51856 7855 51862 7907
rect 51914 7895 51920 7907
rect 53008 7895 53014 7907
rect 51914 7867 53014 7895
rect 51914 7855 51920 7867
rect 53008 7855 53014 7867
rect 53066 7855 53072 7907
rect 46058 7793 46430 7821
rect 46058 7781 46064 7793
rect 46480 7781 46486 7833
rect 46538 7821 46544 7833
rect 46675 7824 46733 7830
rect 46675 7821 46687 7824
rect 46538 7793 46687 7821
rect 46538 7781 46544 7793
rect 46675 7790 46687 7793
rect 46721 7821 46733 7824
rect 46771 7824 46829 7830
rect 46771 7821 46783 7824
rect 46721 7793 46783 7821
rect 46721 7790 46733 7793
rect 46675 7784 46733 7790
rect 46771 7790 46783 7793
rect 46817 7790 46829 7824
rect 59344 7821 59350 7833
rect 46771 7784 46829 7790
rect 47170 7793 49502 7821
rect 44755 7750 44813 7756
rect 44755 7716 44767 7750
rect 44801 7716 44813 7750
rect 44755 7710 44813 7716
rect 45523 7750 45581 7756
rect 45523 7716 45535 7750
rect 45569 7716 45581 7750
rect 45523 7710 45581 7716
rect 45811 7750 45869 7756
rect 45811 7716 45823 7750
rect 45857 7747 45869 7750
rect 47170 7747 47198 7793
rect 45857 7719 47198 7747
rect 45857 7716 45869 7719
rect 45811 7710 45869 7716
rect 47248 7707 47254 7759
rect 47306 7747 47312 7759
rect 47923 7750 47981 7756
rect 47923 7747 47935 7750
rect 47306 7719 47935 7747
rect 47306 7707 47312 7719
rect 47923 7716 47935 7719
rect 47969 7716 47981 7750
rect 47923 7710 47981 7716
rect 48400 7707 48406 7759
rect 48458 7747 48464 7759
rect 49363 7750 49421 7756
rect 49363 7747 49375 7750
rect 48458 7719 49375 7747
rect 48458 7707 48464 7719
rect 49363 7716 49375 7719
rect 49409 7716 49421 7750
rect 49363 7710 49421 7716
rect 35248 7673 35254 7685
rect 28586 7645 34142 7673
rect 34210 7645 35254 7673
rect 28586 7633 28592 7645
rect 8518 7627 8570 7633
rect 2227 7602 2285 7608
rect 2227 7568 2239 7602
rect 2273 7599 2285 7602
rect 2512 7599 2518 7611
rect 2273 7571 2518 7599
rect 2273 7568 2285 7571
rect 2227 7562 2285 7568
rect 2512 7559 2518 7571
rect 2570 7559 2576 7611
rect 13651 7602 13709 7608
rect 13651 7568 13663 7602
rect 13697 7599 13709 7602
rect 13936 7599 13942 7611
rect 13697 7571 13942 7599
rect 13697 7568 13709 7571
rect 13651 7562 13709 7568
rect 13936 7559 13942 7571
rect 13994 7559 14000 7611
rect 14608 7559 14614 7611
rect 14666 7599 14672 7611
rect 18832 7599 18838 7611
rect 14666 7571 18838 7599
rect 14666 7559 14672 7571
rect 18832 7559 18838 7571
rect 18890 7559 18896 7611
rect 19315 7602 19373 7608
rect 19315 7568 19327 7602
rect 19361 7599 19373 7602
rect 26995 7602 27053 7608
rect 26995 7599 27007 7602
rect 19361 7571 27007 7599
rect 19361 7568 19373 7571
rect 19315 7562 19373 7568
rect 26995 7568 27007 7571
rect 27041 7568 27053 7602
rect 26995 7562 27053 7568
rect 27088 7559 27094 7611
rect 27146 7599 27152 7611
rect 29680 7599 29686 7611
rect 27146 7571 29686 7599
rect 27146 7559 27152 7571
rect 29680 7559 29686 7571
rect 29738 7559 29744 7611
rect 33808 7599 33814 7611
rect 33769 7571 33814 7599
rect 33808 7559 33814 7571
rect 33866 7559 33872 7611
rect 34114 7599 34142 7645
rect 35248 7633 35254 7645
rect 35306 7633 35312 7685
rect 35440 7633 35446 7685
rect 35498 7673 35504 7685
rect 48979 7676 49037 7682
rect 48979 7673 48991 7676
rect 35498 7645 48991 7673
rect 35498 7633 35504 7645
rect 48979 7642 48991 7645
rect 49025 7673 49037 7676
rect 49267 7676 49325 7682
rect 49267 7673 49279 7676
rect 49025 7645 49279 7673
rect 49025 7642 49037 7645
rect 48979 7636 49037 7642
rect 49267 7642 49279 7645
rect 49313 7642 49325 7676
rect 49267 7636 49325 7642
rect 35152 7599 35158 7611
rect 34114 7571 35158 7599
rect 35152 7559 35158 7571
rect 35210 7559 35216 7611
rect 35347 7602 35405 7608
rect 35347 7568 35359 7602
rect 35393 7568 35405 7602
rect 35347 7562 35405 7568
rect 8371 7528 8429 7534
rect 8371 7525 8383 7528
rect 8256 7497 8383 7525
rect 8371 7494 8383 7497
rect 8417 7494 8429 7528
rect 8371 7488 8429 7494
rect 8752 7485 8758 7537
rect 8810 7525 8816 7537
rect 9347 7528 9405 7534
rect 9347 7525 9359 7528
rect 8810 7497 9359 7525
rect 8810 7485 8816 7497
rect 9347 7494 9359 7497
rect 9393 7494 9405 7528
rect 9347 7488 9405 7494
rect 9904 7485 9910 7537
rect 9962 7525 9968 7537
rect 9962 7497 10910 7525
rect 9962 7485 9968 7497
rect 2320 7411 2326 7463
rect 2378 7451 2384 7463
rect 2419 7454 2477 7460
rect 2419 7451 2431 7454
rect 2378 7423 2431 7451
rect 2378 7411 2384 7423
rect 2419 7420 2431 7423
rect 2465 7420 2477 7454
rect 2419 7414 2477 7420
rect 2992 7411 2998 7463
rect 3050 7451 3056 7463
rect 3187 7454 3245 7460
rect 3187 7451 3199 7454
rect 3050 7423 3199 7451
rect 3050 7411 3056 7423
rect 3187 7420 3199 7423
rect 3233 7420 3245 7454
rect 3952 7451 3958 7463
rect 3913 7423 3958 7451
rect 3187 7414 3245 7420
rect 3952 7411 3958 7423
rect 4010 7411 4016 7463
rect 4048 7411 4054 7463
rect 4106 7451 4112 7463
rect 4723 7454 4781 7460
rect 4723 7451 4735 7454
rect 4106 7423 4735 7451
rect 4106 7411 4112 7423
rect 4723 7420 4735 7423
rect 4769 7420 4781 7454
rect 4723 7414 4781 7420
rect 5296 7411 5302 7463
rect 5354 7451 5360 7463
rect 5491 7454 5549 7460
rect 5491 7451 5503 7454
rect 5354 7423 5503 7451
rect 5354 7411 5360 7423
rect 5491 7420 5503 7423
rect 5537 7420 5549 7454
rect 7600 7451 7606 7463
rect 7561 7423 7606 7451
rect 5491 7414 5549 7420
rect 7600 7411 7606 7423
rect 7658 7411 7664 7463
rect 8560 7411 8566 7463
rect 8618 7411 8624 7463
rect 9136 7411 9142 7463
rect 9194 7451 9200 7463
rect 10882 7460 10910 7497
rect 11728 7485 11734 7537
rect 11786 7525 11792 7537
rect 11786 7497 12542 7525
rect 11786 7485 11792 7497
rect 10099 7454 10157 7460
rect 10099 7451 10111 7454
rect 9194 7423 10111 7451
rect 9194 7411 9200 7423
rect 10099 7420 10111 7423
rect 10145 7420 10157 7454
rect 10099 7414 10157 7420
rect 10867 7454 10925 7460
rect 10867 7420 10879 7454
rect 10913 7420 10925 7454
rect 10867 7414 10925 7420
rect 11056 7411 11062 7463
rect 11114 7451 11120 7463
rect 12403 7454 12461 7460
rect 12403 7451 12415 7454
rect 11114 7423 12415 7451
rect 11114 7411 11120 7423
rect 12403 7420 12415 7423
rect 12449 7420 12461 7454
rect 12514 7451 12542 7497
rect 12592 7485 12598 7537
rect 12650 7525 12656 7537
rect 13859 7528 13917 7534
rect 13859 7525 13871 7528
rect 12650 7497 13871 7525
rect 12650 7485 12656 7497
rect 13859 7494 13871 7497
rect 13905 7494 13917 7528
rect 13859 7488 13917 7494
rect 15280 7485 15286 7537
rect 15338 7525 15344 7537
rect 28528 7525 28534 7537
rect 15338 7497 28534 7525
rect 15338 7485 15344 7497
rect 28528 7485 28534 7497
rect 28586 7485 28592 7537
rect 28915 7528 28973 7534
rect 28915 7494 28927 7528
rect 28961 7525 28973 7528
rect 34003 7528 34061 7534
rect 34003 7525 34015 7528
rect 28961 7497 34015 7525
rect 28961 7494 28973 7497
rect 28915 7488 28973 7494
rect 34003 7494 34015 7497
rect 34049 7494 34061 7528
rect 35362 7525 35390 7562
rect 35536 7559 35542 7611
rect 35594 7599 35600 7611
rect 44083 7602 44141 7608
rect 35594 7571 41150 7599
rect 35594 7559 35600 7571
rect 37075 7528 37133 7534
rect 37075 7525 37087 7528
rect 35362 7497 37087 7525
rect 34003 7488 34061 7494
rect 37075 7494 37087 7497
rect 37121 7494 37133 7528
rect 37075 7488 37133 7494
rect 40048 7485 40054 7537
rect 40106 7525 40112 7537
rect 41122 7525 41150 7571
rect 44083 7568 44095 7602
rect 44129 7599 44141 7602
rect 45811 7602 45869 7608
rect 45811 7599 45823 7602
rect 44129 7571 45823 7599
rect 44129 7568 44141 7571
rect 44083 7562 44141 7568
rect 45811 7568 45823 7571
rect 45857 7568 45869 7602
rect 46000 7599 46006 7611
rect 45961 7571 46006 7599
rect 45811 7562 45869 7568
rect 46000 7559 46006 7571
rect 46058 7599 46064 7611
rect 46291 7602 46349 7608
rect 46291 7599 46303 7602
rect 46058 7571 46303 7599
rect 46058 7559 46064 7571
rect 46291 7568 46303 7571
rect 46337 7568 46349 7602
rect 46291 7562 46349 7568
rect 46675 7602 46733 7608
rect 46675 7568 46687 7602
rect 46721 7599 46733 7602
rect 47059 7602 47117 7608
rect 47059 7599 47071 7602
rect 46721 7571 47071 7599
rect 46721 7568 46733 7571
rect 46675 7562 46733 7568
rect 47059 7568 47071 7571
rect 47105 7568 47117 7602
rect 47059 7562 47117 7568
rect 47632 7559 47638 7611
rect 47690 7599 47696 7611
rect 47827 7602 47885 7608
rect 47827 7599 47839 7602
rect 47690 7571 47839 7599
rect 47690 7559 47696 7571
rect 47827 7568 47839 7571
rect 47873 7568 47885 7602
rect 49474 7599 49502 7793
rect 51010 7793 59350 7821
rect 50128 7747 50134 7759
rect 50089 7719 50134 7747
rect 50128 7707 50134 7719
rect 50186 7707 50192 7759
rect 51010 7756 51038 7793
rect 59344 7781 59350 7793
rect 59402 7781 59408 7833
rect 50995 7750 51053 7756
rect 50995 7716 51007 7750
rect 51041 7716 51053 7750
rect 50995 7710 51053 7716
rect 51571 7750 51629 7756
rect 51571 7716 51583 7750
rect 51617 7747 51629 7750
rect 51760 7747 51766 7759
rect 51617 7719 51766 7747
rect 51617 7716 51629 7719
rect 51571 7710 51629 7716
rect 51760 7707 51766 7719
rect 51818 7707 51824 7759
rect 52816 7707 52822 7759
rect 52874 7747 52880 7759
rect 53395 7750 53453 7756
rect 53395 7747 53407 7750
rect 52874 7719 53407 7747
rect 52874 7707 52880 7719
rect 53395 7716 53407 7719
rect 53441 7716 53453 7750
rect 58768 7747 58774 7759
rect 53395 7710 53453 7716
rect 55138 7719 58774 7747
rect 51091 7676 51149 7682
rect 51091 7642 51103 7676
rect 51137 7673 51149 7676
rect 53107 7676 53165 7682
rect 51137 7645 52766 7673
rect 51137 7642 51149 7645
rect 51091 7636 51149 7642
rect 51856 7599 51862 7611
rect 49474 7571 51862 7599
rect 47827 7562 47885 7568
rect 51856 7559 51862 7571
rect 51914 7559 51920 7611
rect 52627 7602 52685 7608
rect 52627 7568 52639 7602
rect 52673 7568 52685 7602
rect 52738 7599 52766 7645
rect 53107 7642 53119 7676
rect 53153 7673 53165 7676
rect 53200 7673 53206 7685
rect 53153 7645 53206 7673
rect 53153 7642 53165 7645
rect 53107 7636 53165 7642
rect 53200 7633 53206 7645
rect 53258 7673 53264 7685
rect 55138 7682 55166 7719
rect 58768 7707 58774 7719
rect 58826 7707 58832 7759
rect 53299 7676 53357 7682
rect 53299 7673 53311 7676
rect 53258 7645 53311 7673
rect 53258 7633 53264 7645
rect 53299 7642 53311 7645
rect 53345 7642 53357 7676
rect 53299 7636 53357 7642
rect 55123 7676 55181 7682
rect 55123 7642 55135 7676
rect 55169 7642 55181 7676
rect 55792 7673 55798 7685
rect 55753 7645 55798 7673
rect 55123 7636 55181 7642
rect 55792 7633 55798 7645
rect 55850 7633 55856 7685
rect 56176 7633 56182 7685
rect 56234 7673 56240 7685
rect 56563 7676 56621 7682
rect 56563 7673 56575 7676
rect 56234 7645 56575 7673
rect 56234 7633 56240 7645
rect 56563 7642 56575 7645
rect 56609 7642 56621 7676
rect 56563 7636 56621 7642
rect 56848 7633 56854 7685
rect 56906 7673 56912 7685
rect 57331 7676 57389 7682
rect 57331 7673 57343 7676
rect 56906 7645 57343 7673
rect 56906 7633 56912 7645
rect 57331 7642 57343 7645
rect 57377 7642 57389 7676
rect 57331 7636 57389 7642
rect 56272 7599 56278 7611
rect 52738 7571 56278 7599
rect 52627 7562 52685 7568
rect 52642 7525 52670 7562
rect 56272 7559 56278 7571
rect 56330 7559 56336 7611
rect 40106 7497 41054 7525
rect 41122 7497 52670 7525
rect 40106 7485 40112 7497
rect 13075 7454 13133 7460
rect 13075 7451 13087 7454
rect 12514 7423 13087 7451
rect 12403 7414 12461 7420
rect 13075 7420 13087 7423
rect 13121 7420 13133 7454
rect 13075 7414 13133 7420
rect 13168 7411 13174 7463
rect 13226 7451 13232 7463
rect 15568 7451 15574 7463
rect 13226 7423 15574 7451
rect 13226 7411 13232 7423
rect 15568 7411 15574 7423
rect 15626 7411 15632 7463
rect 15664 7411 15670 7463
rect 15722 7451 15728 7463
rect 15859 7454 15917 7460
rect 15859 7451 15871 7454
rect 15722 7423 15871 7451
rect 15722 7411 15728 7423
rect 15859 7420 15871 7423
rect 15905 7420 15917 7454
rect 15859 7414 15917 7420
rect 20752 7411 20758 7463
rect 20810 7451 20816 7463
rect 20851 7454 20909 7460
rect 20851 7451 20863 7454
rect 20810 7423 20863 7451
rect 20810 7411 20816 7423
rect 20851 7420 20863 7423
rect 20897 7420 20909 7454
rect 20851 7414 20909 7420
rect 23728 7411 23734 7463
rect 23786 7451 23792 7463
rect 23827 7454 23885 7460
rect 23827 7451 23839 7454
rect 23786 7423 23839 7451
rect 23786 7411 23792 7423
rect 23827 7420 23839 7423
rect 23873 7420 23885 7454
rect 23827 7414 23885 7420
rect 24112 7411 24118 7463
rect 24170 7451 24176 7463
rect 24595 7454 24653 7460
rect 24595 7451 24607 7454
rect 24170 7423 24607 7451
rect 24170 7411 24176 7423
rect 24595 7420 24607 7423
rect 24641 7420 24653 7454
rect 24595 7414 24653 7420
rect 24784 7411 24790 7463
rect 24842 7451 24848 7463
rect 25363 7454 25421 7460
rect 25363 7451 25375 7454
rect 24842 7423 25375 7451
rect 24842 7411 24848 7423
rect 25363 7420 25375 7423
rect 25409 7420 25421 7454
rect 25363 7414 25421 7420
rect 25936 7411 25942 7463
rect 25994 7451 26000 7463
rect 26227 7454 26285 7460
rect 26227 7451 26239 7454
rect 25994 7423 26239 7451
rect 25994 7411 26000 7423
rect 26227 7420 26239 7423
rect 26273 7420 26285 7454
rect 26227 7414 26285 7420
rect 26704 7411 26710 7463
rect 26762 7451 26768 7463
rect 26899 7454 26957 7460
rect 26899 7451 26911 7454
rect 26762 7423 26911 7451
rect 26762 7411 26768 7423
rect 26899 7420 26911 7423
rect 26945 7420 26957 7454
rect 26899 7414 26957 7420
rect 28144 7411 28150 7463
rect 28202 7451 28208 7463
rect 28339 7454 28397 7460
rect 28339 7451 28351 7454
rect 28202 7423 28351 7451
rect 28202 7411 28208 7423
rect 28339 7420 28351 7423
rect 28385 7420 28397 7454
rect 28339 7414 28397 7420
rect 29200 7411 29206 7463
rect 29258 7451 29264 7463
rect 29299 7454 29357 7460
rect 29299 7451 29311 7454
rect 29258 7423 29311 7451
rect 29258 7411 29264 7423
rect 29299 7420 29311 7423
rect 29345 7420 29357 7454
rect 29299 7414 29357 7420
rect 29584 7411 29590 7463
rect 29642 7451 29648 7463
rect 30067 7454 30125 7460
rect 30067 7451 30079 7454
rect 29642 7423 30079 7451
rect 29642 7411 29648 7423
rect 30067 7420 30079 7423
rect 30113 7420 30125 7454
rect 30067 7414 30125 7420
rect 31120 7411 31126 7463
rect 31178 7451 31184 7463
rect 31219 7454 31277 7460
rect 31219 7451 31231 7454
rect 31178 7423 31231 7451
rect 31178 7411 31184 7423
rect 31219 7420 31231 7423
rect 31265 7420 31277 7454
rect 31219 7414 31277 7420
rect 33616 7411 33622 7463
rect 33674 7451 33680 7463
rect 33715 7454 33773 7460
rect 33715 7451 33727 7454
rect 33674 7423 33727 7451
rect 33674 7411 33680 7423
rect 33715 7420 33727 7423
rect 33761 7420 33773 7454
rect 33715 7414 33773 7420
rect 34384 7411 34390 7463
rect 34442 7451 34448 7463
rect 34483 7454 34541 7460
rect 34483 7451 34495 7454
rect 34442 7423 34495 7451
rect 34442 7411 34448 7423
rect 34483 7420 34495 7423
rect 34529 7420 34541 7454
rect 34483 7414 34541 7420
rect 34864 7411 34870 7463
rect 34922 7451 34928 7463
rect 35251 7454 35309 7460
rect 35251 7451 35263 7454
rect 34922 7423 35263 7451
rect 34922 7411 34928 7423
rect 35251 7420 35263 7423
rect 35297 7420 35309 7454
rect 35251 7414 35309 7420
rect 35824 7411 35830 7463
rect 35882 7451 35888 7463
rect 36019 7454 36077 7460
rect 36019 7451 36031 7454
rect 35882 7423 36031 7451
rect 35882 7411 35888 7423
rect 36019 7420 36031 7423
rect 36065 7420 36077 7454
rect 36019 7414 36077 7420
rect 36592 7411 36598 7463
rect 36650 7451 36656 7463
rect 36787 7454 36845 7460
rect 36787 7451 36799 7454
rect 36650 7423 36799 7451
rect 36650 7411 36656 7423
rect 36787 7420 36799 7423
rect 36833 7420 36845 7454
rect 36787 7414 36845 7420
rect 38032 7411 38038 7463
rect 38090 7451 38096 7463
rect 38707 7454 38765 7460
rect 38707 7451 38719 7454
rect 38090 7423 38719 7451
rect 38090 7411 38096 7423
rect 38707 7420 38719 7423
rect 38753 7420 38765 7454
rect 38707 7414 38765 7420
rect 38800 7411 38806 7463
rect 38858 7451 38864 7463
rect 39475 7454 39533 7460
rect 39475 7451 39487 7454
rect 38858 7423 39487 7451
rect 38858 7411 38864 7423
rect 39475 7420 39487 7423
rect 39521 7420 39533 7454
rect 39475 7414 39533 7420
rect 39568 7411 39574 7463
rect 39626 7451 39632 7463
rect 41026 7460 41054 7497
rect 40243 7454 40301 7460
rect 40243 7451 40255 7454
rect 39626 7423 40255 7451
rect 39626 7411 39632 7423
rect 40243 7420 40255 7423
rect 40289 7420 40301 7454
rect 40243 7414 40301 7420
rect 41011 7454 41069 7460
rect 41011 7420 41023 7454
rect 41057 7420 41069 7454
rect 41011 7414 41069 7420
rect 41392 7411 41398 7463
rect 41450 7451 41456 7463
rect 41779 7454 41837 7460
rect 41779 7451 41791 7454
rect 41450 7423 41791 7451
rect 41450 7411 41456 7423
rect 41779 7420 41791 7423
rect 41825 7420 41837 7454
rect 41779 7414 41837 7420
rect 42448 7411 42454 7463
rect 42506 7451 42512 7463
rect 42547 7454 42605 7460
rect 42547 7451 42559 7454
rect 42506 7423 42559 7451
rect 42506 7411 42512 7423
rect 42547 7420 42559 7423
rect 42593 7420 42605 7454
rect 42547 7414 42605 7420
rect 43888 7411 43894 7463
rect 43946 7451 43952 7463
rect 43987 7454 44045 7460
rect 43987 7451 43999 7454
rect 43946 7423 43999 7451
rect 43946 7411 43952 7423
rect 43987 7420 43999 7423
rect 44033 7420 44045 7454
rect 43987 7414 44045 7420
rect 44656 7411 44662 7463
rect 44714 7451 44720 7463
rect 44851 7454 44909 7460
rect 44851 7451 44863 7454
rect 44714 7423 44863 7451
rect 44714 7411 44720 7423
rect 44851 7420 44863 7423
rect 44897 7420 44909 7454
rect 44851 7414 44909 7420
rect 45040 7411 45046 7463
rect 45098 7451 45104 7463
rect 45619 7454 45677 7460
rect 45619 7451 45631 7454
rect 45098 7423 45631 7451
rect 45098 7411 45104 7423
rect 45619 7420 45631 7423
rect 45665 7420 45677 7454
rect 45619 7414 45677 7420
rect 45808 7411 45814 7463
rect 45866 7451 45872 7463
rect 46387 7454 46445 7460
rect 46387 7451 46399 7454
rect 45866 7423 46399 7451
rect 45866 7411 45872 7423
rect 46387 7420 46399 7423
rect 46433 7420 46445 7454
rect 46387 7414 46445 7420
rect 46480 7411 46486 7463
rect 46538 7451 46544 7463
rect 47155 7454 47213 7460
rect 47155 7451 47167 7454
rect 46538 7423 47167 7451
rect 46538 7411 46544 7423
rect 47155 7420 47167 7423
rect 47201 7420 47213 7454
rect 47632 7451 47638 7463
rect 47593 7423 47638 7451
rect 47155 7414 47213 7420
rect 47632 7411 47638 7423
rect 47690 7411 47696 7463
rect 50032 7451 50038 7463
rect 49993 7423 50038 7451
rect 50032 7411 50038 7423
rect 50090 7411 50096 7463
rect 51760 7411 51766 7463
rect 51818 7451 51824 7463
rect 51859 7454 51917 7460
rect 51859 7451 51871 7454
rect 51818 7423 51871 7451
rect 51818 7411 51824 7423
rect 51859 7420 51871 7423
rect 51905 7420 51917 7454
rect 51859 7414 51917 7420
rect 52336 7411 52342 7463
rect 52394 7451 52400 7463
rect 52531 7454 52589 7460
rect 52531 7451 52543 7454
rect 52394 7423 52543 7451
rect 52394 7411 52400 7423
rect 52531 7420 52543 7423
rect 52577 7420 52589 7454
rect 52531 7414 52589 7420
rect 1152 7352 58848 7374
rect 1152 7300 19654 7352
rect 19706 7300 19718 7352
rect 19770 7300 19782 7352
rect 19834 7300 19846 7352
rect 19898 7300 50374 7352
rect 50426 7300 50438 7352
rect 50490 7300 50502 7352
rect 50554 7300 50566 7352
rect 50618 7300 58848 7352
rect 1152 7278 58848 7300
rect 5203 7232 5261 7238
rect 5203 7198 5215 7232
rect 5249 7198 5261 7232
rect 5203 7192 5261 7198
rect 3664 7115 3670 7167
rect 3722 7155 3728 7167
rect 5218 7155 5246 7192
rect 6544 7189 6550 7241
rect 6602 7189 6608 7241
rect 6928 7189 6934 7241
rect 6986 7229 6992 7241
rect 7507 7232 7565 7238
rect 7507 7229 7519 7232
rect 6986 7201 7519 7229
rect 6986 7189 6992 7201
rect 7507 7198 7519 7201
rect 7553 7198 7565 7232
rect 7507 7192 7565 7198
rect 7600 7189 7606 7241
rect 7658 7229 7664 7241
rect 8560 7229 8566 7241
rect 7658 7201 8566 7229
rect 7658 7189 7664 7201
rect 8560 7189 8566 7201
rect 8618 7229 8624 7241
rect 12784 7229 12790 7241
rect 8618 7201 12790 7229
rect 8618 7189 8624 7201
rect 12784 7189 12790 7201
rect 12842 7189 12848 7241
rect 29296 7229 29302 7241
rect 12898 7201 29302 7229
rect 3722 7127 5246 7155
rect 6562 7155 6590 7189
rect 6562 7127 9950 7155
rect 3722 7115 3728 7127
rect 5011 7084 5069 7090
rect 5011 7050 5023 7084
rect 5057 7081 5069 7084
rect 5299 7084 5357 7090
rect 5299 7081 5311 7084
rect 5057 7053 5311 7081
rect 5057 7050 5069 7053
rect 5011 7044 5069 7050
rect 5299 7050 5311 7053
rect 5345 7081 5357 7084
rect 5392 7081 5398 7093
rect 5345 7053 5398 7081
rect 5345 7050 5357 7053
rect 5299 7044 5357 7050
rect 5392 7041 5398 7053
rect 5450 7041 5456 7093
rect 6547 7084 6605 7090
rect 6547 7050 6559 7084
rect 6593 7081 6605 7084
rect 6835 7084 6893 7090
rect 6835 7081 6847 7084
rect 6593 7053 6847 7081
rect 6593 7050 6605 7053
rect 6547 7044 6605 7050
rect 6835 7050 6847 7053
rect 6881 7081 6893 7084
rect 8752 7081 8758 7093
rect 6881 7053 8758 7081
rect 6881 7050 6893 7053
rect 6835 7044 6893 7050
rect 8752 7041 8758 7053
rect 8810 7041 8816 7093
rect 9520 7041 9526 7093
rect 9578 7041 9584 7093
rect 9922 7081 9950 7127
rect 10048 7115 10054 7167
rect 10106 7155 10112 7167
rect 12304 7155 12310 7167
rect 10106 7127 12310 7155
rect 10106 7115 10112 7127
rect 12304 7115 12310 7127
rect 12362 7115 12368 7167
rect 12898 7155 12926 7201
rect 29296 7189 29302 7201
rect 29354 7189 29360 7241
rect 29488 7189 29494 7241
rect 29546 7229 29552 7241
rect 54064 7229 54070 7241
rect 29546 7201 54070 7229
rect 29546 7189 29552 7201
rect 54064 7189 54070 7201
rect 54122 7189 54128 7241
rect 12418 7127 12926 7155
rect 11923 7084 11981 7090
rect 9922 7053 11774 7081
rect 1648 7007 1654 7019
rect 1609 6979 1654 7007
rect 1648 6967 1654 6979
rect 1706 6967 1712 7019
rect 2512 7007 2518 7019
rect 2473 6979 2518 7007
rect 2512 6967 2518 6979
rect 2570 6967 2576 7019
rect 7600 7007 7606 7019
rect 7561 6979 7606 7007
rect 7600 6967 7606 6979
rect 7658 6967 7664 7019
rect 9538 6945 9566 7041
rect 9808 6967 9814 7019
rect 9866 7007 9872 7019
rect 10003 7010 10061 7016
rect 9866 6979 9911 7007
rect 9866 6967 9872 6979
rect 10003 6976 10015 7010
rect 10049 7007 10061 7010
rect 10864 7007 10870 7019
rect 10049 6979 10870 7007
rect 10049 6976 10061 6979
rect 10003 6970 10061 6976
rect 10864 6967 10870 6979
rect 10922 6967 10928 7019
rect 11248 7007 11254 7019
rect 11209 6979 11254 7007
rect 11248 6967 11254 6979
rect 11306 6967 11312 7019
rect 11746 7007 11774 7053
rect 11923 7050 11935 7084
rect 11969 7081 11981 7084
rect 12208 7081 12214 7093
rect 11969 7053 12214 7081
rect 11969 7050 11981 7053
rect 11923 7044 11981 7050
rect 12208 7041 12214 7053
rect 12266 7041 12272 7093
rect 12418 7007 12446 7127
rect 13168 7115 13174 7167
rect 13226 7155 13232 7167
rect 14224 7155 14230 7167
rect 13226 7127 14230 7155
rect 13226 7115 13232 7127
rect 14224 7115 14230 7127
rect 14282 7115 14288 7167
rect 15280 7115 15286 7167
rect 15338 7155 15344 7167
rect 19024 7155 19030 7167
rect 15338 7127 19030 7155
rect 15338 7115 15344 7127
rect 19024 7115 19030 7127
rect 19082 7115 19088 7167
rect 19138 7127 20318 7155
rect 13072 7041 13078 7093
rect 13130 7081 13136 7093
rect 19138 7081 19166 7127
rect 13130 7053 19166 7081
rect 20083 7084 20141 7090
rect 13130 7041 13136 7053
rect 20083 7050 20095 7084
rect 20129 7081 20141 7084
rect 20176 7081 20182 7093
rect 20129 7053 20182 7081
rect 20129 7050 20141 7053
rect 20083 7044 20141 7050
rect 20176 7041 20182 7053
rect 20234 7041 20240 7093
rect 20290 7081 20318 7127
rect 20464 7115 20470 7167
rect 20522 7155 20528 7167
rect 23056 7155 23062 7167
rect 20522 7127 23062 7155
rect 20522 7115 20528 7127
rect 23056 7115 23062 7127
rect 23114 7115 23120 7167
rect 23152 7115 23158 7167
rect 23210 7155 23216 7167
rect 25168 7155 25174 7167
rect 23210 7127 25174 7155
rect 23210 7115 23216 7127
rect 25168 7115 25174 7127
rect 25226 7115 25232 7167
rect 25360 7155 25366 7167
rect 25321 7127 25366 7155
rect 25360 7115 25366 7127
rect 25418 7155 25424 7167
rect 25648 7155 25654 7167
rect 25418 7127 25654 7155
rect 25418 7115 25424 7127
rect 25648 7115 25654 7127
rect 25706 7115 25712 7167
rect 27107 7158 27165 7164
rect 27107 7155 27119 7158
rect 27010 7127 27119 7155
rect 21139 7084 21197 7090
rect 21139 7081 21151 7084
rect 20290 7053 21151 7081
rect 21139 7050 21151 7053
rect 21185 7050 21197 7084
rect 21139 7044 21197 7050
rect 21619 7084 21677 7090
rect 21619 7050 21631 7084
rect 21665 7081 21677 7084
rect 21904 7081 21910 7093
rect 21665 7053 21910 7081
rect 21665 7050 21677 7053
rect 21619 7044 21677 7050
rect 21904 7041 21910 7053
rect 21962 7041 21968 7093
rect 22672 7081 22678 7093
rect 22633 7053 22678 7081
rect 22672 7041 22678 7053
rect 22730 7041 22736 7093
rect 23920 7041 23926 7093
rect 23978 7081 23984 7093
rect 24211 7084 24269 7090
rect 24211 7081 24223 7084
rect 23978 7053 24223 7081
rect 23978 7041 23984 7053
rect 24211 7050 24223 7053
rect 24257 7050 24269 7084
rect 26416 7081 26422 7093
rect 26377 7053 26422 7081
rect 24211 7044 24269 7050
rect 26416 7041 26422 7053
rect 26474 7041 26480 7093
rect 26896 7041 26902 7093
rect 26954 7081 26960 7093
rect 27010 7081 27038 7127
rect 27107 7124 27119 7127
rect 27153 7124 27165 7158
rect 27107 7118 27165 7124
rect 27280 7115 27286 7167
rect 27338 7155 27344 7167
rect 30736 7155 30742 7167
rect 27338 7127 30742 7155
rect 27338 7115 27344 7127
rect 30736 7115 30742 7127
rect 30794 7115 30800 7167
rect 31312 7155 31318 7167
rect 30850 7127 31166 7155
rect 31273 7127 31318 7155
rect 27184 7081 27190 7093
rect 26954 7053 27038 7081
rect 27145 7053 27190 7081
rect 26954 7041 26960 7053
rect 27184 7041 27190 7053
rect 27242 7041 27248 7093
rect 28720 7081 28726 7093
rect 28681 7053 28726 7081
rect 28720 7041 28726 7053
rect 28778 7041 28784 7093
rect 29491 7084 29549 7090
rect 29491 7050 29503 7084
rect 29537 7081 29549 7084
rect 29776 7081 29782 7093
rect 29537 7053 29782 7081
rect 29537 7050 29549 7053
rect 29491 7044 29549 7050
rect 29776 7041 29782 7053
rect 29834 7041 29840 7093
rect 29872 7041 29878 7093
rect 29930 7081 29936 7093
rect 30850 7081 30878 7127
rect 29930 7053 30878 7081
rect 30931 7084 30989 7090
rect 29930 7041 29936 7053
rect 30931 7050 30943 7084
rect 30977 7081 30989 7084
rect 31024 7081 31030 7093
rect 30977 7053 31030 7081
rect 30977 7050 30989 7053
rect 30931 7044 30989 7050
rect 31024 7041 31030 7053
rect 31082 7041 31088 7093
rect 31138 7081 31166 7127
rect 31312 7115 31318 7127
rect 31370 7155 31376 7167
rect 31891 7158 31949 7164
rect 31891 7155 31903 7158
rect 31370 7127 31903 7155
rect 31370 7115 31376 7127
rect 31504 7081 31510 7093
rect 31138 7053 31510 7081
rect 31504 7041 31510 7053
rect 31562 7041 31568 7093
rect 31618 7090 31646 7127
rect 31891 7124 31903 7127
rect 31937 7124 31949 7158
rect 31891 7118 31949 7124
rect 32848 7115 32854 7167
rect 32906 7155 32912 7167
rect 39376 7155 39382 7167
rect 32906 7127 39382 7155
rect 32906 7115 32912 7127
rect 39376 7115 39382 7127
rect 39434 7115 39440 7167
rect 39856 7115 39862 7167
rect 39914 7155 39920 7167
rect 41411 7158 41469 7164
rect 41411 7155 41423 7158
rect 39914 7127 41423 7155
rect 39914 7115 39920 7127
rect 41411 7124 41423 7127
rect 41457 7124 41469 7158
rect 41411 7118 41469 7124
rect 41680 7115 41686 7167
rect 41738 7155 41744 7167
rect 42947 7158 43005 7164
rect 42947 7155 42959 7158
rect 41738 7127 42959 7155
rect 41738 7115 41744 7127
rect 42947 7124 42959 7127
rect 42993 7124 43005 7158
rect 51664 7155 51670 7167
rect 51625 7127 51670 7155
rect 42947 7118 43005 7124
rect 51664 7115 51670 7127
rect 51722 7155 51728 7167
rect 51722 7127 51998 7155
rect 51722 7115 51728 7127
rect 31603 7084 31661 7090
rect 31603 7050 31615 7084
rect 31649 7050 31661 7084
rect 31603 7044 31661 7050
rect 32179 7084 32237 7090
rect 32179 7050 32191 7084
rect 32225 7081 32237 7084
rect 32467 7084 32525 7090
rect 32467 7081 32479 7084
rect 32225 7053 32479 7081
rect 32225 7050 32237 7053
rect 32179 7044 32237 7050
rect 32467 7050 32479 7053
rect 32513 7081 32525 7084
rect 32656 7081 32662 7093
rect 32513 7053 32662 7081
rect 32513 7050 32525 7053
rect 32467 7044 32525 7050
rect 32656 7041 32662 7053
rect 32714 7041 32720 7093
rect 32947 7084 33005 7090
rect 32947 7050 32959 7084
rect 32993 7081 33005 7084
rect 33235 7084 33293 7090
rect 33235 7081 33247 7084
rect 32993 7053 33247 7081
rect 32993 7050 33005 7053
rect 32947 7044 33005 7050
rect 33235 7050 33247 7053
rect 33281 7081 33293 7084
rect 34768 7081 34774 7093
rect 33281 7053 34622 7081
rect 34729 7053 34774 7081
rect 33281 7050 33293 7053
rect 33235 7044 33293 7050
rect 12688 7007 12694 7019
rect 11746 6979 12446 7007
rect 12649 6979 12694 7007
rect 12688 6967 12694 6979
rect 12746 6967 12752 7019
rect 12976 6967 12982 7019
rect 13034 7007 13040 7019
rect 27088 7007 27094 7019
rect 13034 6979 27094 7007
rect 13034 6967 13040 6979
rect 27088 6967 27094 6979
rect 27146 6967 27152 7019
rect 29680 6967 29686 7019
rect 29738 7007 29744 7019
rect 34480 7007 34486 7019
rect 29738 6979 34486 7007
rect 29738 6967 29744 6979
rect 34480 6967 34486 6979
rect 34538 6967 34544 7019
rect 34594 7007 34622 7053
rect 34768 7041 34774 7053
rect 34826 7041 34832 7093
rect 36976 7081 36982 7093
rect 34882 7053 36830 7081
rect 36937 7053 36982 7081
rect 34882 7007 34910 7053
rect 34594 6979 34910 7007
rect 36211 7010 36269 7016
rect 36211 6976 36223 7010
rect 36257 7007 36269 7010
rect 36688 7007 36694 7019
rect 36257 6979 36694 7007
rect 36257 6976 36269 6979
rect 36211 6970 36269 6976
rect 36688 6967 36694 6979
rect 36746 6967 36752 7019
rect 36802 7007 36830 7053
rect 36976 7041 36982 7053
rect 37034 7041 37040 7093
rect 39283 7084 39341 7090
rect 39283 7050 39295 7084
rect 39329 7081 39341 7084
rect 41776 7081 41782 7093
rect 39329 7053 41782 7081
rect 39329 7050 39341 7053
rect 39283 7044 39341 7050
rect 41776 7041 41782 7053
rect 41834 7041 41840 7093
rect 42256 7081 42262 7093
rect 42217 7053 42262 7081
rect 42256 7041 42262 7053
rect 42314 7041 42320 7093
rect 44275 7084 44333 7090
rect 44275 7050 44287 7084
rect 44321 7081 44333 7084
rect 44464 7081 44470 7093
rect 44321 7053 44470 7081
rect 44321 7050 44333 7053
rect 44275 7044 44333 7050
rect 44464 7041 44470 7053
rect 44522 7041 44528 7093
rect 48304 7081 48310 7093
rect 48265 7053 48310 7081
rect 48304 7041 48310 7053
rect 48362 7041 48368 7093
rect 50035 7084 50093 7090
rect 50035 7050 50047 7084
rect 50081 7081 50093 7084
rect 50224 7081 50230 7093
rect 50081 7053 50230 7081
rect 50081 7050 50093 7053
rect 50035 7044 50093 7050
rect 50224 7041 50230 7053
rect 50282 7041 50288 7093
rect 51970 7090 51998 7127
rect 51955 7084 52013 7090
rect 51955 7050 51967 7084
rect 52001 7050 52013 7084
rect 51955 7044 52013 7050
rect 38320 7007 38326 7019
rect 36802 6979 38326 7007
rect 38320 6967 38326 6979
rect 38378 6967 38384 7019
rect 38608 6967 38614 7019
rect 38666 7007 38672 7019
rect 41203 7010 41261 7016
rect 38666 6979 39998 7007
rect 38666 6967 38672 6979
rect 4435 6936 4493 6942
rect 4435 6902 4447 6936
rect 4481 6902 4493 6936
rect 4435 6896 4493 6902
rect 4450 6859 4478 6896
rect 4528 6893 4534 6945
rect 4586 6933 4592 6945
rect 4586 6905 4631 6933
rect 4586 6893 4592 6905
rect 5872 6893 5878 6945
rect 5930 6933 5936 6945
rect 5971 6936 6029 6942
rect 5971 6933 5983 6936
rect 5930 6905 5983 6933
rect 5930 6893 5936 6905
rect 5971 6902 5983 6905
rect 6017 6902 6029 6936
rect 5971 6896 6029 6902
rect 6067 6936 6125 6942
rect 6067 6902 6079 6936
rect 6113 6933 6125 6936
rect 6160 6933 6166 6945
rect 6113 6905 6166 6933
rect 6113 6902 6125 6905
rect 6067 6896 6125 6902
rect 6160 6893 6166 6905
rect 6218 6893 6224 6945
rect 6544 6893 6550 6945
rect 6602 6933 6608 6945
rect 6739 6936 6797 6942
rect 6739 6933 6751 6936
rect 6602 6905 6751 6933
rect 6602 6893 6608 6905
rect 6739 6902 6751 6905
rect 6785 6902 6797 6936
rect 8275 6936 8333 6942
rect 8275 6933 8287 6936
rect 6739 6896 6797 6902
rect 7522 6905 8287 6933
rect 5008 6859 5014 6871
rect 4450 6831 5014 6859
rect 5008 6819 5014 6831
rect 5066 6819 5072 6871
rect 7312 6819 7318 6871
rect 7370 6859 7376 6871
rect 7522 6859 7550 6905
rect 8275 6902 8287 6905
rect 8321 6902 8333 6936
rect 8275 6896 8333 6902
rect 8371 6936 8429 6942
rect 8371 6902 8383 6936
rect 8417 6902 8429 6936
rect 8371 6896 8429 6902
rect 7370 6831 7550 6859
rect 8083 6862 8141 6868
rect 7370 6819 7376 6831
rect 8083 6828 8095 6862
rect 8129 6859 8141 6862
rect 8386 6859 8414 6896
rect 9520 6893 9526 6945
rect 9578 6893 9584 6945
rect 9712 6933 9718 6945
rect 9673 6905 9718 6933
rect 9712 6893 9718 6905
rect 9770 6893 9776 6945
rect 9904 6893 9910 6945
rect 9962 6933 9968 6945
rect 10483 6936 10541 6942
rect 10483 6933 10495 6936
rect 9962 6905 10495 6933
rect 9962 6893 9968 6905
rect 10483 6902 10495 6905
rect 10529 6902 10541 6936
rect 10483 6896 10541 6902
rect 10576 6893 10582 6945
rect 10634 6933 10640 6945
rect 10634 6905 10679 6933
rect 10634 6893 10640 6905
rect 13456 6893 13462 6945
rect 13514 6933 13520 6945
rect 13555 6936 13613 6942
rect 13555 6933 13567 6936
rect 13514 6905 13567 6933
rect 13514 6893 13520 6905
rect 13555 6902 13567 6905
rect 13601 6902 13613 6936
rect 13555 6896 13613 6902
rect 13651 6936 13709 6942
rect 13651 6902 13663 6936
rect 13697 6933 13709 6936
rect 14512 6933 14518 6945
rect 13697 6905 14518 6933
rect 13697 6902 13709 6905
rect 13651 6896 13709 6902
rect 14512 6893 14518 6905
rect 14570 6893 14576 6945
rect 14608 6893 14614 6945
rect 14666 6933 14672 6945
rect 14995 6936 15053 6942
rect 14995 6933 15007 6936
rect 14666 6905 15007 6933
rect 14666 6893 14672 6905
rect 14995 6902 15007 6905
rect 15041 6902 15053 6936
rect 14995 6896 15053 6902
rect 15091 6936 15149 6942
rect 15091 6902 15103 6936
rect 15137 6933 15149 6936
rect 15280 6933 15286 6945
rect 15137 6905 15286 6933
rect 15137 6902 15149 6905
rect 15091 6896 15149 6902
rect 15280 6893 15286 6905
rect 15338 6893 15344 6945
rect 15376 6893 15382 6945
rect 15434 6933 15440 6945
rect 15763 6936 15821 6942
rect 15763 6933 15775 6936
rect 15434 6905 15775 6933
rect 15434 6893 15440 6905
rect 15763 6902 15775 6905
rect 15809 6902 15821 6936
rect 15763 6896 15821 6902
rect 15856 6893 15862 6945
rect 15914 6933 15920 6945
rect 15914 6905 15959 6933
rect 15914 6893 15920 6905
rect 17104 6893 17110 6945
rect 17162 6933 17168 6945
rect 17203 6936 17261 6942
rect 17203 6933 17215 6936
rect 17162 6905 17215 6933
rect 17162 6893 17168 6905
rect 17203 6902 17215 6905
rect 17249 6902 17261 6936
rect 17203 6896 17261 6902
rect 17296 6893 17302 6945
rect 17354 6933 17360 6945
rect 17776 6933 17782 6945
rect 17354 6905 17399 6933
rect 17737 6905 17782 6933
rect 17354 6893 17360 6905
rect 17776 6893 17782 6905
rect 17834 6893 17840 6945
rect 17872 6893 17878 6945
rect 17930 6933 17936 6945
rect 17971 6936 18029 6942
rect 17971 6933 17983 6936
rect 17930 6905 17983 6933
rect 17930 6893 17936 6905
rect 17971 6902 17983 6905
rect 18017 6902 18029 6936
rect 17971 6896 18029 6902
rect 18067 6936 18125 6942
rect 18067 6902 18079 6936
rect 18113 6933 18125 6936
rect 18160 6933 18166 6945
rect 18113 6905 18166 6933
rect 18113 6902 18125 6905
rect 18067 6896 18125 6902
rect 18160 6893 18166 6905
rect 18218 6893 18224 6945
rect 18544 6893 18550 6945
rect 18602 6933 18608 6945
rect 18739 6936 18797 6942
rect 18739 6933 18751 6936
rect 18602 6905 18751 6933
rect 18602 6893 18608 6905
rect 18739 6902 18751 6905
rect 18785 6902 18797 6936
rect 18739 6896 18797 6902
rect 18835 6936 18893 6942
rect 18835 6902 18847 6936
rect 18881 6902 18893 6936
rect 18835 6896 18893 6902
rect 10000 6859 10006 6871
rect 8129 6831 8414 6859
rect 9961 6831 10006 6859
rect 8129 6828 8141 6831
rect 8083 6822 8141 6828
rect 8386 6785 8414 6831
rect 10000 6819 10006 6831
rect 10058 6819 10064 6871
rect 10291 6862 10349 6868
rect 10291 6828 10303 6862
rect 10337 6859 10349 6862
rect 10594 6859 10622 6893
rect 18850 6859 18878 6896
rect 19216 6893 19222 6945
rect 19274 6933 19280 6945
rect 20080 6933 20086 6945
rect 19274 6905 20086 6933
rect 19274 6893 19280 6905
rect 20080 6893 20086 6905
rect 20138 6893 20144 6945
rect 20272 6933 20278 6945
rect 20233 6905 20278 6933
rect 20272 6893 20278 6905
rect 20330 6893 20336 6945
rect 20371 6936 20429 6942
rect 20371 6902 20383 6936
rect 20417 6933 20429 6936
rect 20464 6933 20470 6945
rect 20417 6905 20470 6933
rect 20417 6902 20429 6905
rect 20371 6896 20429 6902
rect 20464 6893 20470 6905
rect 20522 6893 20528 6945
rect 20848 6893 20854 6945
rect 20906 6933 20912 6945
rect 21043 6936 21101 6942
rect 21043 6933 21055 6936
rect 20906 6905 21055 6933
rect 20906 6893 20912 6905
rect 21043 6902 21055 6905
rect 21089 6902 21101 6936
rect 21808 6933 21814 6945
rect 21769 6905 21814 6933
rect 21043 6896 21101 6902
rect 21808 6893 21814 6905
rect 21866 6893 21872 6945
rect 21904 6893 21910 6945
rect 21962 6933 21968 6945
rect 22579 6936 22637 6942
rect 22579 6933 22591 6936
rect 21962 6905 22591 6933
rect 21962 6893 21968 6905
rect 22579 6902 22591 6905
rect 22625 6902 22637 6936
rect 22579 6896 22637 6902
rect 22672 6893 22678 6945
rect 22730 6933 22736 6945
rect 23347 6936 23405 6942
rect 23347 6933 23359 6936
rect 22730 6905 23359 6933
rect 22730 6893 22736 6905
rect 23347 6902 23359 6905
rect 23393 6902 23405 6936
rect 23347 6896 23405 6902
rect 23443 6936 23501 6942
rect 23443 6902 23455 6936
rect 23489 6933 23501 6936
rect 23536 6933 23542 6945
rect 23489 6905 23542 6933
rect 23489 6902 23501 6905
rect 23443 6896 23501 6902
rect 23536 6893 23542 6905
rect 23594 6893 23600 6945
rect 24115 6936 24173 6942
rect 24115 6933 24127 6936
rect 23938 6905 24127 6933
rect 10337 6831 10622 6859
rect 18754 6831 18878 6859
rect 10337 6828 10349 6831
rect 10291 6822 10349 6828
rect 17488 6785 17494 6797
rect 8386 6757 17494 6785
rect 17488 6745 17494 6757
rect 17546 6745 17552 6797
rect 18547 6788 18605 6794
rect 18547 6754 18559 6788
rect 18593 6785 18605 6788
rect 18754 6785 18782 6831
rect 18928 6819 18934 6871
rect 18986 6859 18992 6871
rect 23824 6859 23830 6871
rect 18986 6831 23830 6859
rect 18986 6819 18992 6831
rect 23824 6819 23830 6831
rect 23882 6819 23888 6871
rect 22864 6785 22870 6797
rect 18593 6757 22870 6785
rect 18593 6754 18605 6757
rect 18547 6748 18605 6754
rect 22864 6745 22870 6757
rect 22922 6745 22928 6797
rect 23344 6745 23350 6797
rect 23402 6785 23408 6797
rect 23938 6785 23966 6905
rect 24115 6902 24127 6905
rect 24161 6902 24173 6936
rect 24115 6896 24173 6902
rect 24592 6893 24598 6945
rect 24650 6933 24656 6945
rect 25555 6936 25613 6942
rect 25555 6933 25567 6936
rect 24650 6905 25567 6933
rect 24650 6893 24656 6905
rect 25555 6902 25567 6905
rect 25601 6902 25613 6936
rect 25555 6896 25613 6902
rect 25648 6893 25654 6945
rect 25706 6933 25712 6945
rect 26320 6933 26326 6945
rect 25706 6905 25751 6933
rect 26281 6905 26326 6933
rect 25706 6893 25712 6905
rect 26320 6893 26326 6905
rect 26378 6893 26384 6945
rect 27859 6936 27917 6942
rect 27859 6902 27871 6936
rect 27905 6902 27917 6936
rect 27859 6896 27917 6902
rect 26992 6819 26998 6871
rect 27050 6859 27056 6871
rect 27874 6859 27902 6896
rect 27952 6893 27958 6945
rect 28010 6933 28016 6945
rect 28624 6933 28630 6945
rect 28010 6905 28055 6933
rect 28585 6905 28630 6933
rect 28010 6893 28016 6905
rect 28624 6893 28630 6905
rect 28682 6893 28688 6945
rect 29411 6936 29469 6942
rect 29411 6902 29423 6936
rect 29457 6933 29469 6936
rect 29457 6905 29534 6933
rect 29457 6902 29469 6905
rect 29411 6896 29469 6902
rect 27050 6831 27902 6859
rect 27050 6819 27056 6831
rect 23402 6757 23966 6785
rect 23402 6745 23408 6757
rect 28528 6745 28534 6797
rect 28586 6785 28592 6797
rect 29506 6785 29534 6905
rect 29968 6893 29974 6945
rect 30026 6933 30032 6945
rect 30835 6936 30893 6942
rect 30835 6933 30847 6936
rect 30026 6905 30847 6933
rect 30026 6893 30032 6905
rect 30835 6902 30847 6905
rect 30881 6902 30893 6936
rect 30835 6896 30893 6902
rect 31699 6936 31757 6942
rect 31699 6902 31711 6936
rect 31745 6933 31757 6936
rect 31984 6933 31990 6945
rect 31745 6905 31990 6933
rect 31745 6902 31757 6905
rect 31699 6896 31757 6902
rect 31984 6893 31990 6905
rect 32042 6893 32048 6945
rect 32368 6933 32374 6945
rect 32329 6905 32374 6933
rect 32368 6893 32374 6905
rect 32426 6893 32432 6945
rect 32464 6893 32470 6945
rect 32522 6933 32528 6945
rect 33139 6936 33197 6942
rect 33139 6933 33151 6936
rect 32522 6905 33151 6933
rect 32522 6893 32528 6905
rect 33139 6902 33151 6905
rect 33185 6902 33197 6936
rect 33904 6933 33910 6945
rect 33865 6905 33910 6933
rect 33139 6896 33197 6902
rect 33904 6893 33910 6905
rect 33962 6893 33968 6945
rect 34003 6936 34061 6942
rect 34003 6902 34015 6936
rect 34049 6933 34061 6936
rect 34096 6933 34102 6945
rect 34049 6905 34102 6933
rect 34049 6902 34061 6905
rect 34003 6896 34061 6902
rect 34096 6893 34102 6905
rect 34154 6893 34160 6945
rect 34192 6893 34198 6945
rect 34250 6933 34256 6945
rect 34675 6936 34733 6942
rect 34675 6933 34687 6936
rect 34250 6905 34687 6933
rect 34250 6893 34256 6905
rect 34675 6902 34687 6905
rect 34721 6902 34733 6936
rect 34675 6896 34733 6902
rect 35536 6893 35542 6945
rect 35594 6933 35600 6945
rect 36115 6936 36173 6942
rect 36115 6933 36127 6936
rect 35594 6905 36127 6933
rect 35594 6893 35600 6905
rect 36115 6902 36127 6905
rect 36161 6902 36173 6936
rect 36115 6896 36173 6902
rect 36400 6893 36406 6945
rect 36458 6933 36464 6945
rect 36883 6936 36941 6942
rect 36883 6933 36895 6936
rect 36458 6905 36895 6933
rect 36458 6893 36464 6905
rect 36883 6902 36895 6905
rect 36929 6902 36941 6936
rect 36883 6896 36941 6902
rect 36976 6893 36982 6945
rect 37034 6933 37040 6945
rect 37651 6936 37709 6942
rect 37651 6933 37663 6936
rect 37034 6905 37663 6933
rect 37034 6893 37040 6905
rect 37651 6902 37663 6905
rect 37697 6902 37709 6936
rect 37651 6896 37709 6902
rect 37744 6893 37750 6945
rect 37802 6933 37808 6945
rect 38419 6936 38477 6942
rect 37802 6905 37847 6933
rect 37802 6893 37808 6905
rect 38419 6902 38431 6936
rect 38465 6902 38477 6936
rect 38419 6896 38477 6902
rect 30064 6819 30070 6871
rect 30122 6859 30128 6871
rect 33808 6859 33814 6871
rect 30122 6831 33814 6859
rect 30122 6819 30128 6831
rect 33808 6819 33814 6831
rect 33866 6819 33872 6871
rect 34576 6819 34582 6871
rect 34634 6859 34640 6871
rect 37264 6859 37270 6871
rect 34634 6831 37270 6859
rect 34634 6819 34640 6831
rect 37264 6819 37270 6831
rect 37322 6819 37328 6871
rect 37360 6819 37366 6871
rect 37418 6859 37424 6871
rect 38434 6859 38462 6896
rect 38512 6893 38518 6945
rect 38570 6933 38576 6945
rect 39970 6942 39998 6979
rect 41203 6976 41215 7010
rect 41249 7007 41261 7010
rect 41491 7010 41549 7016
rect 41491 7007 41503 7010
rect 41249 6979 41503 7007
rect 41249 6976 41261 6979
rect 41203 6970 41261 6976
rect 41491 6976 41503 6979
rect 41537 7007 41549 7010
rect 41584 7007 41590 7019
rect 41537 6979 41590 7007
rect 41537 6976 41549 6979
rect 41491 6970 41549 6976
rect 41584 6967 41590 6979
rect 41642 6967 41648 7019
rect 43027 7010 43085 7016
rect 43027 7007 43039 7010
rect 42946 6979 43039 7007
rect 39187 6936 39245 6942
rect 38570 6905 38615 6933
rect 38570 6893 38576 6905
rect 39187 6902 39199 6936
rect 39233 6902 39245 6936
rect 39187 6896 39245 6902
rect 39955 6936 40013 6942
rect 39955 6902 39967 6936
rect 40001 6902 40013 6936
rect 39955 6896 40013 6902
rect 40051 6936 40109 6942
rect 40051 6902 40063 6936
rect 40097 6933 40109 6936
rect 40624 6933 40630 6945
rect 40097 6905 40630 6933
rect 40097 6902 40109 6905
rect 40051 6896 40109 6902
rect 37418 6831 38462 6859
rect 37418 6819 37424 6831
rect 28586 6757 29534 6785
rect 28586 6745 28592 6757
rect 29776 6745 29782 6797
rect 29834 6785 29840 6797
rect 33232 6785 33238 6797
rect 29834 6757 33238 6785
rect 29834 6745 29840 6757
rect 33232 6745 33238 6757
rect 33290 6745 33296 6797
rect 33715 6788 33773 6794
rect 33715 6754 33727 6788
rect 33761 6785 33773 6788
rect 34096 6785 34102 6797
rect 33761 6757 34102 6785
rect 33761 6754 33773 6757
rect 33715 6748 33773 6754
rect 34096 6745 34102 6757
rect 34154 6785 34160 6797
rect 35440 6785 35446 6797
rect 34154 6757 35446 6785
rect 34154 6745 34160 6757
rect 35440 6745 35446 6757
rect 35498 6745 35504 6797
rect 37648 6745 37654 6797
rect 37706 6785 37712 6797
rect 39202 6785 39230 6896
rect 40624 6893 40630 6905
rect 40682 6893 40688 6945
rect 42064 6933 42070 6945
rect 41218 6905 42070 6933
rect 39280 6819 39286 6871
rect 39338 6859 39344 6871
rect 41218 6859 41246 6905
rect 42064 6893 42070 6905
rect 42122 6893 42128 6945
rect 42163 6936 42221 6942
rect 42163 6902 42175 6936
rect 42209 6902 42221 6936
rect 42163 6896 42221 6902
rect 39338 6831 41246 6859
rect 39338 6819 39344 6831
rect 41584 6819 41590 6871
rect 41642 6859 41648 6871
rect 42178 6859 42206 6896
rect 41642 6831 42206 6859
rect 41642 6819 41648 6831
rect 37706 6757 39230 6785
rect 37706 6745 37712 6757
rect 39376 6745 39382 6797
rect 39434 6785 39440 6797
rect 42352 6785 42358 6797
rect 39434 6757 42358 6785
rect 39434 6745 39440 6757
rect 42352 6745 42358 6757
rect 42410 6745 42416 6797
rect 42640 6745 42646 6797
rect 42698 6785 42704 6797
rect 42946 6785 42974 6979
rect 43027 6976 43039 6979
rect 43073 6976 43085 7010
rect 43027 6970 43085 6976
rect 43216 6967 43222 7019
rect 43274 7007 43280 7019
rect 43795 7010 43853 7016
rect 43795 7007 43807 7010
rect 43274 6979 43807 7007
rect 43274 6967 43280 6979
rect 43795 6976 43807 6979
rect 43841 6976 43853 7010
rect 45251 7010 45309 7016
rect 45251 7007 45263 7010
rect 43795 6970 43853 6976
rect 44290 6979 45263 7007
rect 44290 6945 44318 6979
rect 45251 6976 45263 6979
rect 45297 6976 45309 7010
rect 45251 6970 45309 6976
rect 46864 6967 46870 7019
rect 46922 7007 46928 7019
rect 46922 6979 48254 7007
rect 46922 6967 46928 6979
rect 43699 6936 43757 6942
rect 43699 6902 43711 6936
rect 43745 6902 43757 6936
rect 43699 6896 43757 6902
rect 43120 6819 43126 6871
rect 43178 6859 43184 6871
rect 43714 6859 43742 6896
rect 44272 6893 44278 6945
rect 44330 6893 44336 6945
rect 44368 6893 44374 6945
rect 44426 6933 44432 6945
rect 44563 6936 44621 6942
rect 44563 6933 44575 6936
rect 44426 6905 44575 6933
rect 44426 6893 44432 6905
rect 44563 6902 44575 6905
rect 44609 6902 44621 6936
rect 45328 6933 45334 6945
rect 45289 6905 45334 6933
rect 44563 6896 44621 6902
rect 45328 6893 45334 6905
rect 45386 6893 45392 6945
rect 46384 6893 46390 6945
rect 46442 6933 46448 6945
rect 46675 6936 46733 6942
rect 46675 6933 46687 6936
rect 46442 6905 46687 6933
rect 46442 6893 46448 6905
rect 46675 6902 46687 6905
rect 46721 6902 46733 6936
rect 46675 6896 46733 6902
rect 46771 6936 46829 6942
rect 46771 6902 46783 6936
rect 46817 6902 46829 6936
rect 46771 6896 46829 6902
rect 43178 6831 43742 6859
rect 43178 6819 43184 6831
rect 45616 6819 45622 6871
rect 45674 6859 45680 6871
rect 46786 6859 46814 6896
rect 47152 6893 47158 6945
rect 47210 6933 47216 6945
rect 48226 6942 48254 6979
rect 48496 6967 48502 7019
rect 48554 7007 48560 7019
rect 49075 7010 49133 7016
rect 49075 7007 49087 7010
rect 48554 6979 49087 7007
rect 48554 6967 48560 6979
rect 49075 6976 49087 6979
rect 49121 6976 49133 7010
rect 49075 6970 49133 6976
rect 54067 7010 54125 7016
rect 54067 6976 54079 7010
rect 54113 6976 54125 7010
rect 54736 7007 54742 7019
rect 54697 6979 54742 7007
rect 54067 6970 54125 6976
rect 47443 6936 47501 6942
rect 47443 6933 47455 6936
rect 47210 6905 47455 6933
rect 47210 6893 47216 6905
rect 47443 6902 47455 6905
rect 47489 6902 47501 6936
rect 47443 6896 47501 6902
rect 47539 6936 47597 6942
rect 47539 6902 47551 6936
rect 47585 6902 47597 6936
rect 47539 6896 47597 6902
rect 48211 6936 48269 6942
rect 48211 6902 48223 6936
rect 48257 6902 48269 6936
rect 48211 6896 48269 6902
rect 45674 6831 46814 6859
rect 45674 6819 45680 6831
rect 47056 6819 47062 6871
rect 47114 6859 47120 6871
rect 47554 6859 47582 6896
rect 48304 6893 48310 6945
rect 48362 6933 48368 6945
rect 48979 6936 49037 6942
rect 48979 6933 48991 6936
rect 48362 6905 48991 6933
rect 48362 6893 48368 6905
rect 48979 6902 48991 6905
rect 49025 6902 49037 6936
rect 48979 6896 49037 6902
rect 50323 6936 50381 6942
rect 50323 6902 50335 6936
rect 50369 6902 50381 6936
rect 50323 6896 50381 6902
rect 47114 6831 47582 6859
rect 47114 6819 47120 6831
rect 50128 6819 50134 6871
rect 50186 6859 50192 6871
rect 50338 6859 50366 6896
rect 51472 6893 51478 6945
rect 51530 6933 51536 6945
rect 52051 6936 52109 6942
rect 52051 6933 52063 6936
rect 51530 6905 52063 6933
rect 51530 6893 51536 6905
rect 52051 6902 52063 6905
rect 52097 6902 52109 6936
rect 52720 6933 52726 6945
rect 52681 6905 52726 6933
rect 52051 6896 52109 6902
rect 52720 6893 52726 6905
rect 52778 6893 52784 6945
rect 52819 6936 52877 6942
rect 52819 6902 52831 6936
rect 52865 6902 52877 6936
rect 54082 6933 54110 6970
rect 54736 6967 54742 6979
rect 54794 6967 54800 7019
rect 55408 6967 55414 7019
rect 55466 7007 55472 7019
rect 55507 7010 55565 7016
rect 55507 7007 55519 7010
rect 55466 6979 55519 7007
rect 55466 6967 55472 6979
rect 55507 6976 55519 6979
rect 55553 6976 55565 7010
rect 55507 6970 55565 6976
rect 57811 7010 57869 7016
rect 57811 6976 57823 7010
rect 57857 7007 57869 7010
rect 58480 7007 58486 7019
rect 57857 6979 58486 7007
rect 57857 6976 57869 6979
rect 57811 6970 57869 6976
rect 58480 6967 58486 6979
rect 58538 6967 58544 7019
rect 56272 6933 56278 6945
rect 54082 6905 56278 6933
rect 52819 6896 52877 6902
rect 50186 6831 50366 6859
rect 50186 6819 50192 6831
rect 50416 6819 50422 6871
rect 50474 6859 50480 6871
rect 52834 6859 52862 6896
rect 56272 6893 56278 6905
rect 56330 6893 56336 6945
rect 50474 6831 52862 6859
rect 50474 6819 50480 6831
rect 46384 6785 46390 6797
rect 42698 6757 42974 6785
rect 46345 6757 46390 6785
rect 42698 6745 42704 6757
rect 46384 6745 46390 6757
rect 46442 6745 46448 6797
rect 47152 6785 47158 6797
rect 47113 6757 47158 6785
rect 47152 6745 47158 6757
rect 47210 6745 47216 6797
rect 1152 6686 58848 6708
rect 1152 6634 4294 6686
rect 4346 6634 4358 6686
rect 4410 6634 4422 6686
rect 4474 6634 4486 6686
rect 4538 6634 35014 6686
rect 35066 6634 35078 6686
rect 35130 6634 35142 6686
rect 35194 6634 35206 6686
rect 35258 6634 58848 6686
rect 1152 6612 58848 6634
rect 6832 6563 6838 6575
rect 6793 6535 6838 6563
rect 6832 6523 6838 6535
rect 6890 6563 6896 6575
rect 6890 6535 7166 6563
rect 6890 6523 6896 6535
rect 5680 6415 5686 6427
rect 5641 6387 5686 6415
rect 5680 6375 5686 6387
rect 5738 6375 5744 6427
rect 7138 6424 7166 6535
rect 7954 6535 8270 6563
rect 7603 6492 7661 6498
rect 7603 6458 7615 6492
rect 7649 6489 7661 6492
rect 7954 6489 7982 6535
rect 7649 6461 7982 6489
rect 8242 6489 8270 6535
rect 8848 6523 8854 6575
rect 8906 6563 8912 6575
rect 10576 6563 10582 6575
rect 8906 6535 10582 6563
rect 8906 6523 8912 6535
rect 10576 6523 10582 6535
rect 10634 6523 10640 6575
rect 10960 6523 10966 6575
rect 11018 6563 11024 6575
rect 13555 6566 13613 6572
rect 13555 6563 13567 6566
rect 11018 6535 13567 6563
rect 11018 6523 11024 6535
rect 13555 6532 13567 6535
rect 13601 6563 13613 6566
rect 13840 6563 13846 6575
rect 13601 6535 13846 6563
rect 13601 6532 13613 6535
rect 13555 6526 13613 6532
rect 13840 6523 13846 6535
rect 13898 6523 13904 6575
rect 14512 6523 14518 6575
rect 14570 6563 14576 6575
rect 14570 6535 17438 6563
rect 14570 6523 14576 6535
rect 8944 6489 8950 6501
rect 8242 6461 8950 6489
rect 7649 6458 7661 6461
rect 7603 6452 7661 6458
rect 8944 6449 8950 6461
rect 9002 6449 9008 6501
rect 11152 6449 11158 6501
rect 11210 6489 11216 6501
rect 17410 6489 17438 6535
rect 17488 6523 17494 6575
rect 17546 6563 17552 6575
rect 24016 6563 24022 6575
rect 17546 6535 24022 6563
rect 17546 6523 17552 6535
rect 24016 6523 24022 6535
rect 24074 6523 24080 6575
rect 24226 6535 27806 6563
rect 18163 6492 18221 6498
rect 18163 6489 18175 6492
rect 11210 6461 16286 6489
rect 17410 6461 18175 6489
rect 11210 6449 11216 6461
rect 7123 6418 7181 6424
rect 7123 6384 7135 6418
rect 7169 6384 7181 6418
rect 8368 6415 8374 6427
rect 7123 6378 7181 6384
rect 7234 6387 7968 6415
rect 8256 6387 8374 6415
rect 1552 6341 1558 6353
rect 1513 6313 1558 6341
rect 1552 6301 1558 6313
rect 1610 6301 1616 6353
rect 2032 6301 2038 6353
rect 2090 6341 2096 6353
rect 2323 6344 2381 6350
rect 2323 6341 2335 6344
rect 2090 6313 2335 6341
rect 2090 6301 2096 6313
rect 2323 6310 2335 6313
rect 2369 6310 2381 6344
rect 3184 6341 3190 6353
rect 3145 6313 3190 6341
rect 2323 6304 2381 6310
rect 3184 6301 3190 6313
rect 3242 6301 3248 6353
rect 3856 6301 3862 6353
rect 3914 6341 3920 6353
rect 3955 6344 4013 6350
rect 3955 6341 3967 6344
rect 3914 6313 3967 6341
rect 3914 6301 3920 6313
rect 3955 6310 3967 6313
rect 4001 6310 4013 6344
rect 3955 6304 4013 6310
rect 4624 6301 4630 6353
rect 4682 6341 4688 6353
rect 4723 6344 4781 6350
rect 4723 6341 4735 6344
rect 4682 6313 4735 6341
rect 4682 6301 4688 6313
rect 4723 6310 4735 6313
rect 4769 6310 4781 6344
rect 4723 6304 4781 6310
rect 5104 6301 5110 6353
rect 5162 6341 5168 6353
rect 7234 6341 7262 6387
rect 8368 6375 8374 6387
rect 8426 6375 8432 6427
rect 9616 6375 9622 6427
rect 9674 6415 9680 6427
rect 9674 6387 13790 6415
rect 9674 6375 9680 6387
rect 9424 6341 9430 6353
rect 5162 6313 7262 6341
rect 9385 6313 9430 6341
rect 5162 6301 5168 6313
rect 9424 6301 9430 6313
rect 9482 6301 9488 6353
rect 10096 6301 10102 6353
rect 10154 6341 10160 6353
rect 10195 6344 10253 6350
rect 10195 6341 10207 6344
rect 10154 6313 10207 6341
rect 10154 6301 10160 6313
rect 10195 6310 10207 6313
rect 10241 6310 10253 6344
rect 10195 6304 10253 6310
rect 10864 6301 10870 6353
rect 10922 6341 10928 6353
rect 10963 6344 11021 6350
rect 10963 6341 10975 6344
rect 10922 6313 10975 6341
rect 10922 6301 10928 6313
rect 10963 6310 10975 6313
rect 11009 6310 11021 6344
rect 10963 6304 11021 6310
rect 11632 6301 11638 6353
rect 11690 6341 11696 6353
rect 12211 6344 12269 6350
rect 12211 6341 12223 6344
rect 11690 6313 12223 6341
rect 11690 6301 11696 6313
rect 12211 6310 12223 6313
rect 12257 6310 12269 6344
rect 12211 6304 12269 6310
rect 12304 6301 12310 6353
rect 12362 6341 12368 6353
rect 13075 6344 13133 6350
rect 13075 6341 13087 6344
rect 12362 6313 13087 6341
rect 12362 6301 12368 6313
rect 13075 6310 13087 6313
rect 13121 6310 13133 6344
rect 13762 6341 13790 6387
rect 13840 6375 13846 6427
rect 13898 6415 13904 6427
rect 14704 6415 14710 6427
rect 13898 6387 13943 6415
rect 14665 6387 14710 6415
rect 13898 6375 13904 6387
rect 14704 6375 14710 6387
rect 14762 6375 14768 6427
rect 15088 6415 15094 6427
rect 15049 6387 15094 6415
rect 15088 6375 15094 6387
rect 15146 6415 15152 6427
rect 16258 6424 16286 6461
rect 18163 6458 18175 6461
rect 18209 6458 18221 6492
rect 18163 6452 18221 6458
rect 18274 6461 18974 6489
rect 15475 6418 15533 6424
rect 15475 6415 15487 6418
rect 15146 6387 15487 6415
rect 15146 6375 15152 6387
rect 15475 6384 15487 6387
rect 15521 6384 15533 6418
rect 15475 6378 15533 6384
rect 16243 6418 16301 6424
rect 16243 6384 16255 6418
rect 16289 6384 16301 6418
rect 16243 6378 16301 6384
rect 16720 6375 16726 6427
rect 16778 6415 16784 6427
rect 17587 6418 17645 6424
rect 17587 6415 17599 6418
rect 16778 6387 17599 6415
rect 16778 6375 16784 6387
rect 17587 6384 17599 6387
rect 17633 6384 17645 6418
rect 17587 6378 17645 6384
rect 17680 6375 17686 6427
rect 17738 6415 17744 6427
rect 18274 6415 18302 6461
rect 18448 6415 18454 6427
rect 17738 6387 18302 6415
rect 18409 6387 18454 6415
rect 17738 6375 17744 6387
rect 18448 6375 18454 6387
rect 18506 6375 18512 6427
rect 18946 6415 18974 6461
rect 19024 6449 19030 6501
rect 19082 6489 19088 6501
rect 24226 6489 24254 6535
rect 19082 6461 24254 6489
rect 19082 6449 19088 6461
rect 25168 6449 25174 6501
rect 25226 6489 25232 6501
rect 27664 6489 27670 6501
rect 25226 6461 27670 6489
rect 25226 6449 25232 6461
rect 27664 6449 27670 6461
rect 27722 6449 27728 6501
rect 27778 6498 27806 6535
rect 27952 6523 27958 6575
rect 28010 6563 28016 6575
rect 28624 6563 28630 6575
rect 28010 6535 28630 6563
rect 28010 6523 28016 6535
rect 28624 6523 28630 6535
rect 28682 6523 28688 6575
rect 28723 6566 28781 6572
rect 28723 6532 28735 6566
rect 28769 6563 28781 6566
rect 28816 6563 28822 6575
rect 28769 6535 28822 6563
rect 28769 6532 28781 6535
rect 28723 6526 28781 6532
rect 28816 6523 28822 6535
rect 28874 6523 28880 6575
rect 29104 6523 29110 6575
rect 29162 6563 29168 6575
rect 32272 6563 32278 6575
rect 29162 6535 32278 6563
rect 29162 6523 29168 6535
rect 32272 6523 32278 6535
rect 32330 6523 32336 6575
rect 32386 6535 32606 6563
rect 27763 6492 27821 6498
rect 27763 6458 27775 6492
rect 27809 6458 27821 6492
rect 27763 6452 27821 6458
rect 28435 6492 28493 6498
rect 28435 6458 28447 6492
rect 28481 6489 28493 6492
rect 32386 6489 32414 6535
rect 28481 6461 32414 6489
rect 32578 6489 32606 6535
rect 33520 6523 33526 6575
rect 33578 6563 33584 6575
rect 36883 6566 36941 6572
rect 36883 6563 36895 6566
rect 33578 6535 36895 6563
rect 33578 6523 33584 6535
rect 36883 6532 36895 6535
rect 36929 6563 36941 6566
rect 36929 6535 37214 6563
rect 36929 6532 36941 6535
rect 36883 6526 36941 6532
rect 36211 6492 36269 6498
rect 36211 6489 36223 6492
rect 32578 6461 36223 6489
rect 28481 6458 28493 6461
rect 28435 6452 28493 6458
rect 36211 6458 36223 6461
rect 36257 6458 36269 6492
rect 36211 6452 36269 6458
rect 19600 6415 19606 6427
rect 18946 6387 19606 6415
rect 19600 6375 19606 6387
rect 19658 6375 19664 6427
rect 19699 6418 19757 6424
rect 19699 6384 19711 6418
rect 19745 6415 19757 6418
rect 19984 6415 19990 6427
rect 19745 6387 19990 6415
rect 19745 6384 19757 6387
rect 19699 6378 19757 6384
rect 19984 6375 19990 6387
rect 20042 6375 20048 6427
rect 20080 6375 20086 6427
rect 20138 6415 20144 6427
rect 24496 6415 24502 6427
rect 20138 6387 21182 6415
rect 24457 6387 24502 6415
rect 20138 6375 20144 6387
rect 17296 6341 17302 6353
rect 13762 6313 17302 6341
rect 13075 6304 13133 6310
rect 17296 6301 17302 6313
rect 17354 6301 17360 6353
rect 19219 6344 19277 6350
rect 19219 6341 19231 6344
rect 17410 6313 19231 6341
rect 9040 6227 9046 6279
rect 9098 6267 9104 6279
rect 12976 6267 12982 6279
rect 9098 6239 12982 6267
rect 9098 6227 9104 6239
rect 12976 6227 12982 6239
rect 13034 6227 13040 6279
rect 17410 6267 17438 6313
rect 19219 6310 19231 6313
rect 19265 6310 19277 6344
rect 19219 6304 19277 6310
rect 19312 6301 19318 6353
rect 19370 6341 19376 6353
rect 20675 6344 20733 6350
rect 20675 6341 20687 6344
rect 19370 6313 20687 6341
rect 19370 6301 19376 6313
rect 20675 6310 20687 6313
rect 20721 6310 20733 6344
rect 21154 6341 21182 6387
rect 24496 6375 24502 6387
rect 24554 6375 24560 6427
rect 27955 6418 28013 6424
rect 27955 6384 27967 6418
rect 28001 6415 28013 6418
rect 28240 6415 28246 6427
rect 28001 6387 28246 6415
rect 28001 6384 28013 6387
rect 27955 6378 28013 6384
rect 28240 6375 28246 6387
rect 28298 6375 28304 6427
rect 29008 6415 29014 6427
rect 28969 6387 29014 6415
rect 29008 6375 29014 6387
rect 29066 6375 29072 6427
rect 30355 6418 30413 6424
rect 30355 6384 30367 6418
rect 30401 6415 30413 6418
rect 30640 6415 30646 6427
rect 30401 6387 30646 6415
rect 30401 6384 30413 6387
rect 30355 6378 30413 6384
rect 30640 6375 30646 6387
rect 30698 6375 30704 6427
rect 30736 6375 30742 6427
rect 30794 6415 30800 6427
rect 31891 6418 31949 6424
rect 30794 6387 31358 6415
rect 30794 6375 30800 6387
rect 25648 6341 25654 6353
rect 21154 6313 25502 6341
rect 25609 6313 25654 6341
rect 20675 6304 20733 6310
rect 13186 6239 17438 6267
rect 17683 6270 17741 6276
rect 8752 6153 8758 6205
rect 8810 6193 8816 6205
rect 13072 6193 13078 6205
rect 8810 6165 13078 6193
rect 8810 6153 8816 6165
rect 13072 6153 13078 6165
rect 13130 6153 13136 6205
rect 5488 6079 5494 6131
rect 5546 6119 5552 6131
rect 5587 6122 5645 6128
rect 5587 6119 5599 6122
rect 5546 6091 5599 6119
rect 5546 6079 5552 6091
rect 5587 6088 5599 6091
rect 5633 6088 5645 6122
rect 5587 6082 5645 6088
rect 6256 6079 6262 6131
rect 6314 6119 6320 6131
rect 7027 6122 7085 6128
rect 7027 6119 7039 6122
rect 6314 6091 7039 6119
rect 6314 6079 6320 6091
rect 7027 6088 7039 6091
rect 7073 6088 7085 6122
rect 7027 6082 7085 6088
rect 9232 6079 9238 6131
rect 9290 6119 9296 6131
rect 13186 6119 13214 6239
rect 17683 6236 17695 6270
rect 17729 6236 17741 6270
rect 17683 6230 17741 6236
rect 18163 6270 18221 6276
rect 18163 6236 18175 6270
rect 18209 6267 18221 6270
rect 20464 6267 20470 6279
rect 18209 6239 20470 6267
rect 18209 6236 18221 6239
rect 18163 6230 18221 6236
rect 14896 6153 14902 6205
rect 14954 6193 14960 6205
rect 17395 6196 17453 6202
rect 14954 6165 16190 6193
rect 14954 6153 14960 6165
rect 9290 6091 13214 6119
rect 9290 6079 9296 6091
rect 13264 6079 13270 6131
rect 13322 6119 13328 6131
rect 13939 6122 13997 6128
rect 13939 6119 13951 6122
rect 13322 6091 13951 6119
rect 13322 6079 13328 6091
rect 13939 6088 13951 6091
rect 13985 6088 13997 6122
rect 13939 6082 13997 6088
rect 14512 6079 14518 6131
rect 14570 6119 14576 6131
rect 14611 6122 14669 6128
rect 14611 6119 14623 6122
rect 14570 6091 14623 6119
rect 14570 6079 14576 6091
rect 14611 6088 14623 6091
rect 14657 6088 14669 6122
rect 14611 6082 14669 6088
rect 14704 6079 14710 6131
rect 14762 6119 14768 6131
rect 16162 6128 16190 6165
rect 17395 6162 17407 6196
rect 17441 6193 17453 6196
rect 17698 6193 17726 6230
rect 20464 6227 20470 6239
rect 20522 6227 20528 6279
rect 20560 6227 20566 6279
rect 20618 6267 20624 6279
rect 20755 6270 20813 6276
rect 20755 6267 20767 6270
rect 20618 6239 20767 6267
rect 20618 6227 20624 6239
rect 20755 6236 20767 6239
rect 20801 6236 20813 6270
rect 20755 6230 20813 6236
rect 21523 6270 21581 6276
rect 21523 6236 21535 6270
rect 21569 6267 21581 6270
rect 22768 6267 22774 6279
rect 21569 6239 22774 6267
rect 21569 6236 21581 6239
rect 21523 6230 21581 6236
rect 22768 6227 22774 6239
rect 22826 6227 22832 6279
rect 22960 6267 22966 6279
rect 22921 6239 22966 6267
rect 22960 6227 22966 6239
rect 23018 6227 23024 6279
rect 23731 6270 23789 6276
rect 23731 6236 23743 6270
rect 23777 6267 23789 6270
rect 24400 6267 24406 6279
rect 23777 6239 24406 6267
rect 23777 6236 23789 6239
rect 23731 6230 23789 6236
rect 24400 6227 24406 6239
rect 24458 6227 24464 6279
rect 25474 6267 25502 6313
rect 25648 6301 25654 6313
rect 25706 6301 25712 6353
rect 26800 6341 26806 6353
rect 26761 6313 26806 6341
rect 26800 6301 26806 6313
rect 26858 6301 26864 6353
rect 27763 6344 27821 6350
rect 27763 6310 27775 6344
rect 27809 6341 27821 6344
rect 29680 6341 29686 6353
rect 27809 6313 29342 6341
rect 29641 6313 29686 6341
rect 27809 6310 27821 6313
rect 27763 6304 27821 6310
rect 28435 6270 28493 6276
rect 28435 6267 28447 6270
rect 25474 6239 28447 6267
rect 28435 6236 28447 6239
rect 28481 6236 28493 6270
rect 28435 6230 28493 6236
rect 29314 6193 29342 6313
rect 29680 6301 29686 6313
rect 29738 6301 29744 6353
rect 31216 6341 31222 6353
rect 31177 6313 31222 6341
rect 31216 6301 31222 6313
rect 31274 6301 31280 6353
rect 31330 6341 31358 6387
rect 31891 6384 31903 6418
rect 31937 6415 31949 6418
rect 32080 6415 32086 6427
rect 31937 6387 32086 6415
rect 31937 6384 31949 6387
rect 31891 6378 31949 6384
rect 32080 6375 32086 6387
rect 32138 6415 32144 6427
rect 32371 6418 32429 6424
rect 32371 6415 32383 6418
rect 32138 6387 32383 6415
rect 32138 6375 32144 6387
rect 32371 6384 32383 6387
rect 32417 6384 32429 6418
rect 34288 6415 34294 6427
rect 34249 6387 34294 6415
rect 32371 6378 32429 6384
rect 34288 6375 34294 6387
rect 34346 6375 34352 6427
rect 34672 6415 34678 6427
rect 34633 6387 34678 6415
rect 34672 6375 34678 6387
rect 34730 6415 34736 6427
rect 37186 6424 37214 6535
rect 38512 6523 38518 6575
rect 38570 6563 38576 6575
rect 41200 6563 41206 6575
rect 38570 6535 41206 6563
rect 38570 6523 38576 6535
rect 41200 6523 41206 6535
rect 41258 6523 41264 6575
rect 43216 6563 43222 6575
rect 42082 6535 43222 6563
rect 37264 6449 37270 6501
rect 37322 6489 37328 6501
rect 42082 6489 42110 6535
rect 43216 6523 43222 6535
rect 43274 6523 43280 6575
rect 44560 6563 44566 6575
rect 44521 6535 44566 6563
rect 44560 6523 44566 6535
rect 44618 6523 44624 6575
rect 46576 6563 46582 6575
rect 44866 6535 46582 6563
rect 37322 6461 42110 6489
rect 37322 6449 37328 6461
rect 42256 6449 42262 6501
rect 42314 6489 42320 6501
rect 44866 6489 44894 6535
rect 46576 6523 46582 6535
rect 46634 6523 46640 6575
rect 51280 6563 51286 6575
rect 51241 6535 51286 6563
rect 51280 6523 51286 6535
rect 51338 6563 51344 6575
rect 51338 6535 51614 6563
rect 51338 6523 51344 6535
rect 42314 6461 44894 6489
rect 42314 6449 42320 6461
rect 44944 6449 44950 6501
rect 45002 6489 45008 6501
rect 45002 6461 50942 6489
rect 45002 6449 45008 6461
rect 34963 6418 35021 6424
rect 34963 6415 34975 6418
rect 34730 6387 34975 6415
rect 34730 6375 34736 6387
rect 34963 6384 34975 6387
rect 35009 6384 35021 6418
rect 34963 6378 35021 6384
rect 36019 6418 36077 6424
rect 36019 6384 36031 6418
rect 36065 6415 36077 6418
rect 37171 6418 37229 6424
rect 36065 6387 36446 6415
rect 36065 6384 36077 6387
rect 36019 6378 36077 6384
rect 32755 6344 32813 6350
rect 32755 6341 32767 6344
rect 31330 6313 32767 6341
rect 32755 6310 32767 6313
rect 32801 6310 32813 6344
rect 36304 6341 36310 6353
rect 32755 6304 32813 6310
rect 33106 6313 36158 6341
rect 36265 6313 36310 6341
rect 29587 6270 29645 6276
rect 29587 6236 29599 6270
rect 29633 6267 29645 6270
rect 33106 6267 33134 6313
rect 29633 6239 33134 6267
rect 33235 6270 33293 6276
rect 29633 6236 29645 6239
rect 29587 6230 29645 6236
rect 33235 6236 33247 6270
rect 33281 6267 33293 6270
rect 33427 6270 33485 6276
rect 33427 6267 33439 6270
rect 33281 6239 33439 6267
rect 33281 6236 33293 6239
rect 33235 6230 33293 6236
rect 33427 6236 33439 6239
rect 33473 6267 33485 6270
rect 33715 6270 33773 6276
rect 33715 6267 33727 6270
rect 33473 6239 33727 6267
rect 33473 6236 33485 6239
rect 33427 6230 33485 6236
rect 33715 6236 33727 6239
rect 33761 6236 33773 6270
rect 36019 6270 36077 6276
rect 36019 6267 36031 6270
rect 33715 6230 33773 6236
rect 33826 6239 36031 6267
rect 33136 6193 33142 6205
rect 17441 6165 20030 6193
rect 17441 6162 17453 6165
rect 17395 6156 17453 6162
rect 15379 6122 15437 6128
rect 15379 6119 15391 6122
rect 14762 6091 15391 6119
rect 14762 6079 14768 6091
rect 15379 6088 15391 6091
rect 15425 6088 15437 6122
rect 15379 6082 15437 6088
rect 16147 6122 16205 6128
rect 16147 6088 16159 6122
rect 16193 6088 16205 6122
rect 16147 6082 16205 6088
rect 17488 6079 17494 6131
rect 17546 6119 17552 6131
rect 18355 6122 18413 6128
rect 18355 6119 18367 6122
rect 17546 6091 18367 6119
rect 17546 6079 17552 6091
rect 18355 6088 18367 6091
rect 18401 6088 18413 6122
rect 18355 6082 18413 6088
rect 18448 6079 18454 6131
rect 18506 6119 18512 6131
rect 19123 6122 19181 6128
rect 19123 6119 19135 6122
rect 18506 6091 19135 6119
rect 18506 6079 18512 6091
rect 19123 6088 19135 6091
rect 19169 6088 19181 6122
rect 19123 6082 19181 6088
rect 19504 6079 19510 6131
rect 19562 6119 19568 6131
rect 19891 6122 19949 6128
rect 19891 6119 19903 6122
rect 19562 6091 19903 6119
rect 19562 6079 19568 6091
rect 19891 6088 19903 6091
rect 19937 6088 19949 6122
rect 20002 6119 20030 6165
rect 20674 6165 29054 6193
rect 29314 6165 33142 6193
rect 20674 6119 20702 6165
rect 21424 6119 21430 6131
rect 20002 6091 20702 6119
rect 21385 6091 21430 6119
rect 19891 6082 19949 6088
rect 21424 6079 21430 6091
rect 21482 6079 21488 6131
rect 21520 6079 21526 6131
rect 21578 6119 21584 6131
rect 22867 6122 22925 6128
rect 22867 6119 22879 6122
rect 21578 6091 22879 6119
rect 21578 6079 21584 6091
rect 22867 6088 22879 6091
rect 22913 6088 22925 6122
rect 22867 6082 22925 6088
rect 22960 6079 22966 6131
rect 23018 6119 23024 6131
rect 23635 6122 23693 6128
rect 23635 6119 23647 6122
rect 23018 6091 23647 6119
rect 23018 6079 23024 6091
rect 23635 6088 23647 6091
rect 23681 6088 23693 6122
rect 23635 6082 23693 6088
rect 24304 6079 24310 6131
rect 24362 6119 24368 6131
rect 24403 6122 24461 6128
rect 24403 6119 24415 6122
rect 24362 6091 24415 6119
rect 24362 6079 24368 6091
rect 24403 6088 24415 6091
rect 24449 6088 24461 6122
rect 24403 6082 24461 6088
rect 27568 6079 27574 6131
rect 27626 6119 27632 6131
rect 28147 6122 28205 6128
rect 28147 6119 28159 6122
rect 27626 6091 28159 6119
rect 27626 6079 27632 6091
rect 28147 6088 28159 6091
rect 28193 6088 28205 6122
rect 28147 6082 28205 6088
rect 28432 6079 28438 6131
rect 28490 6119 28496 6131
rect 28915 6122 28973 6128
rect 28915 6119 28927 6122
rect 28490 6091 28927 6119
rect 28490 6079 28496 6091
rect 28915 6088 28927 6091
rect 28961 6088 28973 6122
rect 29026 6119 29054 6165
rect 33136 6153 33142 6165
rect 33194 6153 33200 6205
rect 29587 6122 29645 6128
rect 29587 6119 29599 6122
rect 29026 6091 29599 6119
rect 28915 6082 28973 6088
rect 29587 6088 29599 6091
rect 29633 6088 29645 6122
rect 29587 6082 29645 6088
rect 29776 6079 29782 6131
rect 29834 6119 29840 6131
rect 30547 6122 30605 6128
rect 30547 6119 30559 6122
rect 29834 6091 30559 6119
rect 29834 6079 29840 6091
rect 30547 6088 30559 6091
rect 30593 6088 30605 6122
rect 30547 6082 30605 6088
rect 30640 6079 30646 6131
rect 30698 6119 30704 6131
rect 32179 6122 32237 6128
rect 32179 6119 32191 6122
rect 30698 6091 32191 6119
rect 30698 6079 30704 6091
rect 32179 6088 32191 6091
rect 32225 6088 32237 6122
rect 32179 6082 32237 6088
rect 32755 6122 32813 6128
rect 32755 6088 32767 6122
rect 32801 6119 32813 6122
rect 33250 6119 33278 6230
rect 33328 6153 33334 6205
rect 33386 6193 33392 6205
rect 33826 6193 33854 6239
rect 36019 6236 36031 6239
rect 36065 6236 36077 6270
rect 36019 6230 36077 6236
rect 33386 6165 33854 6193
rect 33386 6153 33392 6165
rect 34480 6153 34486 6205
rect 34538 6193 34544 6205
rect 35920 6193 35926 6205
rect 34538 6165 35926 6193
rect 34538 6153 34544 6165
rect 35920 6153 35926 6165
rect 35978 6153 35984 6205
rect 36130 6193 36158 6313
rect 36304 6301 36310 6313
rect 36362 6301 36368 6353
rect 36418 6341 36446 6387
rect 37171 6384 37183 6418
rect 37217 6384 37229 6418
rect 39472 6415 39478 6427
rect 37171 6378 37229 6384
rect 37282 6387 39478 6415
rect 37282 6341 37310 6387
rect 39472 6375 39478 6387
rect 39530 6375 39536 6427
rect 41296 6415 41302 6427
rect 41257 6387 41302 6415
rect 41296 6375 41302 6387
rect 41354 6375 41360 6427
rect 42640 6415 42646 6427
rect 41410 6387 42646 6415
rect 38896 6341 38902 6353
rect 36418 6313 37310 6341
rect 38857 6313 38902 6341
rect 38896 6301 38902 6313
rect 38954 6301 38960 6353
rect 40336 6341 40342 6353
rect 40297 6313 40342 6341
rect 40336 6301 40342 6313
rect 40394 6301 40400 6353
rect 41410 6341 41438 6387
rect 42640 6375 42646 6387
rect 42698 6375 42704 6427
rect 44083 6418 44141 6424
rect 44083 6384 44095 6418
rect 44129 6415 44141 6418
rect 44176 6415 44182 6427
rect 44129 6387 44182 6415
rect 44129 6384 44141 6387
rect 44083 6378 44141 6384
rect 44176 6375 44182 6387
rect 44234 6375 44240 6427
rect 44560 6375 44566 6427
rect 44618 6415 44624 6427
rect 44755 6418 44813 6424
rect 44755 6415 44767 6418
rect 44618 6387 44767 6415
rect 44618 6375 44624 6387
rect 44755 6384 44767 6387
rect 44801 6384 44813 6418
rect 50416 6415 50422 6427
rect 44755 6378 44813 6384
rect 45346 6387 50422 6415
rect 41872 6341 41878 6353
rect 40546 6313 41438 6341
rect 41833 6313 41878 6341
rect 36211 6270 36269 6276
rect 36211 6236 36223 6270
rect 36257 6267 36269 6270
rect 40546 6267 40574 6313
rect 41872 6301 41878 6313
rect 41930 6301 41936 6353
rect 45346 6341 45374 6387
rect 50416 6375 50422 6387
rect 50474 6375 50480 6427
rect 50914 6424 50942 6461
rect 51586 6424 51614 6535
rect 50899 6418 50957 6424
rect 50899 6384 50911 6418
rect 50945 6384 50957 6418
rect 50899 6378 50957 6384
rect 51571 6418 51629 6424
rect 51571 6384 51583 6418
rect 51617 6384 51629 6418
rect 51571 6378 51629 6384
rect 52147 6418 52205 6424
rect 52147 6384 52159 6418
rect 52193 6415 52205 6418
rect 52240 6415 52246 6427
rect 52193 6387 52246 6415
rect 52193 6384 52205 6387
rect 52147 6378 52205 6384
rect 52240 6375 52246 6387
rect 52298 6415 52304 6427
rect 52339 6418 52397 6424
rect 52339 6415 52351 6418
rect 52298 6387 52351 6415
rect 52298 6375 52304 6387
rect 52339 6384 52351 6387
rect 52385 6384 52397 6418
rect 56368 6415 56374 6427
rect 52339 6378 52397 6384
rect 53314 6387 56374 6415
rect 45520 6341 45526 6353
rect 42274 6313 45374 6341
rect 45481 6313 45526 6341
rect 36257 6239 40574 6267
rect 36257 6236 36269 6239
rect 36211 6230 36269 6236
rect 40624 6227 40630 6279
rect 40682 6267 40688 6279
rect 41296 6267 41302 6279
rect 40682 6239 41302 6267
rect 40682 6227 40688 6239
rect 41296 6227 41302 6239
rect 41354 6227 41360 6279
rect 41488 6227 41494 6279
rect 41546 6267 41552 6279
rect 42274 6267 42302 6313
rect 45520 6301 45526 6313
rect 45578 6301 45584 6353
rect 46960 6341 46966 6353
rect 46921 6313 46966 6341
rect 46960 6301 46966 6313
rect 47018 6301 47024 6353
rect 47728 6341 47734 6353
rect 47689 6313 47734 6341
rect 47728 6301 47734 6313
rect 47786 6301 47792 6353
rect 48784 6301 48790 6353
rect 48842 6341 48848 6353
rect 49171 6344 49229 6350
rect 49171 6341 49183 6344
rect 48842 6313 49183 6341
rect 48842 6301 48848 6313
rect 49171 6310 49183 6313
rect 49217 6310 49229 6344
rect 49171 6304 49229 6310
rect 49552 6301 49558 6353
rect 49610 6341 49616 6353
rect 53314 6350 53342 6387
rect 56368 6375 56374 6387
rect 56426 6375 56432 6427
rect 49939 6344 49997 6350
rect 49939 6341 49951 6344
rect 49610 6313 49951 6341
rect 49610 6301 49616 6313
rect 49939 6310 49951 6313
rect 49985 6310 49997 6344
rect 49939 6304 49997 6310
rect 53299 6344 53357 6350
rect 53299 6310 53311 6344
rect 53345 6310 53357 6344
rect 53299 6304 53357 6310
rect 53968 6301 53974 6353
rect 54026 6341 54032 6353
rect 54451 6344 54509 6350
rect 54451 6341 54463 6344
rect 54026 6313 54463 6341
rect 54026 6301 54032 6313
rect 54451 6310 54463 6313
rect 54497 6310 54509 6344
rect 54451 6304 54509 6310
rect 55219 6344 55277 6350
rect 55219 6310 55231 6344
rect 55265 6310 55277 6344
rect 55219 6304 55277 6310
rect 55987 6344 56045 6350
rect 55987 6310 55999 6344
rect 56033 6310 56045 6344
rect 55987 6304 56045 6310
rect 57043 6344 57101 6350
rect 57043 6310 57055 6344
rect 57089 6310 57101 6344
rect 57043 6304 57101 6310
rect 57811 6344 57869 6350
rect 57811 6310 57823 6344
rect 57857 6341 57869 6344
rect 58096 6341 58102 6353
rect 57857 6313 58102 6341
rect 57857 6310 57869 6313
rect 57811 6304 57869 6310
rect 41546 6239 42302 6267
rect 41546 6227 41552 6239
rect 42352 6227 42358 6279
rect 42410 6267 42416 6279
rect 42451 6270 42509 6276
rect 42451 6267 42463 6270
rect 42410 6239 42463 6267
rect 42410 6227 42416 6239
rect 42451 6236 42463 6239
rect 42497 6267 42509 6270
rect 42739 6270 42797 6276
rect 42739 6267 42751 6270
rect 42497 6239 42751 6267
rect 42497 6236 42509 6239
rect 42451 6230 42509 6236
rect 42739 6236 42751 6239
rect 42785 6236 42797 6270
rect 43696 6267 43702 6279
rect 43657 6239 43702 6267
rect 42739 6230 42797 6236
rect 43696 6227 43702 6239
rect 43754 6267 43760 6279
rect 43987 6270 44045 6276
rect 43987 6267 43999 6270
rect 43754 6239 43999 6267
rect 43754 6227 43760 6239
rect 43987 6236 43999 6239
rect 44033 6236 44045 6270
rect 43987 6230 44045 6236
rect 46291 6270 46349 6276
rect 46291 6236 46303 6270
rect 46337 6236 46349 6270
rect 52240 6267 52246 6279
rect 46291 6230 46349 6236
rect 50386 6239 52246 6267
rect 46099 6196 46157 6202
rect 46099 6193 46111 6196
rect 36130 6165 37406 6193
rect 32801 6091 33278 6119
rect 32801 6088 32813 6091
rect 32755 6082 32813 6088
rect 33424 6079 33430 6131
rect 33482 6119 33488 6131
rect 33523 6122 33581 6128
rect 33523 6119 33535 6122
rect 33482 6091 33535 6119
rect 33482 6079 33488 6091
rect 33523 6088 33535 6091
rect 33569 6088 33581 6122
rect 33523 6082 33581 6088
rect 33712 6079 33718 6131
rect 33770 6119 33776 6131
rect 34195 6122 34253 6128
rect 34195 6119 34207 6122
rect 33770 6091 34207 6119
rect 33770 6079 33776 6091
rect 34195 6088 34207 6091
rect 34241 6088 34253 6122
rect 34195 6082 34253 6088
rect 34288 6079 34294 6131
rect 34346 6119 34352 6131
rect 35059 6122 35117 6128
rect 35059 6119 35071 6122
rect 34346 6091 35071 6119
rect 34346 6079 34352 6091
rect 35059 6088 35071 6091
rect 35105 6088 35117 6122
rect 35059 6082 35117 6088
rect 35440 6079 35446 6131
rect 35498 6119 35504 6131
rect 37267 6122 37325 6128
rect 37267 6119 37279 6122
rect 35498 6091 37279 6119
rect 35498 6079 35504 6091
rect 37267 6088 37279 6091
rect 37313 6088 37325 6122
rect 37378 6119 37406 6165
rect 39106 6165 46111 6193
rect 39106 6119 39134 6165
rect 46099 6162 46111 6165
rect 46145 6193 46157 6196
rect 46306 6193 46334 6230
rect 46145 6165 46334 6193
rect 46145 6162 46157 6165
rect 46099 6156 46157 6162
rect 46576 6153 46582 6205
rect 46634 6193 46640 6205
rect 50386 6193 50414 6239
rect 52240 6227 52246 6239
rect 52298 6227 52304 6279
rect 54352 6227 54358 6279
rect 54410 6267 54416 6279
rect 55234 6267 55262 6304
rect 54410 6239 55262 6267
rect 54410 6227 54416 6239
rect 46634 6165 50414 6193
rect 46634 6153 46640 6165
rect 51568 6153 51574 6205
rect 51626 6193 51632 6205
rect 51626 6165 52478 6193
rect 51626 6153 51632 6165
rect 37378 6091 39134 6119
rect 37267 6082 37325 6088
rect 39184 6079 39190 6131
rect 39242 6119 39248 6131
rect 41203 6122 41261 6128
rect 41203 6119 41215 6122
rect 39242 6091 41215 6119
rect 39242 6079 39248 6091
rect 41203 6088 41215 6091
rect 41249 6088 41261 6122
rect 41203 6082 41261 6088
rect 41296 6079 41302 6131
rect 41354 6119 41360 6131
rect 42835 6122 42893 6128
rect 42835 6119 42847 6122
rect 41354 6091 42847 6119
rect 41354 6079 41360 6091
rect 42835 6088 42847 6091
rect 42881 6088 42893 6122
rect 42835 6082 42893 6088
rect 43984 6079 43990 6131
rect 44042 6119 44048 6131
rect 44851 6122 44909 6128
rect 44851 6119 44863 6122
rect 44042 6091 44863 6119
rect 44042 6079 44048 6091
rect 44851 6088 44863 6091
rect 44897 6088 44909 6122
rect 44851 6082 44909 6088
rect 49840 6079 49846 6131
rect 49898 6119 49904 6131
rect 50803 6122 50861 6128
rect 50803 6119 50815 6122
rect 49898 6091 50815 6119
rect 49898 6079 49904 6091
rect 50803 6088 50815 6091
rect 50849 6088 50861 6122
rect 50803 6082 50861 6088
rect 51088 6079 51094 6131
rect 51146 6119 51152 6131
rect 52450 6128 52478 6165
rect 55120 6153 55126 6205
rect 55178 6193 55184 6205
rect 56002 6193 56030 6304
rect 57058 6267 57086 6304
rect 58096 6301 58102 6313
rect 58154 6301 58160 6353
rect 58864 6267 58870 6279
rect 57058 6239 58870 6267
rect 58864 6227 58870 6239
rect 58922 6227 58928 6279
rect 55178 6165 56030 6193
rect 55178 6153 55184 6165
rect 51667 6122 51725 6128
rect 51667 6119 51679 6122
rect 51146 6091 51679 6119
rect 51146 6079 51152 6091
rect 51667 6088 51679 6091
rect 51713 6088 51725 6122
rect 51667 6082 51725 6088
rect 52435 6122 52493 6128
rect 52435 6088 52447 6122
rect 52481 6088 52493 6122
rect 52435 6082 52493 6088
rect 1152 6020 58848 6042
rect 1152 5968 19654 6020
rect 19706 5968 19718 6020
rect 19770 5968 19782 6020
rect 19834 5968 19846 6020
rect 19898 5968 50374 6020
rect 50426 5968 50438 6020
rect 50490 5968 50502 6020
rect 50554 5968 50566 6020
rect 50618 5968 58848 6020
rect 1152 5946 58848 5968
rect 5200 5857 5206 5909
rect 5258 5897 5264 5909
rect 42736 5897 42742 5909
rect 5258 5869 42742 5897
rect 5258 5857 5264 5869
rect 42736 5857 42742 5869
rect 42794 5857 42800 5909
rect 43312 5857 43318 5909
rect 43370 5897 43376 5909
rect 47152 5897 47158 5909
rect 43370 5869 47158 5897
rect 43370 5857 43376 5869
rect 47152 5857 47158 5869
rect 47210 5857 47216 5909
rect 55024 5897 55030 5909
rect 54985 5869 55030 5897
rect 55024 5857 55030 5869
rect 55082 5897 55088 5909
rect 55411 5900 55469 5906
rect 55411 5897 55423 5900
rect 55082 5869 55423 5897
rect 55082 5857 55088 5869
rect 55411 5866 55423 5869
rect 55457 5866 55469 5900
rect 55411 5860 55469 5866
rect 7600 5783 7606 5835
rect 7658 5823 7664 5835
rect 20560 5823 20566 5835
rect 7658 5795 13310 5823
rect 7658 5783 7664 5795
rect 5779 5752 5837 5758
rect 5779 5718 5791 5752
rect 5825 5749 5837 5752
rect 6067 5752 6125 5758
rect 6067 5749 6079 5752
rect 5825 5721 6079 5749
rect 5825 5718 5837 5721
rect 5779 5712 5837 5718
rect 6067 5718 6079 5721
rect 6113 5749 6125 5752
rect 12016 5749 12022 5761
rect 6113 5721 12022 5749
rect 6113 5718 6125 5721
rect 6067 5712 6125 5718
rect 12016 5709 12022 5721
rect 12074 5709 12080 5761
rect 13282 5749 13310 5795
rect 14338 5795 20566 5823
rect 14224 5749 14230 5761
rect 13282 5721 14230 5749
rect 14224 5709 14230 5721
rect 14282 5709 14288 5761
rect 1072 5635 1078 5687
rect 1130 5675 1136 5687
rect 1555 5678 1613 5684
rect 1555 5675 1567 5678
rect 1130 5647 1567 5675
rect 1130 5635 1136 5647
rect 1555 5644 1567 5647
rect 1601 5644 1613 5678
rect 1555 5638 1613 5644
rect 2896 5635 2902 5687
rect 2954 5675 2960 5687
rect 4435 5678 4493 5684
rect 2954 5647 2999 5675
rect 2954 5635 2960 5647
rect 4435 5644 4447 5678
rect 4481 5675 4493 5678
rect 4912 5675 4918 5687
rect 4481 5647 4918 5675
rect 4481 5644 4493 5647
rect 4435 5638 4493 5644
rect 4912 5635 4918 5647
rect 4970 5635 4976 5687
rect 5200 5675 5206 5687
rect 5161 5647 5206 5675
rect 5200 5635 5206 5647
rect 5258 5635 5264 5687
rect 6832 5675 6838 5687
rect 6793 5647 6838 5675
rect 6832 5635 6838 5647
rect 6890 5635 6896 5687
rect 7216 5635 7222 5687
rect 7274 5675 7280 5687
rect 7603 5678 7661 5684
rect 7603 5675 7615 5678
rect 7274 5647 7615 5675
rect 7274 5635 7280 5647
rect 7603 5644 7615 5647
rect 7649 5644 7661 5678
rect 7603 5638 7661 5644
rect 8371 5678 8429 5684
rect 8371 5644 8383 5678
rect 8417 5644 8429 5678
rect 8371 5638 8429 5644
rect 5776 5561 5782 5613
rect 5834 5601 5840 5613
rect 5971 5604 6029 5610
rect 5971 5601 5983 5604
rect 5834 5573 5983 5601
rect 5834 5561 5840 5573
rect 5971 5570 5983 5573
rect 6017 5570 6029 5604
rect 5971 5564 6029 5570
rect 7600 5487 7606 5539
rect 7658 5527 7664 5539
rect 8386 5527 8414 5638
rect 8752 5635 8758 5687
rect 8810 5675 8816 5687
rect 9619 5678 9677 5684
rect 9619 5675 9631 5678
rect 8810 5647 9631 5675
rect 8810 5635 8816 5647
rect 9619 5644 9631 5647
rect 9665 5644 9677 5678
rect 9619 5638 9677 5644
rect 10192 5635 10198 5687
rect 10250 5675 10256 5687
rect 10387 5678 10445 5684
rect 10387 5675 10399 5678
rect 10250 5647 10399 5675
rect 10250 5635 10256 5647
rect 10387 5644 10399 5647
rect 10433 5644 10445 5678
rect 10387 5638 10445 5644
rect 10480 5635 10486 5687
rect 10538 5675 10544 5687
rect 11155 5678 11213 5684
rect 11155 5675 11167 5678
rect 10538 5647 11167 5675
rect 10538 5635 10544 5647
rect 11155 5644 11167 5647
rect 11201 5644 11213 5678
rect 12592 5675 12598 5687
rect 12553 5647 12598 5675
rect 11155 5638 11213 5644
rect 12592 5635 12598 5647
rect 12650 5635 12656 5687
rect 13360 5675 13366 5687
rect 13321 5647 13366 5675
rect 13360 5635 13366 5647
rect 13418 5635 13424 5687
rect 10576 5561 10582 5613
rect 10634 5601 10640 5613
rect 14338 5601 14366 5795
rect 20560 5783 20566 5795
rect 20618 5783 20624 5835
rect 33136 5823 33142 5835
rect 23170 5795 33142 5823
rect 22864 5709 22870 5761
rect 22922 5749 22928 5761
rect 23170 5749 23198 5795
rect 33136 5783 33142 5795
rect 33194 5783 33200 5835
rect 37744 5823 37750 5835
rect 33250 5795 37750 5823
rect 22922 5721 23198 5749
rect 22922 5709 22928 5721
rect 23536 5709 23542 5761
rect 23594 5749 23600 5761
rect 29872 5749 29878 5761
rect 23594 5721 29878 5749
rect 23594 5709 23600 5721
rect 29872 5709 29878 5721
rect 29930 5709 29936 5761
rect 32944 5709 32950 5761
rect 33002 5749 33008 5761
rect 33250 5749 33278 5795
rect 37744 5783 37750 5795
rect 37802 5783 37808 5835
rect 37858 5795 41054 5823
rect 33002 5721 33278 5749
rect 33002 5709 33008 5721
rect 35920 5709 35926 5761
rect 35978 5749 35984 5761
rect 37858 5749 37886 5795
rect 35978 5721 37886 5749
rect 41026 5749 41054 5795
rect 41968 5749 41974 5761
rect 41026 5721 41974 5749
rect 35978 5709 35984 5721
rect 41968 5709 41974 5721
rect 42026 5709 42032 5761
rect 14992 5675 14998 5687
rect 14953 5647 14998 5675
rect 14992 5635 14998 5647
rect 15050 5635 15056 5687
rect 15856 5675 15862 5687
rect 15817 5647 15862 5675
rect 15856 5635 15862 5647
rect 15914 5635 15920 5687
rect 16144 5635 16150 5687
rect 16202 5675 16208 5687
rect 16531 5678 16589 5684
rect 16531 5675 16543 5678
rect 16202 5647 16543 5675
rect 16202 5635 16208 5647
rect 16531 5644 16543 5647
rect 16577 5644 16589 5678
rect 17392 5675 17398 5687
rect 17353 5647 17398 5675
rect 16531 5638 16589 5644
rect 17392 5635 17398 5647
rect 17450 5635 17456 5687
rect 18736 5675 18742 5687
rect 18697 5647 18742 5675
rect 18736 5635 18742 5647
rect 18794 5635 18800 5687
rect 20176 5675 20182 5687
rect 20137 5647 20182 5675
rect 20176 5635 20182 5647
rect 20234 5635 20240 5687
rect 20560 5635 20566 5687
rect 20618 5675 20624 5687
rect 20947 5678 21005 5684
rect 20947 5675 20959 5678
rect 20618 5647 20959 5675
rect 20618 5635 20624 5647
rect 20947 5644 20959 5647
rect 20993 5644 21005 5678
rect 21712 5675 21718 5687
rect 21673 5647 21718 5675
rect 20947 5638 21005 5644
rect 21712 5635 21718 5647
rect 21770 5635 21776 5687
rect 22483 5678 22541 5684
rect 22483 5644 22495 5678
rect 22529 5644 22541 5678
rect 22483 5638 22541 5644
rect 10634 5573 14366 5601
rect 10634 5561 10640 5573
rect 21616 5561 21622 5613
rect 21674 5601 21680 5613
rect 22498 5601 22526 5638
rect 23056 5635 23062 5687
rect 23114 5675 23120 5687
rect 23251 5678 23309 5684
rect 23251 5675 23263 5678
rect 23114 5647 23263 5675
rect 23114 5635 23120 5647
rect 23251 5644 23263 5647
rect 23297 5644 23309 5678
rect 23251 5638 23309 5644
rect 23440 5635 23446 5687
rect 23498 5675 23504 5687
rect 24019 5678 24077 5684
rect 24019 5675 24031 5678
rect 23498 5647 24031 5675
rect 23498 5635 23504 5647
rect 24019 5644 24031 5647
rect 24065 5644 24077 5678
rect 24019 5638 24077 5644
rect 24592 5635 24598 5687
rect 24650 5675 24656 5687
rect 25459 5678 25517 5684
rect 25459 5675 25471 5678
rect 24650 5647 25471 5675
rect 24650 5635 24656 5647
rect 25459 5644 25471 5647
rect 25505 5644 25517 5678
rect 26224 5675 26230 5687
rect 26185 5647 26230 5675
rect 25459 5638 25517 5644
rect 26224 5635 26230 5647
rect 26282 5635 26288 5687
rect 26995 5678 27053 5684
rect 26995 5644 27007 5678
rect 27041 5644 27053 5678
rect 26995 5638 27053 5644
rect 21674 5573 22526 5601
rect 21674 5561 21680 5573
rect 26032 5561 26038 5613
rect 26090 5601 26096 5613
rect 27010 5601 27038 5638
rect 27376 5635 27382 5687
rect 27434 5675 27440 5687
rect 27763 5678 27821 5684
rect 27763 5675 27775 5678
rect 27434 5647 27775 5675
rect 27434 5635 27440 5647
rect 27763 5644 27775 5647
rect 27809 5644 27821 5678
rect 27763 5638 27821 5644
rect 27856 5635 27862 5687
rect 27914 5675 27920 5687
rect 28531 5678 28589 5684
rect 28531 5675 28543 5678
rect 27914 5647 28543 5675
rect 27914 5635 27920 5647
rect 28531 5644 28543 5647
rect 28577 5644 28589 5678
rect 28531 5638 28589 5644
rect 28816 5635 28822 5687
rect 28874 5675 28880 5687
rect 29299 5678 29357 5684
rect 29299 5675 29311 5678
rect 28874 5647 29311 5675
rect 28874 5635 28880 5647
rect 29299 5644 29311 5647
rect 29345 5644 29357 5678
rect 29299 5638 29357 5644
rect 30256 5635 30262 5687
rect 30314 5675 30320 5687
rect 30739 5678 30797 5684
rect 30739 5675 30751 5678
rect 30314 5647 30751 5675
rect 30314 5635 30320 5647
rect 30739 5644 30751 5647
rect 30785 5644 30797 5678
rect 30739 5638 30797 5644
rect 30832 5635 30838 5687
rect 30890 5675 30896 5687
rect 31507 5678 31565 5684
rect 31507 5675 31519 5678
rect 30890 5647 31519 5675
rect 30890 5635 30896 5647
rect 31507 5644 31519 5647
rect 31553 5644 31565 5678
rect 31507 5638 31565 5644
rect 31696 5635 31702 5687
rect 31754 5675 31760 5687
rect 32275 5678 32333 5684
rect 32275 5675 32287 5678
rect 31754 5647 32287 5675
rect 31754 5635 31760 5647
rect 32275 5644 32287 5647
rect 32321 5644 32333 5678
rect 32275 5638 32333 5644
rect 33136 5635 33142 5687
rect 33194 5675 33200 5687
rect 33811 5678 33869 5684
rect 33194 5647 33239 5675
rect 33194 5635 33200 5647
rect 33811 5644 33823 5678
rect 33857 5644 33869 5678
rect 34672 5675 34678 5687
rect 34633 5647 34678 5675
rect 33811 5638 33869 5644
rect 26090 5573 27038 5601
rect 26090 5561 26096 5573
rect 33232 5561 33238 5613
rect 33290 5601 33296 5613
rect 33826 5601 33854 5638
rect 34672 5635 34678 5647
rect 34730 5635 34736 5687
rect 36016 5675 36022 5687
rect 35977 5647 36022 5675
rect 36016 5635 36022 5647
rect 36074 5635 36080 5687
rect 36208 5635 36214 5687
rect 36266 5675 36272 5687
rect 36787 5678 36845 5684
rect 36787 5675 36799 5678
rect 36266 5647 36799 5675
rect 36266 5635 36272 5647
rect 36787 5644 36799 5647
rect 36833 5644 36845 5678
rect 37552 5675 37558 5687
rect 37513 5647 37558 5675
rect 36787 5638 36845 5644
rect 37552 5635 37558 5647
rect 37610 5635 37616 5687
rect 38323 5678 38381 5684
rect 38323 5644 38335 5678
rect 38369 5644 38381 5678
rect 39088 5675 39094 5687
rect 39049 5647 39094 5675
rect 38323 5638 38381 5644
rect 33290 5573 33854 5601
rect 33290 5561 33296 5573
rect 37456 5561 37462 5613
rect 37514 5601 37520 5613
rect 38338 5601 38366 5638
rect 39088 5635 39094 5647
rect 39146 5635 39152 5687
rect 39280 5635 39286 5687
rect 39338 5675 39344 5687
rect 39859 5678 39917 5684
rect 39859 5675 39871 5678
rect 39338 5647 39871 5675
rect 39338 5635 39344 5647
rect 39859 5644 39871 5647
rect 39905 5644 39917 5678
rect 39859 5638 39917 5644
rect 40720 5635 40726 5687
rect 40778 5675 40784 5687
rect 41299 5678 41357 5684
rect 41299 5675 41311 5678
rect 40778 5647 41311 5675
rect 40778 5635 40784 5647
rect 41299 5644 41311 5647
rect 41345 5644 41357 5678
rect 41299 5638 41357 5644
rect 41776 5635 41782 5687
rect 41834 5675 41840 5687
rect 42067 5678 42125 5684
rect 42067 5675 42079 5678
rect 41834 5647 42079 5675
rect 41834 5635 41840 5647
rect 42067 5644 42079 5647
rect 42113 5644 42125 5678
rect 42067 5638 42125 5644
rect 42256 5635 42262 5687
rect 42314 5675 42320 5687
rect 42835 5678 42893 5684
rect 42835 5675 42847 5678
rect 42314 5647 42847 5675
rect 42314 5635 42320 5647
rect 42835 5644 42847 5647
rect 42881 5644 42893 5678
rect 42835 5638 42893 5644
rect 43216 5635 43222 5687
rect 43274 5675 43280 5687
rect 43603 5678 43661 5684
rect 43603 5675 43615 5678
rect 43274 5647 43615 5675
rect 43274 5635 43280 5647
rect 43603 5644 43615 5647
rect 43649 5644 43661 5678
rect 43603 5638 43661 5644
rect 43696 5635 43702 5687
rect 43754 5675 43760 5687
rect 44371 5678 44429 5684
rect 44371 5675 44383 5678
rect 43754 5647 44383 5675
rect 43754 5635 43760 5647
rect 44371 5644 44383 5647
rect 44417 5644 44429 5678
rect 45136 5675 45142 5687
rect 45097 5647 45142 5675
rect 44371 5638 44429 5644
rect 45136 5635 45142 5647
rect 45194 5635 45200 5687
rect 46096 5635 46102 5687
rect 46154 5675 46160 5687
rect 46579 5678 46637 5684
rect 46579 5675 46591 5678
rect 46154 5647 46591 5675
rect 46154 5635 46160 5647
rect 46579 5644 46591 5647
rect 46625 5644 46637 5678
rect 46579 5638 46637 5644
rect 46672 5635 46678 5687
rect 46730 5675 46736 5687
rect 47347 5678 47405 5684
rect 47347 5675 47359 5678
rect 46730 5647 47359 5675
rect 46730 5635 46736 5647
rect 47347 5644 47359 5647
rect 47393 5644 47405 5678
rect 47347 5638 47405 5644
rect 47536 5635 47542 5687
rect 47594 5675 47600 5687
rect 48115 5678 48173 5684
rect 48115 5675 48127 5678
rect 47594 5647 48127 5675
rect 47594 5635 47600 5647
rect 48115 5644 48127 5647
rect 48161 5644 48173 5678
rect 48976 5675 48982 5687
rect 48937 5647 48982 5675
rect 48115 5638 48173 5644
rect 48976 5635 48982 5647
rect 49034 5635 49040 5687
rect 49648 5675 49654 5687
rect 49609 5647 49654 5675
rect 49648 5635 49654 5647
rect 49706 5635 49712 5687
rect 50515 5678 50573 5684
rect 50515 5644 50527 5678
rect 50561 5675 50573 5678
rect 50704 5675 50710 5687
rect 50561 5647 50710 5675
rect 50561 5644 50573 5647
rect 50515 5638 50573 5644
rect 50704 5635 50710 5647
rect 50762 5635 50768 5687
rect 52144 5675 52150 5687
rect 52105 5647 52150 5675
rect 52144 5635 52150 5647
rect 52202 5635 52208 5687
rect 52528 5635 52534 5687
rect 52586 5675 52592 5687
rect 52915 5678 52973 5684
rect 52915 5675 52927 5678
rect 52586 5647 52927 5675
rect 52586 5635 52592 5647
rect 52915 5644 52927 5647
rect 52961 5644 52973 5678
rect 53680 5675 53686 5687
rect 53641 5647 53686 5675
rect 52915 5638 52973 5644
rect 53680 5635 53686 5647
rect 53738 5635 53744 5687
rect 54451 5678 54509 5684
rect 54451 5644 54463 5678
rect 54497 5644 54509 5678
rect 54451 5638 54509 5644
rect 55987 5678 56045 5684
rect 55987 5644 55999 5678
rect 56033 5644 56045 5678
rect 57424 5675 57430 5687
rect 57385 5647 57430 5675
rect 55987 5638 56045 5644
rect 37514 5573 38366 5601
rect 37514 5561 37520 5573
rect 42736 5561 42742 5613
rect 42794 5601 42800 5613
rect 43312 5601 43318 5613
rect 42794 5573 43318 5601
rect 42794 5561 42800 5573
rect 43312 5561 43318 5573
rect 43370 5561 43376 5613
rect 53584 5561 53590 5613
rect 53642 5601 53648 5613
rect 54466 5601 54494 5638
rect 53642 5573 54494 5601
rect 56002 5601 56030 5638
rect 57424 5635 57430 5647
rect 57482 5635 57488 5687
rect 59632 5601 59638 5613
rect 56002 5573 59638 5601
rect 53642 5561 53648 5573
rect 59632 5561 59638 5573
rect 59690 5561 59696 5613
rect 7658 5499 8414 5527
rect 7658 5487 7664 5499
rect 20464 5487 20470 5539
rect 20522 5527 20528 5539
rect 29104 5527 29110 5539
rect 20522 5499 29110 5527
rect 20522 5487 20528 5499
rect 29104 5487 29110 5499
rect 29162 5487 29168 5539
rect 7120 5413 7126 5465
rect 7178 5453 7184 5465
rect 11536 5453 11542 5465
rect 7178 5425 11542 5453
rect 7178 5413 7184 5425
rect 11536 5413 11542 5425
rect 11594 5413 11600 5465
rect 12115 5456 12173 5462
rect 12115 5422 12127 5456
rect 12161 5453 12173 5456
rect 47632 5453 47638 5465
rect 12161 5425 47638 5453
rect 12161 5422 12173 5425
rect 12115 5416 12173 5422
rect 47632 5413 47638 5425
rect 47690 5413 47696 5465
rect 1152 5354 58848 5376
rect 1152 5302 4294 5354
rect 4346 5302 4358 5354
rect 4410 5302 4422 5354
rect 4474 5302 4486 5354
rect 4538 5302 35014 5354
rect 35066 5302 35078 5354
rect 35130 5302 35142 5354
rect 35194 5302 35206 5354
rect 35258 5302 58848 5354
rect 1152 5280 58848 5302
rect 4720 5191 4726 5243
rect 4778 5231 4784 5243
rect 7507 5234 7565 5240
rect 7507 5231 7519 5234
rect 4778 5203 7519 5231
rect 4778 5191 4784 5203
rect 7507 5200 7519 5203
rect 7553 5231 7565 5234
rect 7699 5234 7757 5240
rect 7699 5231 7711 5234
rect 7553 5203 7711 5231
rect 7553 5200 7565 5203
rect 7507 5194 7565 5200
rect 7699 5200 7711 5203
rect 7745 5200 7757 5234
rect 7699 5194 7757 5200
rect 7906 5203 8270 5231
rect 1840 5117 1846 5169
rect 1898 5117 1904 5169
rect 3568 5117 3574 5169
rect 3626 5157 3632 5169
rect 7906 5157 7934 5203
rect 3626 5129 7934 5157
rect 3626 5117 3632 5129
rect 1858 5083 1886 5117
rect 1858 5055 7968 5083
rect 8242 5069 8270 5203
rect 8371 5160 8429 5166
rect 8371 5126 8383 5160
rect 8417 5157 8429 5160
rect 8417 5129 8640 5157
rect 8417 5126 8429 5129
rect 8371 5120 8429 5126
rect 304 4969 310 5021
rect 362 5009 368 5021
rect 1555 5012 1613 5018
rect 1555 5009 1567 5012
rect 362 4981 1567 5009
rect 362 4969 368 4981
rect 1555 4978 1567 4981
rect 1601 4978 1613 5012
rect 1555 4972 1613 4978
rect 1840 4969 1846 5021
rect 1898 5009 1904 5021
rect 2323 5012 2381 5018
rect 2323 5009 2335 5012
rect 1898 4981 2335 5009
rect 1898 4969 1904 4981
rect 2323 4978 2335 4981
rect 2369 4978 2381 5012
rect 3088 5009 3094 5021
rect 3049 4981 3094 5009
rect 2323 4972 2381 4978
rect 3088 4969 3094 4981
rect 3146 4969 3152 5021
rect 4144 5009 4150 5021
rect 4105 4981 4150 5009
rect 4144 4969 4150 4981
rect 4202 4969 4208 5021
rect 5392 5009 5398 5021
rect 5353 4981 5398 5009
rect 5392 4969 5398 4981
rect 5450 4969 5456 5021
rect 6064 4969 6070 5021
rect 6122 5009 6128 5021
rect 6931 5012 6989 5018
rect 6931 5009 6943 5012
rect 6122 4981 6943 5009
rect 6122 4969 6128 4981
rect 6931 4978 6943 4981
rect 6977 4978 6989 5012
rect 9232 5009 9238 5021
rect 9193 4981 9238 5009
rect 6931 4972 6989 4978
rect 9232 4969 9238 4981
rect 9290 4969 9296 5021
rect 10099 5012 10157 5018
rect 10099 4978 10111 5012
rect 10145 5009 10157 5012
rect 10576 5009 10582 5021
rect 10145 4981 10582 5009
rect 10145 4978 10157 4981
rect 10099 4972 10157 4978
rect 10576 4969 10582 4981
rect 10634 4969 10640 5021
rect 10867 5012 10925 5018
rect 10867 4978 10879 5012
rect 10913 5009 10925 5012
rect 10960 5009 10966 5021
rect 10913 4981 10966 5009
rect 10913 4978 10925 4981
rect 10867 4972 10925 4978
rect 10960 4969 10966 4981
rect 11018 4969 11024 5021
rect 11824 4969 11830 5021
rect 11882 5009 11888 5021
rect 12211 5012 12269 5018
rect 12211 5009 12223 5012
rect 11882 4981 12223 5009
rect 11882 4969 11888 4981
rect 12211 4978 12223 4981
rect 12257 4978 12269 5012
rect 12211 4972 12269 4978
rect 12979 5012 13037 5018
rect 12979 4978 12991 5012
rect 13025 4978 13037 5012
rect 13936 5009 13942 5021
rect 13897 4981 13942 5009
rect 12979 4972 13037 4978
rect 12208 4821 12214 4873
rect 12266 4861 12272 4873
rect 12994 4861 13022 4972
rect 13936 4969 13942 4981
rect 13994 4969 14000 5021
rect 14416 4969 14422 5021
rect 14474 5009 14480 5021
rect 14707 5012 14765 5018
rect 14707 5009 14719 5012
rect 14474 4981 14719 5009
rect 14474 4969 14480 4981
rect 14707 4978 14719 4981
rect 14753 4978 14765 5012
rect 14707 4972 14765 4978
rect 14800 4969 14806 5021
rect 14858 5009 14864 5021
rect 15475 5012 15533 5018
rect 15475 5009 15487 5012
rect 14858 4981 15487 5009
rect 14858 4969 14864 4981
rect 15475 4978 15487 4981
rect 15521 4978 15533 5012
rect 15475 4972 15533 4978
rect 16339 5012 16397 5018
rect 16339 4978 16351 5012
rect 16385 5009 16397 5012
rect 16432 5009 16438 5021
rect 16385 4981 16438 5009
rect 16385 4978 16397 4981
rect 16339 4972 16397 4978
rect 16432 4969 16438 4981
rect 16490 4969 16496 5021
rect 17296 4969 17302 5021
rect 17354 5009 17360 5021
rect 17491 5012 17549 5018
rect 17491 5009 17503 5012
rect 17354 4981 17503 5009
rect 17354 4969 17360 4981
rect 17491 4978 17503 4981
rect 17537 4978 17549 5012
rect 17491 4972 17549 4978
rect 17968 4969 17974 5021
rect 18026 5009 18032 5021
rect 18259 5012 18317 5018
rect 18259 5009 18271 5012
rect 18026 4981 18271 5009
rect 18026 4969 18032 4981
rect 18259 4978 18271 4981
rect 18305 4978 18317 5012
rect 19024 5009 19030 5021
rect 18985 4981 19030 5009
rect 18259 4972 18317 4978
rect 19024 4969 19030 4981
rect 19082 4969 19088 5021
rect 19120 4969 19126 5021
rect 19178 5009 19184 5021
rect 19795 5012 19853 5018
rect 19795 5009 19807 5012
rect 19178 4981 19807 5009
rect 19178 4969 19184 4981
rect 19795 4978 19807 4981
rect 19841 4978 19853 5012
rect 19795 4972 19853 4978
rect 20464 4969 20470 5021
rect 20522 5009 20528 5021
rect 20563 5012 20621 5018
rect 20563 5009 20575 5012
rect 20522 4981 20575 5009
rect 20522 4969 20528 4981
rect 20563 4978 20575 4981
rect 20609 4978 20621 5012
rect 20563 4972 20621 4978
rect 20944 4969 20950 5021
rect 21002 5009 21008 5021
rect 21331 5012 21389 5018
rect 21331 5009 21343 5012
rect 21002 4981 21343 5009
rect 21002 4969 21008 4981
rect 21331 4978 21343 4981
rect 21377 4978 21389 5012
rect 21331 4972 21389 4978
rect 22096 4969 22102 5021
rect 22154 5009 22160 5021
rect 22771 5012 22829 5018
rect 22771 5009 22783 5012
rect 22154 4981 22783 5009
rect 22154 4969 22160 4981
rect 22771 4978 22783 4981
rect 22817 4978 22829 5012
rect 23536 5009 23542 5021
rect 23497 4981 23542 5009
rect 22771 4972 22829 4978
rect 23536 4969 23542 4981
rect 23594 4969 23600 5021
rect 24307 5012 24365 5018
rect 24307 4978 24319 5012
rect 24353 4978 24365 5012
rect 25072 5009 25078 5021
rect 25033 4981 25078 5009
rect 24307 4972 24365 4978
rect 23152 4895 23158 4947
rect 23210 4935 23216 4947
rect 24322 4935 24350 4972
rect 25072 4969 25078 4981
rect 25130 4969 25136 5021
rect 25840 5009 25846 5021
rect 25801 4981 25846 5009
rect 25840 4969 25846 4981
rect 25898 4969 25904 5021
rect 26608 5009 26614 5021
rect 26569 4981 26614 5009
rect 26608 4969 26614 4981
rect 26666 4969 26672 5021
rect 28048 5009 28054 5021
rect 28009 4981 28054 5009
rect 28048 4969 28054 4981
rect 28106 4969 28112 5021
rect 28912 5009 28918 5021
rect 28873 4981 28918 5009
rect 28912 4969 28918 4981
rect 28970 4969 28976 5021
rect 29008 4969 29014 5021
rect 29066 5009 29072 5021
rect 29587 5012 29645 5018
rect 29587 5009 29599 5012
rect 29066 4981 29599 5009
rect 29066 4969 29072 4981
rect 29587 4978 29599 4981
rect 29633 4978 29645 5012
rect 30352 5009 30358 5021
rect 30313 4981 30358 5009
rect 29587 4972 29645 4978
rect 30352 4969 30358 4981
rect 30410 4969 30416 5021
rect 30448 4969 30454 5021
rect 30506 5009 30512 5021
rect 31123 5012 31181 5018
rect 31123 5009 31135 5012
rect 30506 4981 31135 5009
rect 30506 4969 30512 4981
rect 31123 4978 31135 4981
rect 31169 4978 31181 5012
rect 31888 5009 31894 5021
rect 31849 4981 31894 5009
rect 31123 4972 31181 4978
rect 31888 4969 31894 4981
rect 31946 4969 31952 5021
rect 33328 5009 33334 5021
rect 33289 4981 33334 5009
rect 33328 4969 33334 4981
rect 33386 4969 33392 5021
rect 34096 5009 34102 5021
rect 34057 4981 34102 5009
rect 34096 4969 34102 4981
rect 34154 4969 34160 5021
rect 34768 4969 34774 5021
rect 34826 5009 34832 5021
rect 34867 5012 34925 5018
rect 34867 5009 34879 5012
rect 34826 4981 34879 5009
rect 34826 4969 34832 4981
rect 34867 4978 34879 4981
rect 34913 4978 34925 5012
rect 34867 4972 34925 4978
rect 35635 5012 35693 5018
rect 35635 4978 35647 5012
rect 35681 4978 35693 5012
rect 35635 4972 35693 4978
rect 36403 5012 36461 5018
rect 36403 4978 36415 5012
rect 36449 4978 36461 5012
rect 36403 4972 36461 4978
rect 23210 4907 24350 4935
rect 23210 4895 23216 4907
rect 34576 4895 34582 4947
rect 34634 4935 34640 4947
rect 35650 4935 35678 4972
rect 34634 4907 35678 4935
rect 36418 4935 36446 4972
rect 36496 4969 36502 5021
rect 36554 5009 36560 5021
rect 37171 5012 37229 5018
rect 37171 5009 37183 5012
rect 36554 4981 37183 5009
rect 36554 4969 36560 4981
rect 37171 4978 37183 4981
rect 37217 4978 37229 5012
rect 38608 5009 38614 5021
rect 38569 4981 38614 5009
rect 37171 4972 37229 4978
rect 38608 4969 38614 4981
rect 38666 4969 38672 5021
rect 39376 5009 39382 5021
rect 39337 4981 39382 5009
rect 39376 4969 39382 4981
rect 39434 4969 39440 5021
rect 40144 5009 40150 5021
rect 40105 4981 40150 5009
rect 40144 4969 40150 4981
rect 40202 4969 40208 5021
rect 40912 5009 40918 5021
rect 40873 4981 40918 5009
rect 40912 4969 40918 4981
rect 40970 4969 40976 5021
rect 41008 4969 41014 5021
rect 41066 5009 41072 5021
rect 41683 5012 41741 5018
rect 41683 5009 41695 5012
rect 41066 4981 41695 5009
rect 41066 4969 41072 4981
rect 41683 4978 41695 4981
rect 41729 4978 41741 5012
rect 41683 4972 41741 4978
rect 42064 4969 42070 5021
rect 42122 5009 42128 5021
rect 42451 5012 42509 5018
rect 42451 5009 42463 5012
rect 42122 4981 42463 5009
rect 42122 4969 42128 4981
rect 42451 4978 42463 4981
rect 42497 4978 42509 5012
rect 42451 4972 42509 4978
rect 43504 4969 43510 5021
rect 43562 5009 43568 5021
rect 43891 5012 43949 5018
rect 43891 5009 43903 5012
rect 43562 4981 43903 5009
rect 43562 4969 43568 4981
rect 43891 4978 43903 4981
rect 43937 4978 43949 5012
rect 44752 5009 44758 5021
rect 44713 4981 44758 5009
rect 43891 4972 43949 4978
rect 44752 4969 44758 4981
rect 44810 4969 44816 5021
rect 45424 5009 45430 5021
rect 45385 4981 45430 5009
rect 45424 4969 45430 4981
rect 45482 4969 45488 5021
rect 46192 5009 46198 5021
rect 46153 4981 46198 5009
rect 46192 4969 46198 4981
rect 46250 4969 46256 5021
rect 46384 4969 46390 5021
rect 46442 5009 46448 5021
rect 46963 5012 47021 5018
rect 46963 5009 46975 5012
rect 46442 4981 46975 5009
rect 46442 4969 46448 4981
rect 46963 4978 46975 4981
rect 47009 4978 47021 5012
rect 46963 4972 47021 4978
rect 47632 4969 47638 5021
rect 47690 5009 47696 5021
rect 47731 5012 47789 5018
rect 47731 5009 47743 5012
rect 47690 4981 47743 5009
rect 47690 4969 47696 4981
rect 47731 4978 47743 4981
rect 47777 4978 47789 5012
rect 49360 5009 49366 5021
rect 49321 4981 49366 5009
rect 47731 4972 47789 4978
rect 49360 4969 49366 4981
rect 49418 4969 49424 5021
rect 50416 5009 50422 5021
rect 50377 4981 50422 5009
rect 50416 4969 50422 4981
rect 50474 4969 50480 5021
rect 50896 4969 50902 5021
rect 50954 5009 50960 5021
rect 51091 5012 51149 5018
rect 51091 5009 51103 5012
rect 50954 4981 51103 5009
rect 50954 4969 50960 4981
rect 51091 4978 51103 4981
rect 51137 4978 51149 5012
rect 51856 5009 51862 5021
rect 51817 4981 51862 5009
rect 51091 4972 51149 4978
rect 51856 4969 51862 4981
rect 51914 4969 51920 5021
rect 51952 4969 51958 5021
rect 52010 5009 52016 5021
rect 52627 5012 52685 5018
rect 52627 5009 52639 5012
rect 52010 4981 52639 5009
rect 52010 4969 52016 4981
rect 52627 4978 52639 4981
rect 52673 4978 52685 5012
rect 52627 4972 52685 4978
rect 53296 4969 53302 5021
rect 53354 5009 53360 5021
rect 54451 5012 54509 5018
rect 54451 5009 54463 5012
rect 53354 4981 54463 5009
rect 53354 4969 53360 4981
rect 54451 4978 54463 4981
rect 54497 4978 54509 5012
rect 54451 4972 54509 4978
rect 55603 5012 55661 5018
rect 55603 4978 55615 5012
rect 55649 4978 55661 5012
rect 55603 4972 55661 4978
rect 56371 5012 56429 5018
rect 56371 4978 56383 5012
rect 56417 4978 56429 5012
rect 57040 5009 57046 5021
rect 57001 4981 57046 5009
rect 56371 4972 56429 4978
rect 36880 4935 36886 4947
rect 36418 4907 36886 4935
rect 34634 4895 34640 4907
rect 36880 4895 36886 4907
rect 36938 4895 36944 4947
rect 12266 4833 13022 4861
rect 55618 4861 55646 4972
rect 56386 4935 56414 4972
rect 57040 4969 57046 4981
rect 57098 4969 57104 5021
rect 57808 4935 57814 4947
rect 56386 4907 57814 4935
rect 57808 4895 57814 4907
rect 57866 4895 57872 4947
rect 59248 4861 59254 4873
rect 55618 4833 59254 4861
rect 12266 4821 12272 4833
rect 59248 4821 59254 4833
rect 59306 4821 59312 4873
rect 8848 4747 8854 4799
rect 8906 4787 8912 4799
rect 9904 4787 9910 4799
rect 8906 4759 9910 4787
rect 8906 4747 8912 4759
rect 9904 4747 9910 4759
rect 9962 4747 9968 4799
rect 39952 4747 39958 4799
rect 40010 4787 40016 4799
rect 57715 4790 57773 4796
rect 57715 4787 57727 4790
rect 40010 4759 57727 4787
rect 40010 4747 40016 4759
rect 57715 4756 57727 4759
rect 57761 4787 57773 4790
rect 57811 4790 57869 4796
rect 57811 4787 57823 4790
rect 57761 4759 57823 4787
rect 57761 4756 57773 4759
rect 57715 4750 57773 4756
rect 57811 4756 57823 4759
rect 57857 4756 57869 4790
rect 57811 4750 57869 4756
rect 1152 4688 58848 4710
rect 1152 4636 19654 4688
rect 19706 4636 19718 4688
rect 19770 4636 19782 4688
rect 19834 4636 19846 4688
rect 19898 4636 50374 4688
rect 50426 4636 50438 4688
rect 50490 4636 50502 4688
rect 50554 4636 50566 4688
rect 50618 4636 58848 4688
rect 1152 4614 58848 4636
rect 7408 4525 7414 4577
rect 7466 4565 7472 4577
rect 15763 4568 15821 4574
rect 15763 4565 15775 4568
rect 7466 4537 15775 4565
rect 7466 4525 7472 4537
rect 15763 4534 15775 4537
rect 15809 4534 15821 4568
rect 15763 4528 15821 4534
rect 43792 4525 43798 4577
rect 43850 4565 43856 4577
rect 44083 4568 44141 4574
rect 44083 4565 44095 4568
rect 43850 4537 44095 4565
rect 43850 4525 43856 4537
rect 44083 4534 44095 4537
rect 44129 4565 44141 4568
rect 44129 4537 44318 4565
rect 44129 4534 44141 4537
rect 44083 4528 44141 4534
rect 8080 4451 8086 4503
rect 8138 4491 8144 4503
rect 8944 4491 8950 4503
rect 8138 4463 8950 4491
rect 8138 4451 8144 4463
rect 8944 4451 8950 4463
rect 9002 4451 9008 4503
rect 10768 4451 10774 4503
rect 10826 4491 10832 4503
rect 11440 4491 11446 4503
rect 10826 4463 11446 4491
rect 10826 4451 10832 4463
rect 11440 4451 11446 4463
rect 11498 4451 11504 4503
rect 11536 4451 11542 4503
rect 11594 4491 11600 4503
rect 16531 4494 16589 4500
rect 16531 4491 16543 4494
rect 11594 4463 16543 4491
rect 11594 4451 11600 4463
rect 16531 4460 16543 4463
rect 16577 4460 16589 4494
rect 16531 4454 16589 4460
rect 17299 4494 17357 4500
rect 17299 4460 17311 4494
rect 17345 4460 17357 4494
rect 17299 4454 17357 4460
rect 784 4377 790 4429
rect 842 4417 848 4429
rect 842 4389 2366 4417
rect 842 4377 848 4389
rect 1168 4303 1174 4355
rect 1226 4343 1232 4355
rect 2338 4352 2366 4389
rect 8272 4377 8278 4429
rect 8330 4417 8336 4429
rect 17314 4417 17342 4454
rect 32944 4451 32950 4503
rect 33002 4491 33008 4503
rect 33904 4491 33910 4503
rect 33002 4463 33910 4491
rect 33002 4451 33008 4463
rect 33904 4451 33910 4463
rect 33962 4451 33968 4503
rect 8330 4389 17342 4417
rect 8330 4377 8336 4389
rect 17584 4377 17590 4429
rect 17642 4417 17648 4429
rect 17642 4389 18590 4417
rect 17642 4377 17648 4389
rect 1555 4346 1613 4352
rect 1555 4343 1567 4346
rect 1226 4315 1567 4343
rect 1226 4303 1232 4315
rect 1555 4312 1567 4315
rect 1601 4312 1613 4346
rect 1555 4306 1613 4312
rect 2323 4346 2381 4352
rect 2323 4312 2335 4346
rect 2369 4312 2381 4346
rect 3091 4346 3149 4352
rect 3091 4343 3103 4346
rect 2323 4306 2381 4312
rect 2866 4315 3103 4343
rect 1360 4229 1366 4281
rect 1418 4269 1424 4281
rect 2866 4269 2894 4315
rect 3091 4312 3103 4315
rect 3137 4312 3149 4346
rect 3091 4306 3149 4312
rect 4339 4346 4397 4352
rect 4339 4312 4351 4346
rect 4385 4312 4397 4346
rect 4339 4306 4397 4312
rect 1418 4241 2894 4269
rect 1418 4229 1424 4241
rect 3760 4229 3766 4281
rect 3818 4269 3824 4281
rect 4354 4269 4382 4306
rect 4720 4303 4726 4355
rect 4778 4343 4784 4355
rect 5107 4346 5165 4352
rect 5107 4343 5119 4346
rect 4778 4315 5119 4343
rect 4778 4303 4784 4315
rect 5107 4312 5119 4315
rect 5153 4312 5165 4346
rect 5875 4346 5933 4352
rect 5875 4343 5887 4346
rect 5107 4306 5165 4312
rect 5602 4315 5887 4343
rect 3818 4241 4382 4269
rect 3818 4229 3824 4241
rect 3472 4155 3478 4207
rect 3530 4195 3536 4207
rect 4912 4195 4918 4207
rect 3530 4167 4918 4195
rect 3530 4155 3536 4167
rect 4912 4155 4918 4167
rect 4970 4155 4976 4207
rect 5104 4155 5110 4207
rect 5162 4195 5168 4207
rect 5602 4195 5630 4315
rect 5875 4312 5887 4315
rect 5921 4312 5933 4346
rect 5875 4306 5933 4312
rect 6643 4346 6701 4352
rect 6643 4312 6655 4346
rect 6689 4312 6701 4346
rect 7408 4343 7414 4355
rect 7369 4315 7414 4343
rect 6643 4306 6701 4312
rect 5680 4229 5686 4281
rect 5738 4269 5744 4281
rect 6658 4269 6686 4306
rect 7408 4303 7414 4315
rect 7466 4303 7472 4355
rect 8179 4346 8237 4352
rect 8179 4343 8191 4346
rect 7522 4315 8191 4343
rect 5738 4241 6686 4269
rect 5738 4229 5744 4241
rect 5162 4167 5630 4195
rect 5162 4155 5168 4167
rect 6448 4155 6454 4207
rect 6506 4195 6512 4207
rect 7522 4195 7550 4315
rect 8179 4312 8191 4315
rect 8225 4312 8237 4346
rect 9616 4343 9622 4355
rect 9577 4315 9622 4343
rect 8179 4306 8237 4312
rect 9616 4303 9622 4315
rect 9674 4303 9680 4355
rect 10384 4343 10390 4355
rect 10345 4315 10390 4343
rect 10384 4303 10390 4315
rect 10442 4303 10448 4355
rect 10768 4303 10774 4355
rect 10826 4343 10832 4355
rect 11155 4346 11213 4352
rect 11155 4343 11167 4346
rect 10826 4315 11167 4343
rect 10826 4303 10832 4315
rect 11155 4312 11167 4315
rect 11201 4312 11213 4346
rect 11923 4346 11981 4352
rect 11923 4343 11935 4346
rect 11155 4306 11213 4312
rect 11266 4315 11935 4343
rect 7888 4229 7894 4281
rect 7946 4269 7952 4281
rect 9808 4269 9814 4281
rect 7946 4241 9814 4269
rect 7946 4229 7952 4241
rect 9808 4229 9814 4241
rect 9866 4229 9872 4281
rect 6506 4167 7550 4195
rect 6506 4155 6512 4167
rect 9328 4155 9334 4207
rect 9386 4195 9392 4207
rect 9386 4167 11102 4195
rect 9386 4155 9392 4167
rect 976 4081 982 4133
rect 1034 4121 1040 4133
rect 2320 4121 2326 4133
rect 1034 4093 2326 4121
rect 1034 4081 1040 4093
rect 2320 4081 2326 4093
rect 2378 4081 2384 4133
rect 2416 4081 2422 4133
rect 2474 4121 2480 4133
rect 5008 4121 5014 4133
rect 2474 4093 5014 4121
rect 2474 4081 2480 4093
rect 5008 4081 5014 4093
rect 5066 4081 5072 4133
rect 9040 4081 9046 4133
rect 9098 4121 9104 4133
rect 10960 4121 10966 4133
rect 9098 4093 10966 4121
rect 9098 4081 9104 4093
rect 10960 4081 10966 4093
rect 11018 4081 11024 4133
rect 11074 4121 11102 4167
rect 11152 4155 11158 4207
rect 11210 4195 11216 4207
rect 11266 4195 11294 4315
rect 11923 4312 11935 4315
rect 11969 4312 11981 4346
rect 11923 4306 11981 4312
rect 12691 4346 12749 4352
rect 12691 4312 12703 4346
rect 12737 4312 12749 4346
rect 13552 4343 13558 4355
rect 13513 4315 13558 4343
rect 12691 4306 12749 4312
rect 11440 4229 11446 4281
rect 11498 4269 11504 4281
rect 12706 4269 12734 4306
rect 13552 4303 13558 4315
rect 13610 4303 13616 4355
rect 15472 4343 15478 4355
rect 15433 4315 15478 4343
rect 15472 4303 15478 4315
rect 15530 4303 15536 4355
rect 15952 4303 15958 4355
rect 16010 4343 16016 4355
rect 18562 4352 18590 4389
rect 24400 4377 24406 4429
rect 24458 4417 24464 4429
rect 44290 4426 44318 4537
rect 56752 4451 56758 4503
rect 56810 4491 56816 4503
rect 57328 4491 57334 4503
rect 56810 4463 57334 4491
rect 56810 4451 56816 4463
rect 57328 4451 57334 4463
rect 57386 4451 57392 4503
rect 44275 4420 44333 4426
rect 24458 4389 25598 4417
rect 24458 4377 24464 4389
rect 16243 4346 16301 4352
rect 16243 4343 16255 4346
rect 16010 4315 16255 4343
rect 16010 4303 16016 4315
rect 16243 4312 16255 4315
rect 16289 4312 16301 4346
rect 16243 4306 16301 4312
rect 17011 4346 17069 4352
rect 17011 4312 17023 4346
rect 17057 4312 17069 4346
rect 17011 4306 17069 4312
rect 17779 4346 17837 4352
rect 17779 4312 17791 4346
rect 17825 4312 17837 4346
rect 17779 4306 17837 4312
rect 18547 4346 18605 4352
rect 18547 4312 18559 4346
rect 18593 4312 18605 4346
rect 20272 4343 20278 4355
rect 20233 4315 20278 4343
rect 18547 4306 18605 4312
rect 11498 4241 12734 4269
rect 11498 4229 11504 4241
rect 13840 4229 13846 4281
rect 13898 4269 13904 4281
rect 14512 4269 14518 4281
rect 13898 4241 14518 4269
rect 13898 4229 13904 4241
rect 14512 4229 14518 4241
rect 14570 4229 14576 4281
rect 11210 4167 11294 4195
rect 11362 4167 14078 4195
rect 11210 4155 11216 4167
rect 11362 4121 11390 4167
rect 11074 4093 11390 4121
rect 11920 4081 11926 4133
rect 11978 4121 11984 4133
rect 13072 4121 13078 4133
rect 11978 4093 13078 4121
rect 11978 4081 11984 4093
rect 13072 4081 13078 4093
rect 13130 4081 13136 4133
rect 14050 4121 14078 4167
rect 14128 4155 14134 4207
rect 14186 4195 14192 4207
rect 14704 4195 14710 4207
rect 14186 4167 14710 4195
rect 14186 4155 14192 4167
rect 14704 4155 14710 4167
rect 14762 4155 14768 4207
rect 16240 4155 16246 4207
rect 16298 4195 16304 4207
rect 17026 4195 17054 4306
rect 16298 4167 17054 4195
rect 16298 4155 16304 4167
rect 16816 4121 16822 4133
rect 14050 4093 16822 4121
rect 16816 4081 16822 4093
rect 16874 4081 16880 4133
rect 16912 4081 16918 4133
rect 16970 4121 16976 4133
rect 17794 4121 17822 4306
rect 20272 4303 20278 4315
rect 20330 4303 20336 4355
rect 21040 4343 21046 4355
rect 21001 4315 21046 4343
rect 21040 4303 21046 4315
rect 21098 4303 21104 4355
rect 21808 4343 21814 4355
rect 21769 4315 21814 4343
rect 21808 4303 21814 4315
rect 21866 4303 21872 4355
rect 23248 4343 23254 4355
rect 23209 4315 23254 4343
rect 23248 4303 23254 4315
rect 23306 4303 23312 4355
rect 24016 4343 24022 4355
rect 23977 4315 24022 4343
rect 24016 4303 24022 4315
rect 24074 4303 24080 4355
rect 25456 4343 25462 4355
rect 25417 4315 25462 4343
rect 25456 4303 25462 4315
rect 25514 4303 25520 4355
rect 25570 4343 25598 4389
rect 31330 4389 31838 4417
rect 25570 4315 25982 4343
rect 21232 4229 21238 4281
rect 21290 4269 21296 4281
rect 22000 4269 22006 4281
rect 21290 4241 22006 4269
rect 21290 4229 21296 4241
rect 22000 4229 22006 4241
rect 22058 4229 22064 4281
rect 22768 4269 22774 4281
rect 22729 4241 22774 4269
rect 22768 4229 22774 4241
rect 22826 4229 22832 4281
rect 24208 4229 24214 4281
rect 24266 4269 24272 4281
rect 25840 4269 25846 4281
rect 24266 4241 25846 4269
rect 24266 4229 24272 4241
rect 25840 4229 25846 4241
rect 25898 4229 25904 4281
rect 25954 4269 25982 4315
rect 26128 4303 26134 4355
rect 26186 4343 26192 4355
rect 26227 4346 26285 4352
rect 26227 4343 26239 4346
rect 26186 4315 26239 4343
rect 26186 4303 26192 4315
rect 26227 4312 26239 4315
rect 26273 4312 26285 4346
rect 26227 4306 26285 4312
rect 26512 4303 26518 4355
rect 26570 4343 26576 4355
rect 26995 4346 27053 4352
rect 26995 4343 27007 4346
rect 26570 4315 27007 4343
rect 26570 4303 26576 4315
rect 26995 4312 27007 4315
rect 27041 4312 27053 4346
rect 28336 4343 28342 4355
rect 28297 4315 28342 4343
rect 26995 4306 27053 4312
rect 28336 4303 28342 4315
rect 28394 4303 28400 4355
rect 29104 4343 29110 4355
rect 29065 4315 29110 4343
rect 29104 4303 29110 4315
rect 29162 4303 29168 4355
rect 30928 4343 30934 4355
rect 30889 4315 30934 4343
rect 30928 4303 30934 4315
rect 30986 4303 30992 4355
rect 25954 4241 28478 4269
rect 22288 4155 22294 4207
rect 22346 4195 22352 4207
rect 22960 4195 22966 4207
rect 22346 4167 22966 4195
rect 22346 4155 22352 4167
rect 22960 4155 22966 4167
rect 23018 4155 23024 4207
rect 25360 4155 25366 4207
rect 25418 4195 25424 4207
rect 26224 4195 26230 4207
rect 25418 4167 26230 4195
rect 25418 4155 25424 4167
rect 26224 4155 26230 4167
rect 26282 4155 26288 4207
rect 28450 4195 28478 4241
rect 31330 4195 31358 4389
rect 31696 4343 31702 4355
rect 31657 4315 31702 4343
rect 31696 4303 31702 4315
rect 31754 4303 31760 4355
rect 31810 4343 31838 4389
rect 44275 4386 44287 4420
rect 44321 4386 44333 4420
rect 44275 4380 44333 4386
rect 32752 4343 32758 4355
rect 31810 4315 31934 4343
rect 32713 4315 32758 4343
rect 31906 4269 31934 4315
rect 32752 4303 32758 4315
rect 32810 4303 32816 4355
rect 33904 4343 33910 4355
rect 33865 4315 33910 4343
rect 33904 4303 33910 4315
rect 33962 4303 33968 4355
rect 34576 4303 34582 4355
rect 34634 4343 34640 4355
rect 34675 4346 34733 4352
rect 34675 4343 34687 4346
rect 34634 4315 34687 4343
rect 34634 4303 34640 4315
rect 34675 4312 34687 4315
rect 34721 4312 34733 4346
rect 36019 4346 36077 4352
rect 36019 4343 36031 4346
rect 34675 4306 34733 4312
rect 34786 4315 36031 4343
rect 31906 4241 33134 4269
rect 28450 4167 31358 4195
rect 31408 4155 31414 4207
rect 31466 4195 31472 4207
rect 32368 4195 32374 4207
rect 31466 4167 32374 4195
rect 31466 4155 31472 4167
rect 32368 4155 32374 4167
rect 32426 4155 32432 4207
rect 33106 4195 33134 4241
rect 34192 4229 34198 4281
rect 34250 4269 34256 4281
rect 34786 4269 34814 4315
rect 36019 4312 36031 4315
rect 36065 4312 36077 4346
rect 36784 4343 36790 4355
rect 36745 4315 36790 4343
rect 36019 4306 36077 4312
rect 36784 4303 36790 4315
rect 36842 4303 36848 4355
rect 37555 4346 37613 4352
rect 37555 4312 37567 4346
rect 37601 4312 37613 4346
rect 38992 4343 38998 4355
rect 38953 4315 38998 4343
rect 37555 4306 37613 4312
rect 34250 4241 34814 4269
rect 34250 4229 34256 4241
rect 37168 4229 37174 4281
rect 37226 4269 37232 4281
rect 37570 4269 37598 4306
rect 38992 4303 38998 4315
rect 39050 4303 39056 4355
rect 39760 4343 39766 4355
rect 39721 4315 39766 4343
rect 39760 4303 39766 4315
rect 39818 4303 39824 4355
rect 41968 4343 41974 4355
rect 41929 4315 41974 4343
rect 41968 4303 41974 4315
rect 42026 4303 42032 4355
rect 42352 4303 42358 4355
rect 42410 4343 42416 4355
rect 42739 4346 42797 4352
rect 42739 4343 42751 4346
rect 42410 4315 42751 4343
rect 42410 4303 42416 4315
rect 42739 4312 42751 4315
rect 42785 4312 42797 4346
rect 42739 4306 42797 4312
rect 43408 4303 43414 4355
rect 43466 4343 43472 4355
rect 43507 4346 43565 4352
rect 43507 4343 43519 4346
rect 43466 4315 43519 4343
rect 43466 4303 43472 4315
rect 43507 4312 43519 4315
rect 43553 4312 43565 4346
rect 44944 4343 44950 4355
rect 44905 4315 44950 4343
rect 43507 4306 43565 4312
rect 44944 4303 44950 4315
rect 45002 4303 45008 4355
rect 46768 4343 46774 4355
rect 46729 4315 46774 4343
rect 46768 4303 46774 4315
rect 46826 4303 46832 4355
rect 47539 4346 47597 4352
rect 47539 4312 47551 4346
rect 47585 4312 47597 4346
rect 47539 4306 47597 4312
rect 37226 4241 37598 4269
rect 37226 4229 37232 4241
rect 38128 4229 38134 4281
rect 38186 4269 38192 4281
rect 39088 4269 39094 4281
rect 38186 4241 39094 4269
rect 38186 4229 38192 4241
rect 39088 4229 39094 4241
rect 39146 4229 39152 4281
rect 41488 4229 41494 4281
rect 41546 4269 41552 4281
rect 41776 4269 41782 4281
rect 41546 4241 41782 4269
rect 41546 4229 41552 4241
rect 41776 4229 41782 4241
rect 41834 4229 41840 4281
rect 43600 4229 43606 4281
rect 43658 4269 43664 4281
rect 44368 4269 44374 4281
rect 43658 4241 44374 4269
rect 43658 4229 43664 4241
rect 44368 4229 44374 4241
rect 44426 4229 44432 4281
rect 44464 4229 44470 4281
rect 44522 4269 44528 4281
rect 45136 4269 45142 4281
rect 44522 4241 45142 4269
rect 44522 4229 44528 4241
rect 45136 4229 45142 4241
rect 45194 4229 45200 4281
rect 47440 4229 47446 4281
rect 47498 4269 47504 4281
rect 47554 4269 47582 4306
rect 47824 4303 47830 4355
rect 47882 4343 47888 4355
rect 48307 4346 48365 4352
rect 48307 4343 48319 4346
rect 47882 4315 48319 4343
rect 47882 4303 47888 4315
rect 48307 4312 48319 4315
rect 48353 4312 48365 4346
rect 48307 4306 48365 4312
rect 49075 4346 49133 4352
rect 49075 4312 49087 4346
rect 49121 4312 49133 4346
rect 49075 4306 49133 4312
rect 47498 4241 47582 4269
rect 47498 4229 47504 4241
rect 48592 4229 48598 4281
rect 48650 4269 48656 4281
rect 49090 4269 49118 4306
rect 49168 4303 49174 4355
rect 49226 4343 49232 4355
rect 49843 4346 49901 4352
rect 49843 4343 49855 4346
rect 49226 4315 49855 4343
rect 49226 4303 49232 4315
rect 49843 4312 49855 4315
rect 49889 4312 49901 4346
rect 49843 4306 49901 4312
rect 50611 4346 50669 4352
rect 50611 4312 50623 4346
rect 50657 4312 50669 4346
rect 50611 4306 50669 4312
rect 51859 4346 51917 4352
rect 51859 4312 51871 4346
rect 51905 4312 51917 4346
rect 52624 4343 52630 4355
rect 52585 4315 52630 4343
rect 51859 4306 51917 4312
rect 48650 4241 49118 4269
rect 48650 4229 48656 4241
rect 49936 4229 49942 4281
rect 49994 4269 50000 4281
rect 50626 4269 50654 4306
rect 49994 4241 50654 4269
rect 49994 4229 50000 4241
rect 50992 4229 50998 4281
rect 51050 4269 51056 4281
rect 51874 4269 51902 4306
rect 52624 4303 52630 4315
rect 52682 4303 52688 4355
rect 53395 4346 53453 4352
rect 53395 4312 53407 4346
rect 53441 4312 53453 4346
rect 53395 4306 53453 4312
rect 51050 4241 51902 4269
rect 51050 4229 51056 4241
rect 53008 4229 53014 4281
rect 53066 4269 53072 4281
rect 53410 4269 53438 4306
rect 54064 4303 54070 4355
rect 54122 4343 54128 4355
rect 54163 4346 54221 4352
rect 54163 4343 54175 4346
rect 54122 4315 54175 4343
rect 54122 4303 54128 4315
rect 54163 4312 54175 4315
rect 54209 4312 54221 4346
rect 55600 4343 55606 4355
rect 55561 4315 55606 4343
rect 54163 4306 54221 4312
rect 55600 4303 55606 4315
rect 55658 4303 55664 4355
rect 57235 4346 57293 4352
rect 57235 4312 57247 4346
rect 57281 4343 57293 4346
rect 57328 4343 57334 4355
rect 57281 4315 57334 4343
rect 57281 4312 57293 4315
rect 57235 4306 57293 4312
rect 57328 4303 57334 4315
rect 57386 4303 57392 4355
rect 53066 4241 53438 4269
rect 53066 4229 53072 4241
rect 56560 4229 56566 4281
rect 56618 4269 56624 4281
rect 58288 4269 58294 4281
rect 56618 4241 58294 4269
rect 56618 4229 56624 4241
rect 58288 4229 58294 4241
rect 58346 4229 58352 4281
rect 55123 4198 55181 4204
rect 55123 4195 55135 4198
rect 33106 4167 55135 4195
rect 55123 4164 55135 4167
rect 55169 4164 55181 4198
rect 55123 4158 55181 4164
rect 55984 4155 55990 4207
rect 56042 4195 56048 4207
rect 57904 4195 57910 4207
rect 56042 4167 57910 4195
rect 56042 4155 56048 4167
rect 57904 4155 57910 4167
rect 57962 4155 57968 4207
rect 16970 4093 17822 4121
rect 16970 4081 16976 4093
rect 25552 4081 25558 4133
rect 25610 4121 25616 4133
rect 25936 4121 25942 4133
rect 25610 4093 25942 4121
rect 25610 4081 25616 4093
rect 25936 4081 25942 4093
rect 25994 4081 26000 4133
rect 26416 4081 26422 4133
rect 26474 4121 26480 4133
rect 28048 4121 28054 4133
rect 26474 4093 28054 4121
rect 26474 4081 26480 4093
rect 28048 4081 28054 4093
rect 28106 4081 28112 4133
rect 28240 4081 28246 4133
rect 28298 4121 28304 4133
rect 29008 4121 29014 4133
rect 28298 4093 29014 4121
rect 28298 4081 28304 4093
rect 29008 4081 29014 4093
rect 29066 4081 29072 4133
rect 29296 4081 29302 4133
rect 29354 4121 29360 4133
rect 30448 4121 30454 4133
rect 29354 4093 30454 4121
rect 29354 4081 29360 4093
rect 30448 4081 30454 4093
rect 30506 4081 30512 4133
rect 31792 4081 31798 4133
rect 31850 4121 31856 4133
rect 33040 4121 33046 4133
rect 31850 4093 33046 4121
rect 31850 4081 31856 4093
rect 33040 4081 33046 4093
rect 33098 4081 33104 4133
rect 33808 4081 33814 4133
rect 33866 4121 33872 4133
rect 34672 4121 34678 4133
rect 33866 4093 34678 4121
rect 33866 4081 33872 4093
rect 34672 4081 34678 4093
rect 34730 4081 34736 4133
rect 38512 4081 38518 4133
rect 38570 4121 38576 4133
rect 40144 4121 40150 4133
rect 38570 4093 40150 4121
rect 38570 4081 38576 4093
rect 40144 4081 40150 4093
rect 40202 4081 40208 4133
rect 48112 4081 48118 4133
rect 48170 4121 48176 4133
rect 48976 4121 48982 4133
rect 48170 4093 48982 4121
rect 48170 4081 48176 4093
rect 48976 4081 48982 4093
rect 49034 4081 49040 4133
rect 49264 4081 49270 4133
rect 49322 4121 49328 4133
rect 50704 4121 50710 4133
rect 49322 4093 50710 4121
rect 49322 4081 49328 4093
rect 50704 4081 50710 4093
rect 50762 4081 50768 4133
rect 1152 4022 58848 4044
rect 1152 3970 4294 4022
rect 4346 3970 4358 4022
rect 4410 3970 4422 4022
rect 4474 3970 4486 4022
rect 4538 3970 35014 4022
rect 35066 3970 35078 4022
rect 35130 3970 35142 4022
rect 35194 3970 35206 4022
rect 35258 3970 58848 4022
rect 1152 3948 58848 3970
rect 1936 3859 1942 3911
rect 1994 3899 2000 3911
rect 2992 3899 2998 3911
rect 1994 3871 2998 3899
rect 1994 3859 2000 3871
rect 2992 3859 2998 3871
rect 3050 3859 3056 3911
rect 7888 3859 7894 3911
rect 7946 3899 7952 3911
rect 9232 3899 9238 3911
rect 7946 3871 9238 3899
rect 7946 3859 7952 3871
rect 9232 3859 9238 3871
rect 9290 3859 9296 3911
rect 9808 3859 9814 3911
rect 9866 3899 9872 3911
rect 9866 3871 10718 3899
rect 9866 3859 9872 3871
rect 496 3785 502 3837
rect 554 3825 560 3837
rect 1648 3825 1654 3837
rect 554 3797 1654 3825
rect 554 3785 560 3797
rect 1648 3785 1654 3797
rect 1706 3785 1712 3837
rect 2320 3785 2326 3837
rect 2378 3825 2384 3837
rect 3088 3825 3094 3837
rect 2378 3797 3094 3825
rect 2378 3785 2384 3797
rect 3088 3785 3094 3797
rect 3146 3785 3152 3837
rect 8272 3785 8278 3837
rect 8330 3825 8336 3837
rect 10576 3825 10582 3837
rect 8330 3797 10582 3825
rect 8330 3785 8336 3797
rect 10576 3785 10582 3797
rect 10634 3785 10640 3837
rect 10690 3834 10718 3871
rect 11536 3859 11542 3911
rect 11594 3899 11600 3911
rect 11594 3871 16478 3899
rect 11594 3859 11600 3871
rect 10675 3828 10733 3834
rect 10675 3794 10687 3828
rect 10721 3794 10733 3828
rect 16450 3825 16478 3871
rect 16528 3859 16534 3911
rect 16586 3899 16592 3911
rect 17392 3899 17398 3911
rect 16586 3871 17398 3899
rect 16586 3859 16592 3871
rect 17392 3859 17398 3871
rect 17450 3859 17456 3911
rect 18352 3859 18358 3911
rect 18410 3899 18416 3911
rect 19024 3899 19030 3911
rect 18410 3871 19030 3899
rect 18410 3859 18416 3871
rect 19024 3859 19030 3871
rect 19082 3859 19088 3911
rect 19216 3859 19222 3911
rect 19274 3899 19280 3911
rect 19315 3902 19373 3908
rect 19315 3899 19327 3902
rect 19274 3871 19327 3899
rect 19274 3859 19280 3871
rect 19315 3868 19327 3871
rect 19361 3868 19373 3902
rect 19315 3862 19373 3868
rect 19408 3859 19414 3911
rect 19466 3899 19472 3911
rect 20464 3899 20470 3911
rect 19466 3871 20470 3899
rect 19466 3859 19472 3871
rect 20464 3859 20470 3871
rect 20522 3859 20528 3911
rect 21328 3859 21334 3911
rect 21386 3899 21392 3911
rect 22096 3899 22102 3911
rect 21386 3871 22102 3899
rect 21386 3859 21392 3871
rect 22096 3859 22102 3871
rect 22154 3859 22160 3911
rect 23824 3859 23830 3911
rect 23882 3899 23888 3911
rect 25072 3899 25078 3911
rect 23882 3871 25078 3899
rect 23882 3859 23888 3871
rect 25072 3859 25078 3871
rect 25130 3859 25136 3911
rect 25936 3859 25942 3911
rect 25994 3899 26000 3911
rect 26896 3899 26902 3911
rect 25994 3871 26902 3899
rect 25994 3859 26000 3871
rect 26896 3859 26902 3871
rect 26954 3859 26960 3911
rect 27472 3859 27478 3911
rect 27530 3899 27536 3911
rect 28912 3899 28918 3911
rect 27530 3871 28918 3899
rect 27530 3859 27536 3871
rect 28912 3859 28918 3871
rect 28970 3859 28976 3911
rect 29008 3859 29014 3911
rect 29066 3899 29072 3911
rect 30352 3899 30358 3911
rect 29066 3871 30358 3899
rect 29066 3859 29072 3871
rect 30352 3859 30358 3871
rect 30410 3859 30416 3911
rect 30736 3859 30742 3911
rect 30794 3899 30800 3911
rect 31984 3899 31990 3911
rect 30794 3871 31990 3899
rect 30794 3859 30800 3871
rect 31984 3859 31990 3871
rect 32042 3859 32048 3911
rect 33424 3859 33430 3911
rect 33482 3899 33488 3911
rect 34768 3899 34774 3911
rect 33482 3871 34774 3899
rect 33482 3859 33488 3871
rect 34768 3859 34774 3871
rect 34826 3859 34832 3911
rect 37072 3859 37078 3911
rect 37130 3899 37136 3911
rect 38608 3899 38614 3911
rect 37130 3871 38614 3899
rect 37130 3859 37136 3871
rect 38608 3859 38614 3871
rect 38666 3859 38672 3911
rect 39664 3859 39670 3911
rect 39722 3899 39728 3911
rect 40912 3899 40918 3911
rect 39722 3871 40918 3899
rect 39722 3859 39728 3871
rect 40912 3859 40918 3871
rect 40970 3859 40976 3911
rect 41104 3859 41110 3911
rect 41162 3899 41168 3911
rect 42064 3899 42070 3911
rect 41162 3871 42070 3899
rect 41162 3859 41168 3871
rect 42064 3859 42070 3871
rect 42122 3859 42128 3911
rect 43312 3859 43318 3911
rect 43370 3899 43376 3911
rect 44752 3899 44758 3911
rect 43370 3871 44758 3899
rect 43370 3859 43376 3871
rect 44752 3859 44758 3871
rect 44810 3859 44816 3911
rect 44848 3859 44854 3911
rect 44906 3899 44912 3911
rect 46192 3899 46198 3911
rect 44906 3871 46198 3899
rect 44906 3859 44912 3871
rect 46192 3859 46198 3871
rect 46250 3859 46256 3911
rect 46288 3859 46294 3911
rect 46346 3899 46352 3911
rect 47632 3899 47638 3911
rect 46346 3871 47638 3899
rect 46346 3859 46352 3871
rect 47632 3859 47638 3871
rect 47690 3859 47696 3911
rect 48496 3859 48502 3911
rect 48554 3899 48560 3911
rect 49648 3899 49654 3911
rect 48554 3871 49654 3899
rect 48554 3859 48560 3871
rect 49648 3859 49654 3871
rect 49706 3859 49712 3911
rect 51376 3859 51382 3911
rect 51434 3899 51440 3911
rect 51856 3899 51862 3911
rect 51434 3871 51862 3899
rect 51434 3859 51440 3871
rect 51856 3859 51862 3871
rect 51914 3859 51920 3911
rect 56272 3859 56278 3911
rect 56330 3899 56336 3911
rect 56330 3871 57614 3899
rect 56330 3859 56336 3871
rect 18928 3825 18934 3837
rect 10675 3788 10733 3794
rect 10786 3797 11006 3825
rect 16450 3797 18934 3825
rect 2992 3711 2998 3763
rect 3050 3751 3056 3763
rect 3280 3751 3286 3763
rect 3050 3723 3286 3751
rect 3050 3711 3056 3723
rect 3280 3711 3286 3723
rect 3338 3711 3344 3763
rect 3376 3711 3382 3763
rect 3434 3751 3440 3763
rect 10786 3751 10814 3797
rect 3434 3723 4670 3751
rect 3434 3711 3440 3723
rect 112 3637 118 3689
rect 170 3677 176 3689
rect 1555 3680 1613 3686
rect 1555 3677 1567 3680
rect 170 3649 1567 3677
rect 170 3637 176 3649
rect 1555 3646 1567 3649
rect 1601 3646 1613 3680
rect 1555 3640 1613 3646
rect 1648 3637 1654 3689
rect 1706 3677 1712 3689
rect 2323 3680 2381 3686
rect 2323 3677 2335 3680
rect 1706 3649 2335 3677
rect 1706 3637 1712 3649
rect 2323 3646 2335 3649
rect 2369 3646 2381 3680
rect 2323 3640 2381 3646
rect 2704 3637 2710 3689
rect 2762 3677 2768 3689
rect 4642 3686 4670 3723
rect 10498 3723 10814 3751
rect 10978 3751 11006 3797
rect 18928 3785 18934 3797
rect 18986 3785 18992 3837
rect 24211 3828 24269 3834
rect 24211 3794 24223 3828
rect 24257 3825 24269 3828
rect 24257 3797 34526 3825
rect 24257 3794 24269 3797
rect 24211 3788 24269 3794
rect 15475 3754 15533 3760
rect 15475 3751 15487 3754
rect 10978 3723 15487 3751
rect 3091 3680 3149 3686
rect 3091 3677 3103 3680
rect 2762 3649 3103 3677
rect 2762 3637 2768 3649
rect 3091 3646 3103 3649
rect 3137 3646 3149 3680
rect 3091 3640 3149 3646
rect 3859 3680 3917 3686
rect 3859 3646 3871 3680
rect 3905 3646 3917 3680
rect 3859 3640 3917 3646
rect 4627 3680 4685 3686
rect 4627 3646 4639 3680
rect 4673 3646 4685 3680
rect 5584 3677 5590 3689
rect 5545 3649 5590 3677
rect 4627 3640 4685 3646
rect 208 3563 214 3615
rect 266 3603 272 3615
rect 1744 3603 1750 3615
rect 266 3575 1750 3603
rect 266 3563 272 3575
rect 1744 3563 1750 3575
rect 1802 3563 1808 3615
rect 592 3489 598 3541
rect 650 3529 656 3541
rect 1456 3529 1462 3541
rect 650 3501 1462 3529
rect 650 3489 656 3501
rect 1456 3489 1462 3501
rect 1514 3489 1520 3541
rect 3088 3489 3094 3541
rect 3146 3529 3152 3541
rect 3874 3529 3902 3640
rect 5584 3637 5590 3649
rect 5642 3637 5648 3689
rect 6352 3637 6358 3689
rect 6410 3677 6416 3689
rect 6931 3680 6989 3686
rect 6931 3677 6943 3680
rect 6410 3649 6943 3677
rect 6410 3637 6416 3649
rect 6931 3646 6943 3649
rect 6977 3646 6989 3680
rect 6931 3640 6989 3646
rect 7024 3637 7030 3689
rect 7082 3677 7088 3689
rect 7699 3680 7757 3686
rect 7699 3677 7711 3680
rect 7082 3649 7711 3677
rect 7082 3637 7088 3649
rect 7699 3646 7711 3649
rect 7745 3646 7757 3680
rect 7699 3640 7757 3646
rect 7792 3637 7798 3689
rect 7850 3677 7856 3689
rect 8467 3680 8525 3686
rect 8467 3677 8479 3680
rect 7850 3649 8479 3677
rect 7850 3637 7856 3649
rect 8467 3646 8479 3649
rect 8513 3646 8525 3680
rect 8467 3640 8525 3646
rect 8560 3637 8566 3689
rect 8618 3677 8624 3689
rect 9235 3680 9293 3686
rect 9235 3677 9247 3680
rect 8618 3649 9247 3677
rect 8618 3637 8624 3649
rect 9235 3646 9247 3649
rect 9281 3646 9293 3680
rect 9235 3640 9293 3646
rect 9328 3637 9334 3689
rect 9386 3677 9392 3689
rect 10003 3680 10061 3686
rect 10003 3677 10015 3680
rect 9386 3649 10015 3677
rect 9386 3637 9392 3649
rect 10003 3646 10015 3649
rect 10049 3646 10061 3680
rect 10003 3640 10061 3646
rect 7984 3563 7990 3615
rect 8042 3603 8048 3615
rect 10498 3603 10526 3723
rect 15475 3720 15487 3723
rect 15521 3720 15533 3754
rect 15475 3714 15533 3720
rect 20464 3711 20470 3763
rect 20522 3751 20528 3763
rect 20848 3751 20854 3763
rect 20522 3723 20854 3751
rect 20522 3711 20528 3723
rect 20848 3711 20854 3723
rect 20906 3711 20912 3763
rect 25168 3711 25174 3763
rect 25226 3751 25232 3763
rect 26320 3751 26326 3763
rect 25226 3723 26326 3751
rect 25226 3711 25232 3723
rect 26320 3711 26326 3723
rect 26378 3711 26384 3763
rect 27376 3711 27382 3763
rect 27434 3751 27440 3763
rect 28432 3751 28438 3763
rect 27434 3723 28438 3751
rect 27434 3711 27440 3723
rect 28432 3711 28438 3723
rect 28490 3711 28496 3763
rect 28720 3711 28726 3763
rect 28778 3751 28784 3763
rect 34498 3751 34526 3797
rect 34672 3785 34678 3837
rect 34730 3825 34736 3837
rect 35440 3825 35446 3837
rect 34730 3797 35446 3825
rect 34730 3785 34736 3797
rect 35440 3785 35446 3797
rect 35498 3785 35504 3837
rect 35632 3785 35638 3837
rect 35690 3825 35696 3837
rect 36496 3825 36502 3837
rect 35690 3797 36502 3825
rect 35690 3785 35696 3797
rect 36496 3785 36502 3797
rect 36554 3785 36560 3837
rect 37840 3785 37846 3837
rect 37898 3825 37904 3837
rect 39376 3825 39382 3837
rect 37898 3797 39382 3825
rect 37898 3785 37904 3797
rect 39376 3785 39382 3797
rect 39434 3785 39440 3837
rect 39952 3785 39958 3837
rect 40010 3825 40016 3837
rect 41008 3825 41014 3837
rect 40010 3797 41014 3825
rect 40010 3785 40016 3797
rect 41008 3785 41014 3797
rect 41066 3785 41072 3837
rect 44080 3785 44086 3837
rect 44138 3825 44144 3837
rect 45424 3825 45430 3837
rect 44138 3797 45430 3825
rect 44138 3785 44144 3797
rect 45424 3785 45430 3797
rect 45482 3785 45488 3837
rect 56752 3785 56758 3837
rect 56810 3785 56816 3837
rect 57586 3825 57614 3871
rect 59440 3825 59446 3837
rect 57586 3797 59446 3825
rect 59440 3785 59446 3797
rect 59498 3785 59504 3837
rect 36688 3751 36694 3763
rect 28778 3723 29630 3751
rect 34498 3723 36694 3751
rect 28778 3711 28784 3723
rect 10576 3637 10582 3689
rect 10634 3677 10640 3689
rect 10771 3680 10829 3686
rect 10771 3677 10783 3680
rect 10634 3649 10783 3677
rect 10634 3637 10640 3649
rect 10771 3646 10783 3649
rect 10817 3646 10829 3680
rect 10771 3640 10829 3646
rect 12979 3680 13037 3686
rect 12979 3646 12991 3680
rect 13025 3677 13037 3680
rect 13168 3677 13174 3689
rect 13025 3649 13174 3677
rect 13025 3646 13037 3649
rect 12979 3640 13037 3646
rect 13168 3637 13174 3649
rect 13226 3637 13232 3689
rect 13648 3677 13654 3689
rect 13609 3649 13654 3677
rect 13648 3637 13654 3649
rect 13706 3637 13712 3689
rect 14032 3637 14038 3689
rect 14090 3677 14096 3689
rect 14419 3680 14477 3686
rect 14419 3677 14431 3680
rect 14090 3649 14431 3677
rect 14090 3637 14096 3649
rect 14419 3646 14431 3649
rect 14465 3646 14477 3680
rect 14419 3640 14477 3646
rect 14800 3637 14806 3689
rect 14858 3677 14864 3689
rect 15187 3680 15245 3686
rect 15187 3677 15199 3680
rect 14858 3649 15199 3677
rect 14858 3637 14864 3649
rect 15187 3646 15199 3649
rect 15233 3646 15245 3680
rect 15187 3640 15245 3646
rect 15280 3637 15286 3689
rect 15338 3677 15344 3689
rect 15955 3680 16013 3686
rect 15955 3677 15967 3680
rect 15338 3649 15967 3677
rect 15338 3637 15344 3649
rect 15955 3646 15967 3649
rect 16001 3646 16013 3680
rect 15955 3640 16013 3646
rect 17392 3637 17398 3689
rect 17450 3677 17456 3689
rect 17491 3680 17549 3686
rect 17491 3677 17503 3680
rect 17450 3649 17503 3677
rect 17450 3637 17456 3649
rect 17491 3646 17503 3649
rect 17537 3646 17549 3680
rect 17491 3640 17549 3646
rect 18064 3637 18070 3689
rect 18122 3677 18128 3689
rect 18259 3680 18317 3686
rect 18259 3677 18271 3680
rect 18122 3649 18271 3677
rect 18122 3637 18128 3649
rect 18259 3646 18271 3649
rect 18305 3646 18317 3680
rect 18259 3640 18317 3646
rect 18448 3637 18454 3689
rect 18506 3677 18512 3689
rect 19027 3680 19085 3686
rect 19027 3677 19039 3680
rect 18506 3649 19039 3677
rect 18506 3637 18512 3649
rect 19027 3646 19039 3649
rect 19073 3646 19085 3680
rect 19027 3640 19085 3646
rect 19216 3637 19222 3689
rect 19274 3677 19280 3689
rect 19795 3680 19853 3686
rect 19795 3677 19807 3680
rect 19274 3649 19807 3677
rect 19274 3637 19280 3649
rect 19795 3646 19807 3649
rect 19841 3646 19853 3680
rect 19795 3640 19853 3646
rect 19984 3637 19990 3689
rect 20042 3677 20048 3689
rect 20563 3680 20621 3686
rect 20563 3677 20575 3680
rect 20042 3649 20575 3677
rect 20042 3637 20048 3649
rect 20563 3646 20575 3649
rect 20609 3646 20621 3680
rect 20563 3640 20621 3646
rect 20656 3637 20662 3689
rect 20714 3677 20720 3689
rect 21331 3680 21389 3686
rect 21331 3677 21343 3680
rect 20714 3649 21343 3677
rect 20714 3637 20720 3649
rect 21331 3646 21343 3649
rect 21377 3646 21389 3680
rect 21331 3640 21389 3646
rect 22096 3637 22102 3689
rect 22154 3677 22160 3689
rect 22771 3680 22829 3686
rect 22771 3677 22783 3680
rect 22154 3649 22783 3677
rect 22154 3637 22160 3649
rect 22771 3646 22783 3649
rect 22817 3646 22829 3680
rect 22771 3640 22829 3646
rect 22864 3637 22870 3689
rect 22922 3677 22928 3689
rect 23539 3680 23597 3686
rect 23539 3677 23551 3680
rect 22922 3649 23551 3677
rect 22922 3637 22928 3649
rect 23539 3646 23551 3649
rect 23585 3646 23597 3680
rect 23539 3640 23597 3646
rect 23632 3637 23638 3689
rect 23690 3677 23696 3689
rect 24307 3680 24365 3686
rect 24307 3677 24319 3680
rect 23690 3649 24319 3677
rect 23690 3637 23696 3649
rect 24307 3646 24319 3649
rect 24353 3646 24365 3680
rect 24307 3640 24365 3646
rect 24400 3637 24406 3689
rect 24458 3677 24464 3689
rect 25075 3680 25133 3686
rect 25075 3677 25087 3680
rect 24458 3649 25087 3677
rect 24458 3637 24464 3649
rect 25075 3646 25087 3649
rect 25121 3646 25133 3680
rect 25075 3640 25133 3646
rect 25843 3680 25901 3686
rect 25843 3646 25855 3680
rect 25889 3646 25901 3680
rect 25843 3640 25901 3646
rect 26611 3680 26669 3686
rect 26611 3646 26623 3680
rect 26657 3646 26669 3680
rect 26611 3640 26669 3646
rect 8042 3575 10526 3603
rect 10675 3606 10733 3612
rect 8042 3563 8048 3575
rect 10675 3572 10687 3606
rect 10721 3572 10733 3606
rect 10675 3566 10733 3572
rect 12403 3606 12461 3612
rect 12403 3572 12415 3606
rect 12449 3603 12461 3606
rect 24211 3606 24269 3612
rect 24211 3603 24223 3606
rect 12449 3575 24223 3603
rect 12449 3572 12461 3575
rect 12403 3566 12461 3572
rect 24211 3572 24223 3575
rect 24257 3572 24269 3606
rect 24211 3566 24269 3572
rect 3146 3501 3902 3529
rect 3146 3489 3152 3501
rect 10000 3489 10006 3541
rect 10058 3529 10064 3541
rect 10576 3529 10582 3541
rect 10058 3501 10582 3529
rect 10058 3489 10064 3501
rect 10576 3489 10582 3501
rect 10634 3489 10640 3541
rect 10690 3529 10718 3566
rect 24688 3563 24694 3615
rect 24746 3603 24752 3615
rect 25858 3603 25886 3640
rect 24746 3575 25886 3603
rect 24746 3563 24752 3575
rect 14707 3532 14765 3538
rect 14707 3529 14719 3532
rect 10690 3501 14719 3529
rect 14707 3498 14719 3501
rect 14753 3498 14765 3532
rect 14707 3492 14765 3498
rect 19024 3489 19030 3541
rect 19082 3529 19088 3541
rect 19504 3529 19510 3541
rect 19082 3501 19510 3529
rect 19082 3489 19088 3501
rect 19504 3489 19510 3501
rect 19562 3489 19568 3541
rect 25840 3489 25846 3541
rect 25898 3529 25904 3541
rect 26626 3529 26654 3640
rect 27280 3637 27286 3689
rect 27338 3677 27344 3689
rect 29602 3686 29630 3723
rect 36688 3711 36694 3723
rect 36746 3711 36752 3763
rect 41296 3711 41302 3763
rect 41354 3751 41360 3763
rect 41584 3751 41590 3763
rect 41354 3723 41590 3751
rect 41354 3711 41360 3723
rect 41584 3711 41590 3723
rect 41642 3711 41648 3763
rect 45232 3711 45238 3763
rect 45290 3751 45296 3763
rect 45290 3723 46238 3751
rect 45290 3711 45296 3723
rect 28051 3680 28109 3686
rect 28051 3677 28063 3680
rect 27338 3649 28063 3677
rect 27338 3637 27344 3649
rect 28051 3646 28063 3649
rect 28097 3646 28109 3680
rect 28051 3640 28109 3646
rect 28819 3680 28877 3686
rect 28819 3646 28831 3680
rect 28865 3646 28877 3680
rect 28819 3640 28877 3646
rect 29587 3680 29645 3686
rect 29587 3646 29599 3680
rect 29633 3646 29645 3680
rect 29587 3640 29645 3646
rect 30355 3680 30413 3686
rect 30355 3646 30367 3680
rect 30401 3646 30413 3680
rect 30355 3640 30413 3646
rect 25898 3501 26654 3529
rect 25898 3489 25904 3501
rect 28048 3489 28054 3541
rect 28106 3529 28112 3541
rect 28834 3529 28862 3640
rect 29488 3563 29494 3615
rect 29546 3603 29552 3615
rect 30370 3603 30398 3640
rect 30448 3637 30454 3689
rect 30506 3677 30512 3689
rect 31123 3680 31181 3686
rect 31123 3677 31135 3680
rect 30506 3649 31135 3677
rect 30506 3637 30512 3649
rect 31123 3646 31135 3649
rect 31169 3646 31181 3680
rect 31123 3640 31181 3646
rect 31312 3637 31318 3689
rect 31370 3677 31376 3689
rect 31891 3680 31949 3686
rect 31891 3677 31903 3680
rect 31370 3649 31903 3677
rect 31370 3637 31376 3649
rect 31891 3646 31903 3649
rect 31937 3646 31949 3680
rect 31891 3640 31949 3646
rect 32464 3637 32470 3689
rect 32522 3677 32528 3689
rect 33331 3680 33389 3686
rect 33331 3677 33343 3680
rect 32522 3649 33343 3677
rect 32522 3637 32528 3649
rect 33331 3646 33343 3649
rect 33377 3646 33389 3680
rect 33331 3640 33389 3646
rect 33520 3637 33526 3689
rect 33578 3677 33584 3689
rect 34099 3680 34157 3686
rect 34099 3677 34111 3680
rect 33578 3649 34111 3677
rect 33578 3637 33584 3649
rect 34099 3646 34111 3649
rect 34145 3646 34157 3680
rect 34099 3640 34157 3646
rect 34288 3637 34294 3689
rect 34346 3677 34352 3689
rect 34867 3680 34925 3686
rect 34867 3677 34879 3680
rect 34346 3649 34879 3677
rect 34346 3637 34352 3649
rect 34867 3646 34879 3649
rect 34913 3646 34925 3680
rect 34867 3640 34925 3646
rect 35344 3637 35350 3689
rect 35402 3677 35408 3689
rect 35635 3680 35693 3686
rect 35635 3677 35647 3680
rect 35402 3649 35647 3677
rect 35402 3637 35408 3649
rect 35635 3646 35647 3649
rect 35681 3646 35693 3680
rect 35635 3640 35693 3646
rect 35728 3637 35734 3689
rect 35786 3677 35792 3689
rect 36403 3680 36461 3686
rect 36403 3677 36415 3680
rect 35786 3649 36415 3677
rect 35786 3637 35792 3649
rect 36403 3646 36415 3649
rect 36449 3646 36461 3680
rect 36403 3640 36461 3646
rect 36496 3637 36502 3689
rect 36554 3677 36560 3689
rect 37171 3680 37229 3686
rect 37171 3677 37183 3680
rect 36554 3649 37183 3677
rect 36554 3637 36560 3649
rect 37171 3646 37183 3649
rect 37217 3646 37229 3680
rect 37171 3640 37229 3646
rect 37936 3637 37942 3689
rect 37994 3677 38000 3689
rect 38611 3680 38669 3686
rect 38611 3677 38623 3680
rect 37994 3649 38623 3677
rect 37994 3637 38000 3649
rect 38611 3646 38623 3649
rect 38657 3646 38669 3680
rect 38611 3640 38669 3646
rect 38704 3637 38710 3689
rect 38762 3677 38768 3689
rect 39379 3680 39437 3686
rect 39379 3677 39391 3680
rect 38762 3649 39391 3677
rect 38762 3637 38768 3649
rect 39379 3646 39391 3649
rect 39425 3646 39437 3680
rect 39379 3640 39437 3646
rect 39472 3637 39478 3689
rect 39530 3677 39536 3689
rect 40147 3680 40205 3686
rect 40147 3677 40159 3680
rect 39530 3649 40159 3677
rect 39530 3637 39536 3649
rect 40147 3646 40159 3649
rect 40193 3646 40205 3680
rect 40147 3640 40205 3646
rect 40240 3637 40246 3689
rect 40298 3677 40304 3689
rect 40915 3680 40973 3686
rect 40915 3677 40927 3680
rect 40298 3649 40927 3677
rect 40298 3637 40304 3649
rect 40915 3646 40927 3649
rect 40961 3646 40973 3680
rect 40915 3640 40973 3646
rect 41008 3637 41014 3689
rect 41066 3677 41072 3689
rect 41683 3680 41741 3686
rect 41683 3677 41695 3680
rect 41066 3649 41695 3677
rect 41066 3637 41072 3649
rect 41683 3646 41695 3649
rect 41729 3646 41741 3680
rect 41683 3640 41741 3646
rect 42451 3680 42509 3686
rect 42451 3646 42463 3680
rect 42497 3646 42509 3680
rect 42451 3640 42509 3646
rect 29546 3575 30398 3603
rect 29546 3563 29552 3575
rect 36688 3563 36694 3615
rect 36746 3603 36752 3615
rect 37552 3603 37558 3615
rect 36746 3575 37558 3603
rect 36746 3563 36752 3575
rect 37552 3563 37558 3575
rect 37610 3563 37616 3615
rect 41584 3563 41590 3615
rect 41642 3603 41648 3615
rect 42466 3603 42494 3640
rect 42736 3637 42742 3689
rect 42794 3677 42800 3689
rect 46210 3686 46238 3723
rect 47536 3711 47542 3763
rect 47594 3751 47600 3763
rect 48304 3751 48310 3763
rect 47594 3723 48310 3751
rect 47594 3711 47600 3723
rect 48304 3711 48310 3723
rect 48362 3711 48368 3763
rect 55888 3711 55894 3763
rect 55946 3751 55952 3763
rect 56770 3751 56798 3785
rect 59152 3751 59158 3763
rect 55946 3723 56126 3751
rect 56770 3723 59158 3751
rect 55946 3711 55952 3723
rect 43891 3680 43949 3686
rect 43891 3677 43903 3680
rect 42794 3649 43903 3677
rect 42794 3637 42800 3649
rect 43891 3646 43903 3649
rect 43937 3646 43949 3680
rect 43891 3640 43949 3646
rect 44659 3680 44717 3686
rect 44659 3646 44671 3680
rect 44705 3646 44717 3680
rect 44659 3640 44717 3646
rect 45427 3680 45485 3686
rect 45427 3646 45439 3680
rect 45473 3646 45485 3680
rect 45427 3640 45485 3646
rect 46195 3680 46253 3686
rect 46195 3646 46207 3680
rect 46241 3646 46253 3680
rect 46195 3640 46253 3646
rect 46963 3680 47021 3686
rect 46963 3646 46975 3680
rect 47009 3646 47021 3680
rect 46963 3640 47021 3646
rect 41642 3575 42494 3603
rect 41642 3563 41648 3575
rect 43792 3563 43798 3615
rect 43850 3603 43856 3615
rect 44674 3603 44702 3640
rect 43850 3575 44702 3603
rect 43850 3563 43856 3575
rect 28106 3501 28862 3529
rect 28106 3489 28112 3501
rect 30448 3489 30454 3541
rect 30506 3529 30512 3541
rect 31888 3529 31894 3541
rect 30506 3501 31894 3529
rect 30506 3489 30512 3501
rect 31888 3489 31894 3501
rect 31946 3489 31952 3541
rect 44560 3489 44566 3541
rect 44618 3529 44624 3541
rect 45442 3529 45470 3640
rect 46000 3563 46006 3615
rect 46058 3603 46064 3615
rect 46978 3603 47006 3640
rect 47152 3637 47158 3689
rect 47210 3677 47216 3689
rect 47731 3680 47789 3686
rect 47731 3677 47743 3680
rect 47210 3649 47743 3677
rect 47210 3637 47216 3649
rect 47731 3646 47743 3649
rect 47777 3646 47789 3680
rect 47731 3640 47789 3646
rect 48208 3637 48214 3689
rect 48266 3677 48272 3689
rect 49171 3680 49229 3686
rect 49171 3677 49183 3680
rect 48266 3649 49183 3677
rect 48266 3637 48272 3649
rect 49171 3646 49183 3649
rect 49217 3646 49229 3680
rect 49171 3640 49229 3646
rect 50515 3680 50573 3686
rect 50515 3646 50527 3680
rect 50561 3677 50573 3680
rect 50704 3677 50710 3689
rect 50561 3649 50710 3677
rect 50561 3646 50573 3649
rect 50515 3640 50573 3646
rect 50704 3637 50710 3649
rect 50762 3637 50768 3689
rect 50800 3637 50806 3689
rect 50858 3677 50864 3689
rect 51187 3680 51245 3686
rect 51187 3677 51199 3680
rect 50858 3649 51199 3677
rect 50858 3637 50864 3649
rect 51187 3646 51199 3649
rect 51233 3646 51245 3680
rect 51187 3640 51245 3646
rect 51280 3637 51286 3689
rect 51338 3677 51344 3689
rect 51955 3680 52013 3686
rect 51955 3677 51967 3680
rect 51338 3649 51967 3677
rect 51338 3637 51344 3649
rect 51955 3646 51967 3649
rect 52001 3646 52013 3680
rect 51955 3640 52013 3646
rect 52048 3637 52054 3689
rect 52106 3677 52112 3689
rect 52723 3680 52781 3686
rect 52723 3677 52735 3680
rect 52106 3649 52735 3677
rect 52106 3637 52112 3649
rect 52723 3646 52735 3649
rect 52769 3646 52781 3680
rect 52723 3640 52781 3646
rect 53392 3637 53398 3689
rect 53450 3677 53456 3689
rect 54451 3680 54509 3686
rect 54451 3677 54463 3680
rect 53450 3649 54463 3677
rect 53450 3637 53456 3649
rect 54451 3646 54463 3649
rect 54497 3646 54509 3680
rect 54451 3640 54509 3646
rect 55219 3680 55277 3686
rect 55219 3646 55231 3680
rect 55265 3646 55277 3680
rect 55219 3640 55277 3646
rect 55987 3680 56045 3686
rect 55987 3646 55999 3680
rect 56033 3646 56045 3680
rect 56098 3677 56126 3723
rect 59152 3711 59158 3723
rect 59210 3711 59216 3763
rect 56755 3680 56813 3686
rect 56755 3677 56767 3680
rect 56098 3649 56767 3677
rect 55987 3640 56045 3646
rect 56755 3646 56767 3649
rect 56801 3646 56813 3680
rect 56755 3640 56813 3646
rect 57523 3680 57581 3686
rect 57523 3646 57535 3680
rect 57569 3646 57581 3680
rect 57523 3640 57581 3646
rect 46058 3575 47006 3603
rect 46058 3563 46064 3575
rect 44618 3501 45470 3529
rect 44618 3489 44624 3501
rect 45712 3489 45718 3541
rect 45770 3529 45776 3541
rect 46384 3529 46390 3541
rect 45770 3501 46390 3529
rect 45770 3489 45776 3501
rect 46384 3489 46390 3501
rect 46442 3489 46448 3541
rect 49072 3489 49078 3541
rect 49130 3529 49136 3541
rect 50032 3529 50038 3541
rect 49130 3501 50038 3529
rect 49130 3489 49136 3501
rect 50032 3489 50038 3501
rect 50090 3489 50096 3541
rect 51280 3489 51286 3541
rect 51338 3529 51344 3541
rect 51472 3529 51478 3541
rect 51338 3501 51478 3529
rect 51338 3489 51344 3501
rect 51472 3489 51478 3501
rect 51530 3489 51536 3541
rect 52048 3489 52054 3541
rect 52106 3529 52112 3541
rect 52720 3529 52726 3541
rect 52106 3501 52726 3529
rect 52106 3489 52112 3501
rect 52720 3489 52726 3501
rect 52778 3489 52784 3541
rect 54448 3489 54454 3541
rect 54506 3529 54512 3541
rect 55234 3529 55262 3640
rect 54506 3501 55262 3529
rect 54506 3489 54512 3501
rect 3280 3415 3286 3467
rect 3338 3455 3344 3467
rect 3952 3455 3958 3467
rect 3338 3427 3958 3455
rect 3338 3415 3344 3427
rect 3952 3415 3958 3427
rect 4010 3415 4016 3467
rect 7504 3415 7510 3467
rect 7562 3455 7568 3467
rect 11920 3455 11926 3467
rect 7562 3427 11926 3455
rect 7562 3415 7568 3427
rect 11920 3415 11926 3427
rect 11978 3415 11984 3467
rect 12016 3415 12022 3467
rect 12074 3455 12080 3467
rect 13360 3455 13366 3467
rect 12074 3427 13366 3455
rect 12074 3415 12080 3427
rect 13360 3415 13366 3427
rect 13418 3415 13424 3467
rect 14224 3415 14230 3467
rect 14282 3455 14288 3467
rect 17779 3458 17837 3464
rect 17779 3455 17791 3458
rect 14282 3427 17791 3455
rect 14282 3415 14288 3427
rect 17779 3424 17791 3427
rect 17825 3424 17837 3458
rect 20848 3455 20854 3467
rect 20809 3427 20854 3455
rect 17779 3418 17837 3424
rect 20848 3415 20854 3427
rect 20906 3415 20912 3467
rect 26320 3415 26326 3467
rect 26378 3455 26384 3467
rect 27568 3455 27574 3467
rect 26378 3427 27574 3455
rect 26378 3415 26384 3427
rect 27568 3415 27574 3427
rect 27626 3415 27632 3467
rect 28912 3415 28918 3467
rect 28970 3455 28976 3467
rect 29776 3455 29782 3467
rect 28970 3427 29782 3455
rect 28970 3415 28976 3427
rect 29776 3415 29782 3427
rect 29834 3415 29840 3467
rect 32560 3415 32566 3467
rect 32618 3455 32624 3467
rect 33712 3455 33718 3467
rect 32618 3427 33718 3455
rect 32618 3415 32624 3427
rect 33712 3415 33718 3427
rect 33770 3415 33776 3467
rect 45424 3415 45430 3467
rect 45482 3455 45488 3467
rect 45616 3455 45622 3467
rect 45482 3427 45622 3455
rect 45482 3415 45488 3427
rect 45616 3415 45622 3427
rect 45674 3415 45680 3467
rect 55216 3415 55222 3467
rect 55274 3455 55280 3467
rect 56002 3455 56030 3640
rect 56560 3563 56566 3615
rect 56618 3603 56624 3615
rect 56848 3603 56854 3615
rect 56618 3575 56854 3603
rect 56618 3563 56624 3575
rect 56848 3563 56854 3575
rect 56906 3563 56912 3615
rect 56272 3489 56278 3541
rect 56330 3529 56336 3541
rect 57538 3529 57566 3640
rect 58192 3637 58198 3689
rect 58250 3677 58256 3689
rect 59728 3677 59734 3689
rect 58250 3649 59734 3677
rect 58250 3637 58256 3649
rect 59728 3637 59734 3649
rect 59786 3637 59792 3689
rect 56330 3501 57566 3529
rect 56330 3489 56336 3501
rect 55274 3427 56030 3455
rect 55274 3415 55280 3427
rect 1152 3356 58848 3378
rect 1152 3304 19654 3356
rect 19706 3304 19718 3356
rect 19770 3304 19782 3356
rect 19834 3304 19846 3356
rect 19898 3304 50374 3356
rect 50426 3304 50438 3356
rect 50490 3304 50502 3356
rect 50554 3304 50566 3356
rect 50618 3304 58848 3356
rect 1152 3282 58848 3304
rect 1456 3193 1462 3245
rect 1514 3233 1520 3245
rect 2128 3233 2134 3245
rect 1514 3205 2134 3233
rect 1514 3193 1520 3205
rect 2128 3193 2134 3205
rect 2186 3193 2192 3245
rect 3952 3193 3958 3245
rect 4010 3233 4016 3245
rect 5200 3233 5206 3245
rect 4010 3205 5206 3233
rect 4010 3193 4016 3205
rect 5200 3193 5206 3205
rect 5258 3193 5264 3245
rect 8176 3193 8182 3245
rect 8234 3233 8240 3245
rect 12691 3236 12749 3242
rect 12691 3233 12703 3236
rect 8234 3205 12703 3233
rect 8234 3193 8240 3205
rect 12691 3202 12703 3205
rect 12737 3202 12749 3236
rect 12691 3196 12749 3202
rect 12802 3205 13406 3233
rect 7120 3119 7126 3171
rect 7178 3159 7184 3171
rect 12802 3159 12830 3205
rect 7178 3131 12830 3159
rect 7178 3119 7184 3131
rect 13072 3119 13078 3171
rect 13130 3159 13136 3171
rect 13267 3162 13325 3168
rect 13267 3159 13279 3162
rect 13130 3131 13279 3159
rect 13130 3119 13136 3131
rect 13267 3128 13279 3131
rect 13313 3128 13325 3162
rect 13378 3159 13406 3205
rect 13744 3193 13750 3245
rect 13802 3233 13808 3245
rect 14035 3236 14093 3242
rect 14035 3233 14047 3236
rect 13802 3205 14047 3233
rect 13802 3193 13808 3205
rect 14035 3202 14047 3205
rect 14081 3202 14093 3236
rect 15379 3236 15437 3242
rect 15379 3233 15391 3236
rect 14035 3196 14093 3202
rect 14146 3205 15391 3233
rect 14146 3159 14174 3205
rect 15379 3202 15391 3205
rect 15425 3202 15437 3236
rect 16816 3233 16822 3245
rect 16777 3205 16822 3233
rect 15379 3196 15437 3202
rect 16816 3193 16822 3205
rect 16874 3193 16880 3245
rect 18928 3193 18934 3245
rect 18986 3233 18992 3245
rect 19123 3236 19181 3242
rect 19123 3233 19135 3236
rect 18986 3205 19135 3233
rect 18986 3193 18992 3205
rect 19123 3202 19135 3205
rect 19169 3233 19181 3236
rect 19315 3236 19373 3242
rect 19315 3233 19327 3236
rect 19169 3205 19327 3233
rect 19169 3202 19181 3205
rect 19123 3196 19181 3202
rect 19315 3202 19327 3205
rect 19361 3202 19373 3236
rect 19315 3196 19373 3202
rect 19696 3193 19702 3245
rect 19754 3233 19760 3245
rect 20368 3233 20374 3245
rect 19754 3205 20374 3233
rect 19754 3193 19760 3205
rect 20368 3193 20374 3205
rect 20426 3193 20432 3245
rect 20944 3193 20950 3245
rect 21002 3233 21008 3245
rect 21712 3233 21718 3245
rect 21002 3205 21718 3233
rect 21002 3193 21008 3205
rect 21712 3193 21718 3205
rect 21770 3193 21776 3245
rect 22000 3193 22006 3245
rect 22058 3233 22064 3245
rect 24016 3233 24022 3245
rect 22058 3205 24022 3233
rect 22058 3193 22064 3205
rect 24016 3193 24022 3205
rect 24074 3193 24080 3245
rect 24976 3193 24982 3245
rect 25034 3233 25040 3245
rect 26608 3233 26614 3245
rect 25034 3205 26614 3233
rect 25034 3193 25040 3205
rect 26608 3193 26614 3205
rect 26666 3193 26672 3245
rect 32656 3193 32662 3245
rect 32714 3233 32720 3245
rect 34096 3233 34102 3245
rect 32714 3205 34102 3233
rect 32714 3193 32720 3205
rect 34096 3193 34102 3205
rect 34154 3193 34160 3245
rect 40048 3193 40054 3245
rect 40106 3233 40112 3245
rect 40240 3233 40246 3245
rect 40106 3205 40246 3233
rect 40106 3193 40112 3205
rect 40240 3193 40246 3205
rect 40298 3193 40304 3245
rect 41200 3193 41206 3245
rect 41258 3233 41264 3245
rect 48499 3236 48557 3242
rect 48499 3233 48511 3236
rect 41258 3205 48511 3233
rect 41258 3193 41264 3205
rect 48499 3202 48511 3205
rect 48545 3202 48557 3236
rect 48499 3196 48557 3202
rect 56368 3193 56374 3245
rect 56426 3233 56432 3245
rect 58000 3233 58006 3245
rect 56426 3205 58006 3233
rect 56426 3193 56432 3205
rect 58000 3193 58006 3205
rect 58058 3193 58064 3245
rect 18835 3162 18893 3168
rect 18835 3159 18847 3162
rect 13378 3131 14174 3159
rect 14914 3131 18847 3159
rect 13267 3122 13325 3128
rect 8944 3045 8950 3097
rect 9002 3085 9008 3097
rect 12691 3088 12749 3094
rect 9002 3057 10814 3085
rect 9002 3045 9008 3057
rect 16 2971 22 3023
rect 74 3011 80 3023
rect 1555 3014 1613 3020
rect 1555 3011 1567 3014
rect 74 2983 1567 3011
rect 74 2971 80 2983
rect 1555 2980 1567 2983
rect 1601 2980 1613 3014
rect 2323 3014 2381 3020
rect 2323 3011 2335 3014
rect 1555 2974 1613 2980
rect 1666 2983 2335 3011
rect 688 2897 694 2949
rect 746 2937 752 2949
rect 1666 2937 1694 2983
rect 2323 2980 2335 2983
rect 2369 2980 2381 3014
rect 3091 3014 3149 3020
rect 3091 3011 3103 3014
rect 2323 2974 2381 2980
rect 2866 2983 3103 3011
rect 746 2909 1694 2937
rect 746 2897 752 2909
rect 2128 2897 2134 2949
rect 2186 2937 2192 2949
rect 2866 2937 2894 2983
rect 3091 2980 3103 2983
rect 3137 2980 3149 3014
rect 4912 3011 4918 3023
rect 4873 2983 4918 3011
rect 3091 2974 3149 2980
rect 4912 2971 4918 2983
rect 4970 2971 4976 3023
rect 5200 2971 5206 3023
rect 5258 3011 5264 3023
rect 5683 3014 5741 3020
rect 5683 3011 5695 3014
rect 5258 2983 5695 3011
rect 5258 2971 5264 2983
rect 5683 2980 5695 2983
rect 5729 2980 5741 3014
rect 5683 2974 5741 2980
rect 5968 2971 5974 3023
rect 6026 3011 6032 3023
rect 7027 3014 7085 3020
rect 7027 3011 7039 3014
rect 6026 2983 7039 3011
rect 6026 2971 6032 2983
rect 7027 2980 7039 2983
rect 7073 2980 7085 3014
rect 7027 2974 7085 2980
rect 7795 3014 7853 3020
rect 7795 2980 7807 3014
rect 7841 2980 7853 3014
rect 7795 2974 7853 2980
rect 5776 2937 5782 2949
rect 2186 2909 2894 2937
rect 5218 2909 5782 2937
rect 2186 2897 2192 2909
rect 5104 2749 5110 2801
rect 5162 2789 5168 2801
rect 5218 2789 5246 2909
rect 5776 2897 5782 2909
rect 5834 2897 5840 2949
rect 6736 2897 6742 2949
rect 6794 2937 6800 2949
rect 7810 2937 7838 2974
rect 8176 2971 8182 3023
rect 8234 3011 8240 3023
rect 9715 3014 9773 3020
rect 9715 3011 9727 3014
rect 8234 2983 9727 3011
rect 8234 2971 8240 2983
rect 9715 2980 9727 2983
rect 9761 2980 9773 3014
rect 9715 2974 9773 2980
rect 10579 3014 10637 3020
rect 10579 2980 10591 3014
rect 10625 2980 10637 3014
rect 10579 2974 10637 2980
rect 6794 2909 7838 2937
rect 6794 2897 6800 2909
rect 8944 2897 8950 2949
rect 9002 2937 9008 2949
rect 10594 2937 10622 2974
rect 9002 2909 10622 2937
rect 10786 2937 10814 3057
rect 12691 3054 12703 3088
rect 12737 3085 12749 3088
rect 14914 3085 14942 3131
rect 18835 3128 18847 3131
rect 18881 3128 18893 3162
rect 18835 3122 18893 3128
rect 19792 3119 19798 3171
rect 19850 3159 19856 3171
rect 20176 3159 20182 3171
rect 19850 3131 20182 3159
rect 19850 3119 19856 3131
rect 20176 3119 20182 3131
rect 20234 3119 20240 3171
rect 20755 3162 20813 3168
rect 20755 3128 20767 3162
rect 20801 3159 20813 3162
rect 21136 3159 21142 3171
rect 20801 3131 21142 3159
rect 20801 3128 20813 3131
rect 20755 3122 20813 3128
rect 21136 3119 21142 3131
rect 21194 3119 21200 3171
rect 21424 3119 21430 3171
rect 21482 3119 21488 3171
rect 22960 3119 22966 3171
rect 23018 3159 23024 3171
rect 24304 3159 24310 3171
rect 23018 3131 24310 3159
rect 23018 3119 23024 3131
rect 24304 3119 24310 3131
rect 24362 3119 24368 3171
rect 35347 3162 35405 3168
rect 35347 3128 35359 3162
rect 35393 3159 35405 3162
rect 35635 3162 35693 3168
rect 35635 3159 35647 3162
rect 35393 3131 35647 3159
rect 35393 3128 35405 3131
rect 35347 3122 35405 3128
rect 35635 3128 35647 3131
rect 35681 3159 35693 3162
rect 40816 3159 40822 3171
rect 35681 3131 40822 3159
rect 35681 3128 35693 3131
rect 35635 3122 35693 3128
rect 40816 3119 40822 3131
rect 40874 3119 40880 3171
rect 42064 3119 42070 3171
rect 42122 3159 42128 3171
rect 44176 3159 44182 3171
rect 42122 3131 44182 3159
rect 42122 3119 42128 3131
rect 44176 3119 44182 3131
rect 44234 3119 44240 3171
rect 12737 3057 14942 3085
rect 12737 3054 12749 3057
rect 12691 3048 12749 3054
rect 15376 3045 15382 3097
rect 15434 3085 15440 3097
rect 16432 3085 16438 3097
rect 15434 3057 16438 3085
rect 15434 3045 15440 3057
rect 16432 3045 16438 3057
rect 16490 3045 16496 3097
rect 19504 3045 19510 3097
rect 19562 3085 19568 3097
rect 21442 3085 21470 3119
rect 19562 3057 21470 3085
rect 19562 3045 19568 3057
rect 22384 3045 22390 3097
rect 22442 3085 22448 3097
rect 23536 3085 23542 3097
rect 22442 3057 23542 3085
rect 22442 3045 22448 3057
rect 23536 3045 23542 3057
rect 23594 3045 23600 3097
rect 31888 3045 31894 3097
rect 31946 3085 31952 3097
rect 33328 3085 33334 3097
rect 31946 3057 33334 3085
rect 31946 3045 31952 3057
rect 33328 3045 33334 3057
rect 33386 3045 33392 3097
rect 42544 3045 42550 3097
rect 42602 3085 42608 3097
rect 43504 3085 43510 3097
rect 42602 3057 43510 3085
rect 42602 3045 42608 3057
rect 43504 3045 43510 3057
rect 43562 3045 43568 3097
rect 46384 3045 46390 3097
rect 46442 3085 46448 3097
rect 51763 3088 51821 3094
rect 46442 3057 48158 3085
rect 46442 3045 46448 3057
rect 12976 2971 12982 3023
rect 13034 3011 13040 3023
rect 13034 2983 13079 3011
rect 13034 2971 13040 2983
rect 13360 2971 13366 3023
rect 13418 3011 13424 3023
rect 13747 3014 13805 3020
rect 13747 3011 13759 3014
rect 13418 2983 13759 3011
rect 13418 2971 13424 2983
rect 13747 2980 13759 2983
rect 13793 2980 13805 3014
rect 13747 2974 13805 2980
rect 14512 2971 14518 3023
rect 14570 3011 14576 3023
rect 15091 3014 15149 3020
rect 15091 3011 15103 3014
rect 14570 2983 15103 3011
rect 14570 2971 14576 2983
rect 15091 2980 15103 2983
rect 15137 2980 15149 3014
rect 16624 3011 16630 3023
rect 16585 2983 16630 3011
rect 15091 2974 15149 2980
rect 16624 2971 16630 2983
rect 16682 2971 16688 3023
rect 17008 2971 17014 3023
rect 17066 3011 17072 3023
rect 17779 3014 17837 3020
rect 17779 3011 17791 3014
rect 17066 2983 17791 3011
rect 17066 2971 17072 2983
rect 17779 2980 17791 2983
rect 17825 2980 17837 3014
rect 17779 2974 17837 2980
rect 18547 3014 18605 3020
rect 18547 2980 18559 3014
rect 18593 2980 18605 3014
rect 18547 2974 18605 2980
rect 14224 2937 14230 2949
rect 10786 2909 14230 2937
rect 9002 2897 9008 2909
rect 14224 2897 14230 2909
rect 14282 2897 14288 2949
rect 17680 2897 17686 2949
rect 17738 2937 17744 2949
rect 18562 2937 18590 2974
rect 18928 2971 18934 3023
rect 18986 3011 18992 3023
rect 20467 3014 20525 3020
rect 20467 3011 20479 3014
rect 18986 2983 20479 3011
rect 18986 2971 18992 2983
rect 20467 2980 20479 2983
rect 20513 2980 20525 3014
rect 21235 3014 21293 3020
rect 21235 3011 21247 3014
rect 20467 2974 20525 2980
rect 20578 2983 21247 3011
rect 17738 2909 18590 2937
rect 17738 2897 17744 2909
rect 19600 2897 19606 2949
rect 19658 2937 19664 2949
rect 20578 2937 20606 2983
rect 21235 2980 21247 2983
rect 21281 2980 21293 3014
rect 21235 2974 21293 2980
rect 21424 2971 21430 3023
rect 21482 3011 21488 3023
rect 23155 3014 23213 3020
rect 23155 3011 23167 3014
rect 21482 2983 23167 3011
rect 21482 2971 21488 2983
rect 23155 2980 23167 2983
rect 23201 2980 23213 3014
rect 23155 2974 23213 2980
rect 23923 3014 23981 3020
rect 23923 2980 23935 3014
rect 23969 2980 23981 3014
rect 23923 2974 23981 2980
rect 19658 2909 20606 2937
rect 19658 2897 19664 2909
rect 21136 2897 21142 2949
rect 21194 2937 21200 2949
rect 21523 2940 21581 2946
rect 21523 2937 21535 2940
rect 21194 2909 21535 2937
rect 21194 2897 21200 2909
rect 21523 2906 21535 2909
rect 21569 2906 21581 2940
rect 21523 2900 21581 2906
rect 22480 2897 22486 2949
rect 22538 2937 22544 2949
rect 23938 2937 23966 2974
rect 24016 2971 24022 3023
rect 24074 3011 24080 3023
rect 25843 3014 25901 3020
rect 25843 3011 25855 3014
rect 24074 2983 25855 3011
rect 24074 2971 24080 2983
rect 25843 2980 25855 2983
rect 25889 2980 25901 3014
rect 25843 2974 25901 2980
rect 26611 3014 26669 3020
rect 26611 2980 26623 3014
rect 26657 2980 26669 3014
rect 26611 2974 26669 2980
rect 22538 2909 23966 2937
rect 22538 2897 22544 2909
rect 25072 2897 25078 2949
rect 25130 2937 25136 2949
rect 26626 2937 26654 2974
rect 26896 2971 26902 3023
rect 26954 3011 26960 3023
rect 28531 3014 28589 3020
rect 28531 3011 28543 3014
rect 26954 2983 28543 3011
rect 26954 2971 26960 2983
rect 28531 2980 28543 2983
rect 28577 2980 28589 3014
rect 28531 2974 28589 2980
rect 29299 3014 29357 3020
rect 29299 2980 29311 3014
rect 29345 2980 29357 3014
rect 29299 2974 29357 2980
rect 25130 2909 26654 2937
rect 25130 2897 25136 2909
rect 27568 2897 27574 2949
rect 27626 2937 27632 2949
rect 29314 2937 29342 2974
rect 29872 2971 29878 3023
rect 29930 3011 29936 3023
rect 31219 3014 31277 3020
rect 31219 3011 31231 3014
rect 29930 2983 31231 3011
rect 29930 2971 29936 2983
rect 31219 2980 31231 2983
rect 31265 2980 31277 3014
rect 31219 2974 31277 2980
rect 31987 3014 32045 3020
rect 31987 2980 31999 3014
rect 32033 2980 32045 3014
rect 31987 2974 32045 2980
rect 27626 2909 29342 2937
rect 27626 2897 27632 2909
rect 30544 2897 30550 2949
rect 30602 2937 30608 2949
rect 32002 2937 32030 2974
rect 32080 2971 32086 3023
rect 32138 3011 32144 3023
rect 33907 3014 33965 3020
rect 33907 3011 33919 3014
rect 32138 2983 33919 3011
rect 32138 2971 32144 2983
rect 33907 2980 33919 2983
rect 33953 2980 33965 3014
rect 33907 2974 33965 2980
rect 34675 3014 34733 3020
rect 34675 2980 34687 3014
rect 34721 2980 34733 3014
rect 34675 2974 34733 2980
rect 30602 2909 32030 2937
rect 30602 2897 30608 2909
rect 32272 2897 32278 2949
rect 32330 2937 32336 2949
rect 33136 2937 33142 2949
rect 32330 2909 33142 2937
rect 32330 2897 32336 2909
rect 33136 2897 33142 2909
rect 33194 2897 33200 2949
rect 33328 2897 33334 2949
rect 33386 2937 33392 2949
rect 34690 2937 34718 2974
rect 35440 2971 35446 3023
rect 35498 3011 35504 3023
rect 36595 3014 36653 3020
rect 36595 3011 36607 3014
rect 35498 2983 36607 3011
rect 35498 2971 35504 2983
rect 36595 2980 36607 2983
rect 36641 2980 36653 3014
rect 36595 2974 36653 2980
rect 37363 3014 37421 3020
rect 37363 2980 37375 3014
rect 37409 2980 37421 3014
rect 37363 2974 37421 2980
rect 33386 2909 34718 2937
rect 33386 2897 33392 2909
rect 36112 2897 36118 2949
rect 36170 2937 36176 2949
rect 37378 2937 37406 2974
rect 37552 2971 37558 3023
rect 37610 3011 37616 3023
rect 39283 3014 39341 3020
rect 39283 3011 39295 3014
rect 37610 2983 39295 3011
rect 37610 2971 37616 2983
rect 39283 2980 39295 2983
rect 39329 2980 39341 3014
rect 39283 2974 39341 2980
rect 40051 3014 40109 3020
rect 40051 2980 40063 3014
rect 40097 2980 40109 3014
rect 40051 2974 40109 2980
rect 36170 2909 37406 2937
rect 36170 2897 36176 2909
rect 38320 2897 38326 2949
rect 38378 2937 38384 2949
rect 40066 2937 40094 2974
rect 40528 2971 40534 3023
rect 40586 3011 40592 3023
rect 41971 3014 42029 3020
rect 41971 3011 41983 3014
rect 40586 2983 41983 3011
rect 40586 2971 40592 2983
rect 41971 2980 41983 2983
rect 42017 2980 42029 3014
rect 41971 2974 42029 2980
rect 42739 3014 42797 3020
rect 42739 2980 42751 3014
rect 42785 2980 42797 3014
rect 42739 2974 42797 2980
rect 38378 2909 40094 2937
rect 38378 2897 38384 2909
rect 41200 2897 41206 2949
rect 41258 2937 41264 2949
rect 42754 2937 42782 2974
rect 43024 2971 43030 3023
rect 43082 3011 43088 3023
rect 44659 3014 44717 3020
rect 44659 3011 44671 3014
rect 43082 2983 44671 3011
rect 43082 2971 43088 2983
rect 44659 2980 44671 2983
rect 44705 2980 44717 3014
rect 44659 2974 44717 2980
rect 45427 3014 45485 3020
rect 45427 2980 45439 3014
rect 45473 2980 45485 3014
rect 45427 2974 45485 2980
rect 41258 2909 42782 2937
rect 41258 2897 41264 2909
rect 44176 2897 44182 2949
rect 44234 2937 44240 2949
rect 45442 2937 45470 2974
rect 45616 2971 45622 3023
rect 45674 3011 45680 3023
rect 48130 3020 48158 3057
rect 51763 3054 51775 3088
rect 51809 3085 51821 3088
rect 52240 3085 52246 3097
rect 51809 3057 52246 3085
rect 51809 3054 51821 3057
rect 51763 3048 51821 3054
rect 52240 3045 52246 3057
rect 52298 3045 52304 3097
rect 56368 3045 56374 3097
rect 56426 3085 56432 3097
rect 56755 3088 56813 3094
rect 56755 3085 56767 3088
rect 56426 3057 56767 3085
rect 56426 3045 56432 3057
rect 56755 3054 56767 3057
rect 56801 3085 56813 3088
rect 56947 3088 57005 3094
rect 56947 3085 56959 3088
rect 56801 3057 56959 3085
rect 56801 3054 56813 3057
rect 56755 3048 56813 3054
rect 56947 3054 56959 3057
rect 56993 3054 57005 3088
rect 56947 3048 57005 3054
rect 47347 3014 47405 3020
rect 47347 3011 47359 3014
rect 45674 2983 47359 3011
rect 45674 2971 45680 2983
rect 47347 2980 47359 2983
rect 47393 2980 47405 3014
rect 47347 2974 47405 2980
rect 48115 3014 48173 3020
rect 48115 2980 48127 3014
rect 48161 2980 48173 3014
rect 48115 2974 48173 2980
rect 49648 2971 49654 3023
rect 49706 3011 49712 3023
rect 50035 3014 50093 3020
rect 50035 3011 50047 3014
rect 49706 2983 50047 3011
rect 49706 2971 49712 2983
rect 50035 2980 50047 2983
rect 50081 2980 50093 3014
rect 50035 2974 50093 2980
rect 50803 3014 50861 3020
rect 50803 2980 50815 3014
rect 50849 2980 50861 3014
rect 50803 2974 50861 2980
rect 50818 2937 50846 2974
rect 51472 2971 51478 3023
rect 51530 3011 51536 3023
rect 52723 3014 52781 3020
rect 52723 3011 52735 3014
rect 51530 2983 52735 3011
rect 51530 2971 51536 2983
rect 52723 2980 52735 2983
rect 52769 2980 52781 3014
rect 53491 3014 53549 3020
rect 53491 3011 53503 3014
rect 52723 2974 52781 2980
rect 52834 2983 53503 3011
rect 44234 2909 45470 2937
rect 50050 2909 50846 2937
rect 44234 2897 44240 2909
rect 50050 2875 50078 2909
rect 52240 2897 52246 2949
rect 52298 2937 52304 2949
rect 52834 2937 52862 2983
rect 53491 2980 53503 2983
rect 53537 2980 53549 3014
rect 53491 2974 53549 2980
rect 53776 2971 53782 3023
rect 53834 3011 53840 3023
rect 55411 3014 55469 3020
rect 55411 3011 55423 3014
rect 53834 2983 55423 3011
rect 53834 2971 53840 2983
rect 55411 2980 55423 2983
rect 55457 2980 55469 3014
rect 55411 2974 55469 2980
rect 56179 3014 56237 3020
rect 56179 2980 56191 3014
rect 56225 2980 56237 3014
rect 56179 2974 56237 2980
rect 52298 2909 52862 2937
rect 52298 2897 52304 2909
rect 52912 2897 52918 2949
rect 52970 2937 52976 2949
rect 53680 2937 53686 2949
rect 52970 2909 53686 2937
rect 52970 2897 52976 2909
rect 53680 2897 53686 2909
rect 53738 2897 53744 2949
rect 54832 2897 54838 2949
rect 54890 2937 54896 2949
rect 56194 2937 56222 2974
rect 56656 2971 56662 3023
rect 56714 3011 56720 3023
rect 57328 3011 57334 3023
rect 56714 2983 57334 3011
rect 56714 2971 56720 2983
rect 57328 2971 57334 2983
rect 57386 2971 57392 3023
rect 54890 2909 56222 2937
rect 54890 2897 54896 2909
rect 6160 2823 6166 2875
rect 6218 2863 6224 2875
rect 46387 2866 46445 2872
rect 46387 2863 46399 2866
rect 6218 2835 13310 2863
rect 6218 2823 6224 2835
rect 5162 2761 5246 2789
rect 13282 2789 13310 2835
rect 17266 2835 33134 2863
rect 17266 2789 17294 2835
rect 13282 2761 17294 2789
rect 5162 2749 5168 2761
rect 19504 2749 19510 2801
rect 19562 2789 19568 2801
rect 20080 2789 20086 2801
rect 19562 2761 20086 2789
rect 19562 2749 19568 2761
rect 20080 2749 20086 2761
rect 20138 2749 20144 2801
rect 22195 2792 22253 2798
rect 22195 2758 22207 2792
rect 22241 2789 22253 2792
rect 23920 2789 23926 2801
rect 22241 2761 23926 2789
rect 22241 2758 22253 2761
rect 22195 2752 22253 2758
rect 23920 2749 23926 2761
rect 23978 2749 23984 2801
rect 27760 2749 27766 2801
rect 27818 2789 27824 2801
rect 27952 2789 27958 2801
rect 27818 2761 27958 2789
rect 27818 2749 27824 2761
rect 27952 2749 27958 2761
rect 28010 2749 28016 2801
rect 33106 2789 33134 2835
rect 43234 2835 46399 2863
rect 43234 2789 43262 2835
rect 46387 2832 46399 2835
rect 46433 2832 46445 2866
rect 46387 2826 46445 2832
rect 50032 2823 50038 2875
rect 50090 2823 50096 2875
rect 33106 2761 43262 2789
rect 43699 2792 43757 2798
rect 43699 2758 43711 2792
rect 43745 2789 43757 2792
rect 45328 2789 45334 2801
rect 43745 2761 45334 2789
rect 43745 2758 43757 2761
rect 43699 2752 43757 2758
rect 45328 2749 45334 2761
rect 45386 2749 45392 2801
rect 46096 2749 46102 2801
rect 46154 2789 46160 2801
rect 47056 2789 47062 2801
rect 46154 2761 47062 2789
rect 46154 2749 46160 2761
rect 47056 2749 47062 2761
rect 47114 2749 47120 2801
rect 48499 2792 48557 2798
rect 48499 2758 48511 2792
rect 48545 2789 48557 2792
rect 54451 2792 54509 2798
rect 54451 2789 54463 2792
rect 48545 2761 54463 2789
rect 48545 2758 48557 2761
rect 48499 2752 48557 2758
rect 54451 2758 54463 2761
rect 54497 2758 54509 2792
rect 54451 2752 54509 2758
rect 1152 2690 58848 2712
rect 1152 2638 4294 2690
rect 4346 2638 4358 2690
rect 4410 2638 4422 2690
rect 4474 2638 4486 2690
rect 4538 2638 35014 2690
rect 35066 2638 35078 2690
rect 35130 2638 35142 2690
rect 35194 2638 35206 2690
rect 35258 2638 58848 2690
rect 1152 2616 58848 2638
rect 3952 2527 3958 2579
rect 4010 2567 4016 2579
rect 4240 2567 4246 2579
rect 4010 2539 4246 2567
rect 4010 2527 4016 2539
rect 4240 2527 4246 2539
rect 4298 2527 4304 2579
rect 4336 2527 4342 2579
rect 4394 2567 4400 2579
rect 4816 2567 4822 2579
rect 4394 2539 4822 2567
rect 4394 2527 4400 2539
rect 4816 2527 4822 2539
rect 4874 2527 4880 2579
rect 9808 2527 9814 2579
rect 9866 2567 9872 2579
rect 10192 2567 10198 2579
rect 9866 2539 10198 2567
rect 9866 2527 9872 2539
rect 10192 2527 10198 2539
rect 10250 2527 10256 2579
rect 13072 2527 13078 2579
rect 13130 2567 13136 2579
rect 13264 2567 13270 2579
rect 13130 2539 13270 2567
rect 13130 2527 13136 2539
rect 13264 2527 13270 2539
rect 13322 2527 13328 2579
rect 20176 2527 20182 2579
rect 20234 2567 20240 2579
rect 20848 2567 20854 2579
rect 20234 2539 20854 2567
rect 20234 2527 20240 2539
rect 20848 2527 20854 2539
rect 20906 2527 20912 2579
rect 43216 2527 43222 2579
rect 43274 2567 43280 2579
rect 43984 2567 43990 2579
rect 43274 2539 43990 2567
rect 43274 2527 43280 2539
rect 43984 2527 43990 2539
rect 44042 2527 44048 2579
rect 45136 2527 45142 2579
rect 45194 2567 45200 2579
rect 45712 2567 45718 2579
rect 45194 2539 45718 2567
rect 45194 2527 45200 2539
rect 45712 2527 45718 2539
rect 45770 2527 45776 2579
rect 4720 2009 4726 2061
rect 4778 2049 4784 2061
rect 5296 2049 5302 2061
rect 4778 2021 5302 2049
rect 4778 2009 4784 2021
rect 5296 2009 5302 2021
rect 5354 2009 5360 2061
rect 4528 1861 4534 1913
rect 4586 1901 4592 1913
rect 4816 1901 4822 1913
rect 4586 1873 4822 1901
rect 4586 1861 4592 1873
rect 4816 1861 4822 1873
rect 4874 1861 4880 1913
rect 30352 1713 30358 1765
rect 30410 1753 30416 1765
rect 30640 1753 30646 1765
rect 30410 1725 30646 1753
rect 30410 1713 30416 1725
rect 30640 1713 30646 1725
rect 30698 1713 30704 1765
rect 50512 1713 50518 1765
rect 50570 1753 50576 1765
rect 51088 1753 51094 1765
rect 50570 1725 51094 1753
rect 50570 1713 50576 1725
rect 51088 1713 51094 1725
rect 51146 1713 51152 1765
rect 36112 1639 36118 1691
rect 36170 1639 36176 1691
rect 50704 1639 50710 1691
rect 50762 1679 50768 1691
rect 50896 1679 50902 1691
rect 50762 1651 50902 1679
rect 50762 1639 50768 1651
rect 50896 1639 50902 1651
rect 50954 1639 50960 1691
rect 35152 1417 35158 1469
rect 35210 1457 35216 1469
rect 35536 1457 35542 1469
rect 35210 1429 35542 1457
rect 35210 1417 35216 1429
rect 35536 1417 35542 1429
rect 35594 1417 35600 1469
rect 36130 1321 36158 1639
rect 36304 1491 36310 1543
rect 36362 1491 36368 1543
rect 50896 1491 50902 1543
rect 50954 1531 50960 1543
rect 51568 1531 51574 1543
rect 50954 1503 51574 1531
rect 50954 1491 50960 1503
rect 51568 1491 51574 1503
rect 51626 1491 51632 1543
rect 33232 1269 33238 1321
rect 33290 1309 33296 1321
rect 33712 1309 33718 1321
rect 33290 1281 33718 1309
rect 33290 1269 33296 1281
rect 33712 1269 33718 1281
rect 33770 1269 33776 1321
rect 36112 1269 36118 1321
rect 36170 1269 36176 1321
rect 36322 1173 36350 1491
rect 41008 1269 41014 1321
rect 41066 1309 41072 1321
rect 41296 1309 41302 1321
rect 41066 1281 41302 1309
rect 41066 1269 41072 1281
rect 41296 1269 41302 1281
rect 41354 1269 41360 1321
rect 34672 1121 34678 1173
rect 34730 1161 34736 1173
rect 35440 1161 35446 1173
rect 34730 1133 35446 1161
rect 34730 1121 34736 1133
rect 35440 1121 35446 1133
rect 35498 1121 35504 1173
rect 36304 1121 36310 1173
rect 36362 1121 36368 1173
rect 34864 1047 34870 1099
rect 34922 1087 34928 1099
rect 36880 1087 36886 1099
rect 34922 1059 36886 1087
rect 34922 1047 34928 1059
rect 36880 1047 36886 1059
rect 36938 1047 36944 1099
rect 35248 973 35254 1025
rect 35306 1013 35312 1025
rect 35920 1013 35926 1025
rect 35306 985 35926 1013
rect 35306 973 35312 985
rect 35920 973 35926 985
rect 35978 973 35984 1025
<< via1 >>
rect 43990 57361 44042 57413
rect 54550 57361 54602 57413
rect 4294 57250 4346 57302
rect 4358 57250 4410 57302
rect 4422 57250 4474 57302
rect 4486 57250 4538 57302
rect 35014 57250 35066 57302
rect 35078 57250 35130 57302
rect 35142 57250 35194 57302
rect 35206 57250 35258 57302
rect 16630 57139 16682 57191
rect 1750 56991 1802 57043
rect 214 56917 266 56969
rect 3286 56991 3338 57043
rect 4918 56917 4970 56969
rect 9622 56991 9674 57043
rect 11254 56991 11306 57043
rect 6454 56917 6506 56969
rect 8086 56960 8138 56969
rect 8086 56926 8095 56960
rect 8095 56926 8129 56960
rect 8129 56926 8138 56960
rect 8086 56917 8138 56926
rect 16438 56991 16490 57043
rect 29110 56991 29162 57043
rect 39478 56991 39530 57043
rect 43798 56991 43850 57043
rect 44086 56991 44138 57043
rect 52054 56991 52106 57043
rect 12790 56917 12842 56969
rect 14422 56917 14474 56969
rect 15958 56917 16010 56969
rect 17494 56917 17546 56969
rect 19126 56917 19178 56969
rect 20662 56917 20714 56969
rect 22294 56917 22346 56969
rect 23830 56917 23882 56969
rect 25462 56917 25514 56969
rect 26998 56917 27050 56969
rect 28630 56960 28682 56969
rect 28630 56926 28639 56960
rect 28639 56926 28673 56960
rect 28673 56926 28682 56960
rect 28630 56917 28682 56926
rect 30262 56960 30314 56969
rect 30262 56926 30271 56960
rect 30271 56926 30305 56960
rect 30305 56926 30314 56960
rect 30262 56917 30314 56926
rect 31702 56960 31754 56969
rect 31702 56926 31711 56960
rect 31711 56926 31745 56960
rect 31745 56926 31754 56960
rect 31702 56917 31754 56926
rect 33334 56917 33386 56969
rect 34870 56960 34922 56969
rect 34870 56926 34879 56960
rect 34879 56926 34913 56960
rect 34913 56926 34922 56960
rect 34870 56917 34922 56926
rect 38038 56960 38090 56969
rect 38038 56926 38047 56960
rect 38047 56926 38081 56960
rect 38081 56926 38090 56960
rect 38038 56917 38090 56926
rect 38134 56917 38186 56969
rect 1750 56886 1802 56895
rect 1750 56852 1759 56886
rect 1759 56852 1793 56886
rect 1793 56852 1802 56886
rect 1750 56843 1802 56852
rect 3574 56843 3626 56895
rect 5110 56886 5162 56895
rect 5110 56852 5119 56886
rect 5119 56852 5153 56886
rect 5153 56852 5162 56886
rect 5110 56843 5162 56852
rect 8278 56843 8330 56895
rect 11254 56886 11306 56895
rect 11254 56852 11263 56886
rect 11263 56852 11297 56886
rect 11297 56852 11306 56886
rect 11254 56843 11306 56852
rect 12982 56886 13034 56895
rect 12982 56852 12991 56886
rect 12991 56852 13025 56886
rect 13025 56852 13034 56886
rect 12982 56843 13034 56852
rect 15574 56843 15626 56895
rect 16150 56886 16202 56895
rect 16150 56852 16159 56886
rect 16159 56852 16193 56886
rect 16193 56852 16202 56886
rect 16150 56843 16202 56852
rect 17974 56886 18026 56895
rect 17974 56852 17983 56886
rect 17983 56852 18017 56886
rect 18017 56852 18026 56886
rect 17974 56843 18026 56852
rect 19318 56886 19370 56895
rect 19318 56852 19327 56886
rect 19327 56852 19361 56886
rect 19361 56852 19370 56886
rect 19318 56843 19370 56852
rect 20854 56886 20906 56895
rect 20854 56852 20863 56886
rect 20863 56852 20897 56886
rect 20897 56852 20906 56886
rect 20854 56843 20906 56852
rect 25174 56843 25226 56895
rect 30070 56886 30122 56895
rect 30070 56852 30079 56886
rect 30079 56852 30113 56886
rect 30113 56852 30122 56886
rect 30070 56843 30122 56852
rect 32662 56886 32714 56895
rect 32662 56852 32671 56886
rect 32671 56852 32705 56886
rect 32705 56852 32714 56886
rect 32662 56843 32714 56852
rect 22294 56769 22346 56821
rect 25558 56769 25610 56821
rect 36502 56843 36554 56895
rect 39670 56843 39722 56895
rect 41206 56917 41258 56969
rect 47542 56960 47594 56969
rect 47542 56926 47551 56960
rect 47551 56926 47585 56960
rect 47585 56926 47594 56960
rect 47542 56917 47594 56926
rect 52246 56917 52298 56969
rect 41206 56769 41258 56821
rect 42838 56843 42890 56895
rect 44374 56843 44426 56895
rect 45910 56843 45962 56895
rect 49078 56843 49130 56895
rect 50710 56843 50762 56895
rect 53878 56843 53930 56895
rect 55414 56843 55466 56895
rect 57046 56886 57098 56895
rect 57046 56852 57055 56886
rect 57055 56852 57089 56886
rect 57089 56852 57098 56886
rect 57046 56843 57098 56852
rect 55318 56769 55370 56821
rect 9718 56695 9770 56747
rect 36694 56738 36746 56747
rect 36694 56704 36703 56738
rect 36703 56704 36737 56738
rect 36737 56704 36746 56738
rect 36694 56695 36746 56704
rect 39766 56738 39818 56747
rect 39766 56704 39775 56738
rect 39775 56704 39809 56738
rect 39809 56704 39818 56738
rect 39766 56695 39818 56704
rect 40822 56738 40874 56747
rect 40822 56704 40831 56738
rect 40831 56704 40865 56738
rect 40865 56704 40874 56738
rect 40822 56695 40874 56704
rect 42934 56738 42986 56747
rect 42934 56704 42943 56738
rect 42943 56704 42977 56738
rect 42977 56704 42986 56738
rect 42934 56695 42986 56704
rect 44758 56738 44810 56747
rect 44758 56704 44767 56738
rect 44767 56704 44801 56738
rect 44801 56704 44810 56738
rect 44758 56695 44810 56704
rect 46102 56695 46154 56747
rect 48694 56738 48746 56747
rect 48694 56704 48703 56738
rect 48703 56704 48737 56738
rect 48737 56704 48746 56738
rect 48694 56695 48746 56704
rect 50806 56738 50858 56747
rect 50806 56704 50815 56738
rect 50815 56704 50849 56738
rect 50849 56704 50858 56738
rect 50806 56695 50858 56704
rect 53974 56738 54026 56747
rect 53974 56704 53983 56738
rect 53983 56704 54017 56738
rect 54017 56704 54026 56738
rect 53974 56695 54026 56704
rect 55510 56738 55562 56747
rect 55510 56704 55519 56738
rect 55519 56704 55553 56738
rect 55553 56704 55562 56738
rect 55510 56695 55562 56704
rect 19654 56584 19706 56636
rect 19718 56584 19770 56636
rect 19782 56584 19834 56636
rect 19846 56584 19898 56636
rect 50374 56584 50426 56636
rect 50438 56584 50490 56636
rect 50502 56584 50554 56636
rect 50566 56584 50618 56636
rect 694 56473 746 56525
rect 2230 56473 2282 56525
rect 2806 56473 2858 56525
rect 3862 56473 3914 56525
rect 5398 56473 5450 56525
rect 5974 56473 6026 56525
rect 7030 56473 7082 56525
rect 8566 56473 8618 56525
rect 10198 56473 10250 56525
rect 10678 56473 10730 56525
rect 11734 56473 11786 56525
rect 12310 56473 12362 56525
rect 13366 56473 13418 56525
rect 14902 56473 14954 56525
rect 17014 56473 17066 56525
rect 18070 56473 18122 56525
rect 18550 56473 18602 56525
rect 19990 56473 20042 56525
rect 21238 56473 21290 56525
rect 21718 56473 21770 56525
rect 22774 56473 22826 56525
rect 24406 56516 24458 56525
rect 24406 56482 24415 56516
rect 24415 56482 24449 56516
rect 24449 56482 24458 56516
rect 24406 56473 24458 56482
rect 25942 56473 25994 56525
rect 26518 56473 26570 56525
rect 27574 56473 27626 56525
rect 28054 56473 28106 56525
rect 29686 56516 29738 56525
rect 29686 56482 29695 56516
rect 29695 56482 29729 56516
rect 29729 56482 29738 56516
rect 29686 56473 29738 56482
rect 30646 56473 30698 56525
rect 31222 56473 31274 56525
rect 32278 56473 32330 56525
rect 33814 56473 33866 56525
rect 34582 56473 34634 56525
rect 35446 56473 35498 56525
rect 36214 56473 36266 56525
rect 37558 56473 37610 56525
rect 38614 56473 38666 56525
rect 40150 56516 40202 56525
rect 40150 56482 40159 56516
rect 40159 56482 40193 56516
rect 40193 56482 40202 56516
rect 40150 56473 40202 56482
rect 41782 56473 41834 56525
rect 42262 56473 42314 56525
rect 43318 56473 43370 56525
rect 43894 56473 43946 56525
rect 44950 56473 45002 56525
rect 46486 56473 46538 56525
rect 48022 56473 48074 56525
rect 49654 56473 49706 56525
rect 50134 56473 50186 56525
rect 51286 56473 51338 56525
rect 52822 56473 52874 56525
rect 53302 56473 53354 56525
rect 54358 56473 54410 56525
rect 54934 56473 54986 56525
rect 55990 56473 56042 56525
rect 16534 56399 16586 56451
rect 48694 56399 48746 56451
rect 55126 56399 55178 56451
rect 15286 56325 15338 56377
rect 39478 56325 39530 56377
rect 39574 56325 39626 56377
rect 42454 56325 42506 56377
rect 43894 56325 43946 56377
rect 55510 56325 55562 56377
rect 6742 56251 6794 56303
rect 30262 56251 30314 56303
rect 41302 56251 41354 56303
rect 52054 56294 52106 56303
rect 52054 56260 52063 56294
rect 52063 56260 52097 56294
rect 52097 56260 52106 56294
rect 52054 56251 52106 56260
rect 54550 56294 54602 56303
rect 1942 56220 1994 56229
rect 1942 56186 1951 56220
rect 1951 56186 1985 56220
rect 1985 56186 1994 56220
rect 1942 56177 1994 56186
rect 2518 56220 2570 56229
rect 2518 56186 2527 56220
rect 2527 56186 2561 56220
rect 2561 56186 2570 56220
rect 2518 56177 2570 56186
rect 2902 56220 2954 56229
rect 2902 56186 2911 56220
rect 2911 56186 2945 56220
rect 2945 56186 2954 56220
rect 2902 56177 2954 56186
rect 4726 56177 4778 56229
rect 5206 56220 5258 56229
rect 5206 56186 5215 56220
rect 5215 56186 5249 56220
rect 5249 56186 5258 56220
rect 5206 56177 5258 56186
rect 6358 56220 6410 56229
rect 6358 56186 6367 56220
rect 6367 56186 6401 56220
rect 6401 56186 6410 56220
rect 6358 56177 6410 56186
rect 7222 56220 7274 56229
rect 7222 56186 7231 56220
rect 7231 56186 7265 56220
rect 7265 56186 7274 56220
rect 7222 56177 7274 56186
rect 8566 56220 8618 56229
rect 8566 56186 8575 56220
rect 8575 56186 8609 56220
rect 8609 56186 8618 56220
rect 8566 56177 8618 56186
rect 10582 56177 10634 56229
rect 11158 56220 11210 56229
rect 11158 56186 11167 56220
rect 11167 56186 11201 56220
rect 11201 56186 11210 56220
rect 11158 56177 11210 56186
rect 11542 56220 11594 56229
rect 11542 56186 11551 56220
rect 11551 56186 11585 56220
rect 11585 56186 11594 56220
rect 11542 56177 11594 56186
rect 12694 56220 12746 56229
rect 12694 56186 12703 56220
rect 12703 56186 12737 56220
rect 12737 56186 12746 56220
rect 12694 56177 12746 56186
rect 13558 56220 13610 56229
rect 13558 56186 13567 56220
rect 13567 56186 13601 56220
rect 13601 56186 13610 56220
rect 14710 56220 14762 56229
rect 13558 56177 13610 56186
rect 14710 56186 14719 56220
rect 14719 56186 14753 56220
rect 14753 56186 14762 56220
rect 14710 56177 14762 56186
rect 15478 56220 15530 56229
rect 15478 56186 15487 56220
rect 15487 56186 15521 56220
rect 15521 56186 15530 56220
rect 15478 56177 15530 56186
rect 15382 56103 15434 56155
rect 15958 56177 16010 56229
rect 18262 56220 18314 56229
rect 18262 56186 18271 56220
rect 18271 56186 18305 56220
rect 18305 56186 18314 56220
rect 18262 56177 18314 56186
rect 19030 56220 19082 56229
rect 19030 56186 19039 56220
rect 19039 56186 19073 56220
rect 19073 56186 19082 56220
rect 19030 56177 19082 56186
rect 20566 56177 20618 56229
rect 21046 56220 21098 56229
rect 21046 56186 21055 56220
rect 21055 56186 21089 56220
rect 21089 56186 21098 56220
rect 21046 56177 21098 56186
rect 22870 56220 22922 56229
rect 22870 56186 22879 56220
rect 22879 56186 22913 56220
rect 22913 56186 22922 56220
rect 22870 56177 22922 56186
rect 24310 56220 24362 56229
rect 24310 56186 24319 56220
rect 24319 56186 24353 56220
rect 24353 56186 24362 56220
rect 24310 56177 24362 56186
rect 26518 56220 26570 56229
rect 26518 56186 26527 56220
rect 26527 56186 26561 56220
rect 26561 56186 26570 56220
rect 26518 56177 26570 56186
rect 27670 56220 27722 56229
rect 27670 56186 27679 56220
rect 27679 56186 27713 56220
rect 27713 56186 27722 56220
rect 27670 56177 27722 56186
rect 28150 56220 28202 56229
rect 28150 56186 28159 56220
rect 28159 56186 28193 56220
rect 28193 56186 28202 56220
rect 28150 56177 28202 56186
rect 29302 56220 29354 56229
rect 29302 56186 29311 56220
rect 29311 56186 29345 56220
rect 29345 56186 29354 56220
rect 29302 56177 29354 56186
rect 30934 56220 30986 56229
rect 30934 56186 30943 56220
rect 30943 56186 30977 56220
rect 30977 56186 30986 56220
rect 30934 56177 30986 56186
rect 32470 56220 32522 56229
rect 32470 56186 32479 56220
rect 32479 56186 32513 56220
rect 32513 56186 32522 56220
rect 32470 56177 32522 56186
rect 33046 56177 33098 56229
rect 34390 56220 34442 56229
rect 32758 56103 32810 56155
rect 34390 56186 34399 56220
rect 34399 56186 34433 56220
rect 34433 56186 34442 56220
rect 34390 56177 34442 56186
rect 36214 56220 36266 56229
rect 36214 56186 36223 56220
rect 36223 56186 36257 56220
rect 36257 56186 36266 56220
rect 36214 56177 36266 56186
rect 36598 56220 36650 56229
rect 36598 56186 36607 56220
rect 36607 56186 36641 56220
rect 36641 56186 36650 56220
rect 36598 56177 36650 56186
rect 37654 56220 37706 56229
rect 37654 56186 37663 56220
rect 37663 56186 37697 56220
rect 37697 56186 37706 56220
rect 37654 56177 37706 56186
rect 38614 56177 38666 56229
rect 39862 56220 39914 56229
rect 39862 56186 39871 56220
rect 39871 56186 39905 56220
rect 39905 56186 39914 56220
rect 39862 56177 39914 56186
rect 41110 56177 41162 56229
rect 37078 56103 37130 56155
rect 40822 56103 40874 56155
rect 42646 56220 42698 56229
rect 42646 56186 42655 56220
rect 42655 56186 42689 56220
rect 42689 56186 42698 56220
rect 42646 56177 42698 56186
rect 44374 56177 44426 56229
rect 46870 56177 46922 56229
rect 48886 56220 48938 56229
rect 48886 56186 48895 56220
rect 48895 56186 48929 56220
rect 48929 56186 48938 56220
rect 48886 56177 48938 56186
rect 52630 56220 52682 56229
rect 48598 56103 48650 56155
rect 52630 56186 52639 56220
rect 52639 56186 52673 56220
rect 52673 56186 52682 56220
rect 52630 56177 52682 56186
rect 53686 56220 53738 56229
rect 53686 56186 53695 56220
rect 53695 56186 53729 56220
rect 53729 56186 53738 56220
rect 53686 56177 53738 56186
rect 54550 56260 54559 56294
rect 54559 56260 54593 56294
rect 54593 56260 54602 56294
rect 54550 56251 54602 56260
rect 55030 56251 55082 56303
rect 58582 56251 58634 56303
rect 55318 56220 55370 56229
rect 55318 56186 55327 56220
rect 55327 56186 55361 56220
rect 55361 56186 55370 56220
rect 55318 56177 55370 56186
rect 56950 56177 57002 56229
rect 4294 55918 4346 55970
rect 4358 55918 4410 55970
rect 4422 55918 4474 55970
rect 4486 55918 4538 55970
rect 35014 55918 35066 55970
rect 35078 55918 35130 55970
rect 35142 55918 35194 55970
rect 35206 55918 35258 55970
rect 1174 55659 1226 55711
rect 4630 55659 4682 55711
rect 7510 55659 7562 55711
rect 9142 55659 9194 55711
rect 13846 55659 13898 55711
rect 20182 55659 20234 55711
rect 23350 55659 23402 55711
rect 24886 55659 24938 55711
rect 39094 55659 39146 55711
rect 40726 55659 40778 55711
rect 45430 55659 45482 55711
rect 46966 55659 47018 55711
rect 51766 55659 51818 55711
rect 56470 55659 56522 55711
rect 57526 55659 57578 55711
rect 38806 55585 38858 55637
rect 1846 55511 1898 55563
rect 4630 55511 4682 55563
rect 7702 55554 7754 55563
rect 7702 55520 7711 55554
rect 7711 55520 7745 55554
rect 7745 55520 7754 55554
rect 7702 55511 7754 55520
rect 20374 55554 20426 55563
rect 20374 55520 20383 55554
rect 20383 55520 20417 55554
rect 20417 55520 20426 55554
rect 20374 55511 20426 55520
rect 23446 55554 23498 55563
rect 23446 55520 23455 55554
rect 23455 55520 23489 55554
rect 23489 55520 23498 55554
rect 23446 55511 23498 55520
rect 25078 55554 25130 55563
rect 25078 55520 25087 55554
rect 25087 55520 25121 55554
rect 25121 55520 25130 55554
rect 25078 55511 25130 55520
rect 28246 55554 28298 55563
rect 28246 55520 28255 55554
rect 28255 55520 28289 55554
rect 28289 55520 28298 55554
rect 28246 55511 28298 55520
rect 40822 55554 40874 55563
rect 40822 55520 40831 55554
rect 40831 55520 40865 55554
rect 40865 55520 40874 55554
rect 40822 55511 40874 55520
rect 8950 55406 9002 55415
rect 8950 55372 8959 55406
rect 8959 55372 8993 55406
rect 8993 55372 9002 55406
rect 8950 55363 9002 55372
rect 13654 55406 13706 55415
rect 13654 55372 13663 55406
rect 13663 55372 13697 55406
rect 13697 55372 13706 55406
rect 13654 55363 13706 55372
rect 29014 55363 29066 55415
rect 38902 55406 38954 55415
rect 38902 55372 38911 55406
rect 38911 55372 38945 55406
rect 38945 55372 38954 55406
rect 38902 55363 38954 55372
rect 45142 55363 45194 55415
rect 47158 55554 47210 55563
rect 47158 55520 47167 55554
rect 47167 55520 47201 55554
rect 47201 55520 47210 55554
rect 47158 55511 47210 55520
rect 56566 55554 56618 55563
rect 56566 55520 56575 55554
rect 56575 55520 56609 55554
rect 56609 55520 56618 55554
rect 56566 55511 56618 55520
rect 57430 55554 57482 55563
rect 57430 55520 57439 55554
rect 57439 55520 57473 55554
rect 57473 55520 57482 55554
rect 57430 55511 57482 55520
rect 49174 55363 49226 55415
rect 19654 55252 19706 55304
rect 19718 55252 19770 55304
rect 19782 55252 19834 55304
rect 19846 55252 19898 55304
rect 50374 55252 50426 55304
rect 50438 55252 50490 55304
rect 50502 55252 50554 55304
rect 50566 55252 50618 55304
rect 59158 55141 59210 55193
rect 35350 55067 35402 55119
rect 47158 55067 47210 55119
rect 28246 54993 28298 55045
rect 55606 54993 55658 55045
rect 25270 54740 25322 54749
rect 25270 54706 25279 54740
rect 25279 54706 25313 54740
rect 25313 54706 25322 54740
rect 25270 54697 25322 54706
rect 50230 54771 50282 54823
rect 4294 54586 4346 54638
rect 4358 54586 4410 54638
rect 4422 54586 4474 54638
rect 4486 54586 4538 54638
rect 35014 54586 35066 54638
rect 35078 54586 35130 54638
rect 35142 54586 35194 54638
rect 35206 54586 35258 54638
rect 58102 54327 58154 54379
rect 57814 54222 57866 54231
rect 56374 54074 56426 54083
rect 56374 54040 56383 54074
rect 56383 54040 56417 54074
rect 56417 54040 56426 54074
rect 57814 54188 57823 54222
rect 57823 54188 57857 54222
rect 57857 54188 57866 54222
rect 57814 54179 57866 54188
rect 56374 54031 56426 54040
rect 19654 53920 19706 53972
rect 19718 53920 19770 53972
rect 19782 53920 19834 53972
rect 19846 53920 19898 53972
rect 50374 53920 50426 53972
rect 50438 53920 50490 53972
rect 50502 53920 50554 53972
rect 50566 53920 50618 53972
rect 59638 53809 59690 53861
rect 3670 53513 3722 53565
rect 44470 53439 44522 53491
rect 2230 53408 2282 53417
rect 2230 53374 2239 53408
rect 2239 53374 2273 53408
rect 2273 53374 2282 53408
rect 2230 53365 2282 53374
rect 17590 53408 17642 53417
rect 17590 53374 17599 53408
rect 17599 53374 17633 53408
rect 17633 53374 17642 53408
rect 17590 53365 17642 53374
rect 39382 53408 39434 53417
rect 39382 53374 39391 53408
rect 39391 53374 39425 53408
rect 39425 53374 39434 53408
rect 39382 53365 39434 53374
rect 43126 53408 43178 53417
rect 43126 53374 43135 53408
rect 43135 53374 43169 53408
rect 43169 53374 43178 53408
rect 43126 53365 43178 53374
rect 57718 53365 57770 53417
rect 4294 53254 4346 53306
rect 4358 53254 4410 53306
rect 4422 53254 4474 53306
rect 4486 53254 4538 53306
rect 35014 53254 35066 53306
rect 35078 53254 35130 53306
rect 35142 53254 35194 53306
rect 35206 53254 35258 53306
rect 15574 52995 15626 53047
rect 51670 52847 51722 52899
rect 19654 52588 19706 52640
rect 19718 52588 19770 52640
rect 19782 52588 19834 52640
rect 19846 52588 19898 52640
rect 50374 52588 50426 52640
rect 50438 52588 50490 52640
rect 50502 52588 50554 52640
rect 50566 52588 50618 52640
rect 38134 52329 38186 52381
rect 31318 52107 31370 52159
rect 18358 52076 18410 52085
rect 18358 52042 18367 52076
rect 18367 52042 18401 52076
rect 18401 52042 18410 52076
rect 18358 52033 18410 52042
rect 40054 52076 40106 52085
rect 40054 52042 40063 52076
rect 40063 52042 40097 52076
rect 40097 52042 40106 52076
rect 40054 52033 40106 52042
rect 4294 51922 4346 51974
rect 4358 51922 4410 51974
rect 4422 51922 4474 51974
rect 4486 51922 4538 51974
rect 35014 51922 35066 51974
rect 35078 51922 35130 51974
rect 35142 51922 35194 51974
rect 35206 51922 35258 51974
rect 30262 51663 30314 51715
rect 44086 51441 44138 51493
rect 19654 51256 19706 51308
rect 19718 51256 19770 51308
rect 19782 51256 19834 51308
rect 19846 51256 19898 51308
rect 50374 51256 50426 51308
rect 50438 51256 50490 51308
rect 50502 51256 50554 51308
rect 50566 51256 50618 51308
rect 45238 50701 45290 50753
rect 53590 50744 53642 50753
rect 53590 50710 53599 50744
rect 53599 50710 53633 50744
rect 53633 50710 53642 50744
rect 53590 50701 53642 50710
rect 4294 50590 4346 50642
rect 4358 50590 4410 50642
rect 4422 50590 4474 50642
rect 4486 50590 4538 50642
rect 35014 50590 35066 50642
rect 35078 50590 35130 50642
rect 35142 50590 35194 50642
rect 35206 50590 35258 50642
rect 39478 50226 39530 50235
rect 39478 50192 39487 50226
rect 39487 50192 39521 50226
rect 39521 50192 39530 50226
rect 39478 50183 39530 50192
rect 18262 50035 18314 50087
rect 39478 50035 39530 50087
rect 57622 50035 57674 50087
rect 19654 49924 19706 49976
rect 19718 49924 19770 49976
rect 19782 49924 19834 49976
rect 19846 49924 19898 49976
rect 50374 49924 50426 49976
rect 50438 49924 50490 49976
rect 50502 49924 50554 49976
rect 50566 49924 50618 49976
rect 28822 49813 28874 49865
rect 57622 49813 57674 49865
rect 11926 49412 11978 49421
rect 11926 49378 11935 49412
rect 11935 49378 11969 49412
rect 11969 49378 11978 49412
rect 11926 49369 11978 49378
rect 15670 49412 15722 49421
rect 15670 49378 15679 49412
rect 15679 49378 15713 49412
rect 15713 49378 15722 49412
rect 15670 49369 15722 49378
rect 52438 49412 52490 49421
rect 52438 49378 52447 49412
rect 52447 49378 52481 49412
rect 52481 49378 52490 49412
rect 52438 49369 52490 49378
rect 4294 49258 4346 49310
rect 4358 49258 4410 49310
rect 4422 49258 4474 49310
rect 4486 49258 4538 49310
rect 35014 49258 35066 49310
rect 35078 49258 35130 49310
rect 35142 49258 35194 49310
rect 35206 49258 35258 49310
rect 32662 48999 32714 49051
rect 32086 48925 32138 48977
rect 51766 48851 51818 48903
rect 44374 48703 44426 48755
rect 19654 48592 19706 48644
rect 19718 48592 19770 48644
rect 19782 48592 19834 48644
rect 19846 48592 19898 48644
rect 50374 48592 50426 48644
rect 50438 48592 50490 48644
rect 50502 48592 50554 48644
rect 50566 48592 50618 48644
rect 41302 48524 41354 48533
rect 41302 48490 41311 48524
rect 41311 48490 41345 48524
rect 41345 48490 41354 48524
rect 41302 48481 41354 48490
rect 3766 48037 3818 48089
rect 52246 48037 52298 48089
rect 4294 47926 4346 47978
rect 4358 47926 4410 47978
rect 4422 47926 4474 47978
rect 4486 47926 4538 47978
rect 35014 47926 35066 47978
rect 35078 47926 35130 47978
rect 35142 47926 35194 47978
rect 35206 47926 35258 47978
rect 34582 47562 34634 47571
rect 34582 47528 34591 47562
rect 34591 47528 34625 47562
rect 34625 47528 34634 47562
rect 34582 47519 34634 47528
rect 19654 47260 19706 47312
rect 19718 47260 19770 47312
rect 19782 47260 19834 47312
rect 19846 47260 19898 47312
rect 50374 47260 50426 47312
rect 50438 47260 50490 47312
rect 50502 47260 50554 47312
rect 50566 47260 50618 47312
rect 6742 47044 6794 47053
rect 6742 47010 6751 47044
rect 6751 47010 6785 47044
rect 6785 47010 6794 47044
rect 6742 47001 6794 47010
rect 23638 46748 23690 46757
rect 23638 46714 23647 46748
rect 23647 46714 23681 46748
rect 23681 46714 23690 46748
rect 23638 46705 23690 46714
rect 4294 46594 4346 46646
rect 4358 46594 4410 46646
rect 4422 46594 4474 46646
rect 4486 46594 4538 46646
rect 35014 46594 35066 46646
rect 35078 46594 35130 46646
rect 35142 46594 35194 46646
rect 35206 46594 35258 46646
rect 9910 46230 9962 46239
rect 9910 46196 9919 46230
rect 9919 46196 9953 46230
rect 9953 46196 9962 46230
rect 9910 46187 9962 46196
rect 2518 46039 2570 46091
rect 19654 45928 19706 45980
rect 19718 45928 19770 45980
rect 19782 45928 19834 45980
rect 19846 45928 19898 45980
rect 50374 45928 50426 45980
rect 50438 45928 50490 45980
rect 50502 45928 50554 45980
rect 50566 45928 50618 45980
rect 35350 45669 35402 45721
rect 51574 45373 51626 45425
rect 4294 45262 4346 45314
rect 4358 45262 4410 45314
rect 4422 45262 4474 45314
rect 4486 45262 4538 45314
rect 35014 45262 35066 45314
rect 35078 45262 35130 45314
rect 35142 45262 35194 45314
rect 35206 45262 35258 45314
rect 19990 45151 20042 45203
rect 38806 45194 38858 45203
rect 38806 45160 38815 45194
rect 38815 45160 38849 45194
rect 38849 45160 38858 45194
rect 38806 45151 38858 45160
rect 51574 45077 51626 45129
rect 42454 45003 42506 45055
rect 11158 44929 11210 44981
rect 8470 44898 8522 44907
rect 8470 44864 8479 44898
rect 8479 44864 8513 44898
rect 8513 44864 8522 44898
rect 8470 44855 8522 44864
rect 21334 44898 21386 44907
rect 21334 44864 21343 44898
rect 21343 44864 21377 44898
rect 21377 44864 21386 44898
rect 21334 44855 21386 44864
rect 41014 44750 41066 44759
rect 41014 44716 41023 44750
rect 41023 44716 41057 44750
rect 41057 44716 41066 44750
rect 41014 44707 41066 44716
rect 19654 44596 19706 44648
rect 19718 44596 19770 44648
rect 19782 44596 19834 44648
rect 19846 44596 19898 44648
rect 50374 44596 50426 44648
rect 50438 44596 50490 44648
rect 50502 44596 50554 44648
rect 50566 44596 50618 44648
rect 44374 44041 44426 44093
rect 4294 43930 4346 43982
rect 4358 43930 4410 43982
rect 4422 43930 4474 43982
rect 4486 43930 4538 43982
rect 35014 43930 35066 43982
rect 35078 43930 35130 43982
rect 35142 43930 35194 43982
rect 35206 43930 35258 43982
rect 15766 43523 15818 43575
rect 50038 43375 50090 43427
rect 19654 43264 19706 43316
rect 19718 43264 19770 43316
rect 19782 43264 19834 43316
rect 19846 43264 19898 43316
rect 50374 43264 50426 43316
rect 50438 43264 50490 43316
rect 50502 43264 50554 43316
rect 50566 43264 50618 43316
rect 40822 42709 40874 42761
rect 46390 42752 46442 42761
rect 46390 42718 46399 42752
rect 46399 42718 46433 42752
rect 46433 42718 46442 42752
rect 46390 42709 46442 42718
rect 53878 42709 53930 42761
rect 4294 42598 4346 42650
rect 4358 42598 4410 42650
rect 4422 42598 4474 42650
rect 4486 42598 4538 42650
rect 35014 42598 35066 42650
rect 35078 42598 35130 42650
rect 35142 42598 35194 42650
rect 35206 42598 35258 42650
rect 32662 42487 32714 42539
rect 53878 42487 53930 42539
rect 57334 42043 57386 42095
rect 19654 41932 19706 41984
rect 19718 41932 19770 41984
rect 19782 41932 19834 41984
rect 19846 41932 19898 41984
rect 50374 41932 50426 41984
rect 50438 41932 50490 41984
rect 50502 41932 50554 41984
rect 50566 41932 50618 41984
rect 43990 41747 44042 41799
rect 52342 41377 52394 41429
rect 4294 41266 4346 41318
rect 4358 41266 4410 41318
rect 4422 41266 4474 41318
rect 4486 41266 4538 41318
rect 35014 41266 35066 41318
rect 35078 41266 35130 41318
rect 35142 41266 35194 41318
rect 35206 41266 35258 41318
rect 26134 40859 26186 40911
rect 44566 40933 44618 40985
rect 12214 40711 12266 40763
rect 25366 40711 25418 40763
rect 19654 40600 19706 40652
rect 19718 40600 19770 40652
rect 19782 40600 19834 40652
rect 19846 40600 19898 40652
rect 50374 40600 50426 40652
rect 50438 40600 50490 40652
rect 50502 40600 50554 40652
rect 50566 40600 50618 40652
rect 29110 40045 29162 40097
rect 4294 39934 4346 39986
rect 4358 39934 4410 39986
rect 4422 39934 4474 39986
rect 4486 39934 4538 39986
rect 35014 39934 35066 39986
rect 35078 39934 35130 39986
rect 35142 39934 35194 39986
rect 35206 39934 35258 39986
rect 46870 39823 46922 39875
rect 32470 39527 32522 39579
rect 44086 39570 44138 39579
rect 44086 39536 44095 39570
rect 44095 39536 44129 39570
rect 44129 39536 44138 39570
rect 44086 39527 44138 39536
rect 30646 39453 30698 39505
rect 6742 39422 6794 39431
rect 6742 39388 6751 39422
rect 6751 39388 6785 39422
rect 6785 39388 6794 39422
rect 6742 39379 6794 39388
rect 19654 39268 19706 39320
rect 19718 39268 19770 39320
rect 19782 39268 19834 39320
rect 19846 39268 19898 39320
rect 50374 39268 50426 39320
rect 50438 39268 50490 39320
rect 50502 39268 50554 39320
rect 50566 39268 50618 39320
rect 44086 39157 44138 39209
rect 53206 39157 53258 39209
rect 15286 38830 15338 38839
rect 15286 38796 15295 38830
rect 15295 38796 15329 38830
rect 15329 38796 15338 38830
rect 15286 38787 15338 38796
rect 21910 38713 21962 38765
rect 56470 38713 56522 38765
rect 4294 38602 4346 38654
rect 4358 38602 4410 38654
rect 4422 38602 4474 38654
rect 4486 38602 4538 38654
rect 35014 38602 35066 38654
rect 35078 38602 35130 38654
rect 35142 38602 35194 38654
rect 35206 38602 35258 38654
rect 39574 38491 39626 38543
rect 13558 38269 13610 38321
rect 38614 38269 38666 38321
rect 14230 38090 14282 38099
rect 14230 38056 14239 38090
rect 14239 38056 14273 38090
rect 14273 38056 14282 38090
rect 14230 38047 14282 38056
rect 18070 38090 18122 38099
rect 18070 38056 18079 38090
rect 18079 38056 18113 38090
rect 18113 38056 18122 38090
rect 18070 38047 18122 38056
rect 38326 38047 38378 38099
rect 19654 37936 19706 37988
rect 19718 37936 19770 37988
rect 19782 37936 19834 37988
rect 19846 37936 19898 37988
rect 50374 37936 50426 37988
rect 50438 37936 50490 37988
rect 50502 37936 50554 37988
rect 50566 37936 50618 37988
rect 6838 37825 6890 37877
rect 18070 37825 18122 37877
rect 11350 37381 11402 37433
rect 51286 37381 51338 37433
rect 55894 37381 55946 37433
rect 4294 37270 4346 37322
rect 4358 37270 4410 37322
rect 4422 37270 4474 37322
rect 4486 37270 4538 37322
rect 35014 37270 35066 37322
rect 35078 37270 35130 37322
rect 35142 37270 35194 37322
rect 35206 37270 35258 37322
rect 15094 36863 15146 36915
rect 19654 36604 19706 36656
rect 19718 36604 19770 36656
rect 19782 36604 19834 36656
rect 19846 36604 19898 36656
rect 50374 36604 50426 36656
rect 50438 36604 50490 36656
rect 50502 36604 50554 36656
rect 50566 36604 50618 36656
rect 14998 36092 15050 36101
rect 14998 36058 15007 36092
rect 15007 36058 15041 36092
rect 15041 36058 15050 36092
rect 14998 36049 15050 36058
rect 46198 36049 46250 36101
rect 46294 36049 46346 36101
rect 4294 35938 4346 35990
rect 4358 35938 4410 35990
rect 4422 35938 4474 35990
rect 4486 35938 4538 35990
rect 35014 35938 35066 35990
rect 35078 35938 35130 35990
rect 35142 35938 35194 35990
rect 35206 35938 35258 35990
rect 31030 35679 31082 35731
rect 8566 35605 8618 35657
rect 33526 35574 33578 35583
rect 33526 35540 33535 35574
rect 33535 35540 33569 35574
rect 33569 35540 33578 35574
rect 33526 35531 33578 35540
rect 19654 35272 19706 35324
rect 19718 35272 19770 35324
rect 19782 35272 19834 35324
rect 19846 35272 19898 35324
rect 50374 35272 50426 35324
rect 50438 35272 50490 35324
rect 50502 35272 50554 35324
rect 50566 35272 50618 35324
rect 14806 34760 14858 34769
rect 14806 34726 14815 34760
rect 14815 34726 14849 34760
rect 14849 34726 14858 34760
rect 14806 34717 14858 34726
rect 19030 34717 19082 34769
rect 32758 34760 32810 34769
rect 32758 34726 32767 34760
rect 32767 34726 32801 34760
rect 32801 34726 32810 34760
rect 32758 34717 32810 34726
rect 4294 34606 4346 34658
rect 4358 34606 4410 34658
rect 4422 34606 4474 34658
rect 4486 34606 4538 34658
rect 35014 34606 35066 34658
rect 35078 34606 35130 34658
rect 35142 34606 35194 34658
rect 35206 34606 35258 34658
rect 24022 34199 24074 34251
rect 19654 33940 19706 33992
rect 19718 33940 19770 33992
rect 19782 33940 19834 33992
rect 19846 33940 19898 33992
rect 50374 33940 50426 33992
rect 50438 33940 50490 33992
rect 50502 33940 50554 33992
rect 50566 33940 50618 33992
rect 1846 33607 1898 33659
rect 28246 33607 28298 33659
rect 28342 33459 28394 33511
rect 12694 33385 12746 33437
rect 47734 33385 47786 33437
rect 4294 33274 4346 33326
rect 4358 33274 4410 33326
rect 4422 33274 4474 33326
rect 4486 33274 4538 33326
rect 35014 33274 35066 33326
rect 35078 33274 35130 33326
rect 35142 33274 35194 33326
rect 35206 33274 35258 33326
rect 47734 33206 47786 33215
rect 28246 33132 28298 33141
rect 28246 33098 28255 33132
rect 28255 33098 28289 33132
rect 28289 33098 28298 33132
rect 28246 33089 28298 33098
rect 47734 33172 47743 33206
rect 47743 33172 47777 33206
rect 47777 33172 47786 33206
rect 47734 33163 47786 33172
rect 56566 33163 56618 33215
rect 42358 32910 42410 32919
rect 42358 32876 42367 32910
rect 42367 32876 42401 32910
rect 42401 32876 42410 32910
rect 42358 32867 42410 32876
rect 19654 32608 19706 32660
rect 19718 32608 19770 32660
rect 19782 32608 19834 32660
rect 19846 32608 19898 32660
rect 50374 32608 50426 32660
rect 50438 32608 50490 32660
rect 50502 32608 50554 32660
rect 50566 32608 50618 32660
rect 20566 32497 20618 32549
rect 13942 32096 13994 32105
rect 13942 32062 13951 32096
rect 13951 32062 13985 32096
rect 13985 32062 13994 32096
rect 13942 32053 13994 32062
rect 31222 32053 31274 32105
rect 34774 32053 34826 32105
rect 4294 31942 4346 31994
rect 4358 31942 4410 31994
rect 4422 31942 4474 31994
rect 4486 31942 4538 31994
rect 35014 31942 35066 31994
rect 35078 31942 35130 31994
rect 35142 31942 35194 31994
rect 35206 31942 35258 31994
rect 41110 31831 41162 31883
rect 48310 31683 48362 31735
rect 19654 31276 19706 31328
rect 19718 31276 19770 31328
rect 19782 31276 19834 31328
rect 19846 31276 19898 31328
rect 50374 31276 50426 31328
rect 50438 31276 50490 31328
rect 50502 31276 50554 31328
rect 50566 31276 50618 31328
rect 45142 30795 45194 30847
rect 17686 30721 17738 30773
rect 4294 30610 4346 30662
rect 4358 30610 4410 30662
rect 4422 30610 4474 30662
rect 4486 30610 4538 30662
rect 35014 30610 35066 30662
rect 35078 30610 35130 30662
rect 35142 30610 35194 30662
rect 35206 30610 35258 30662
rect 25462 30351 25514 30403
rect 29974 30320 30026 30329
rect 29974 30286 29983 30320
rect 29983 30286 30017 30320
rect 30017 30286 30026 30320
rect 29974 30277 30026 30286
rect 19654 29944 19706 29996
rect 19718 29944 19770 29996
rect 19782 29944 19834 29996
rect 19846 29944 19898 29996
rect 50374 29944 50426 29996
rect 50438 29944 50490 29996
rect 50502 29944 50554 29996
rect 50566 29944 50618 29996
rect 6358 29611 6410 29663
rect 55510 29611 55562 29663
rect 1942 29537 1994 29589
rect 14134 29537 14186 29589
rect 11542 29463 11594 29515
rect 17782 29432 17834 29441
rect 17782 29398 17791 29432
rect 17791 29398 17825 29432
rect 17825 29398 17834 29432
rect 17782 29389 17834 29398
rect 19222 29432 19274 29441
rect 19222 29398 19231 29432
rect 19231 29398 19265 29432
rect 19265 29398 19274 29432
rect 19222 29389 19274 29398
rect 40342 29432 40394 29441
rect 40342 29398 40351 29432
rect 40351 29398 40385 29432
rect 40385 29398 40394 29432
rect 40342 29389 40394 29398
rect 49942 29389 49994 29441
rect 50614 29389 50666 29441
rect 54646 29389 54698 29441
rect 55702 29432 55754 29441
rect 55702 29398 55711 29432
rect 55711 29398 55745 29432
rect 55745 29398 55754 29432
rect 55702 29389 55754 29398
rect 4294 29278 4346 29330
rect 4358 29278 4410 29330
rect 4422 29278 4474 29330
rect 4486 29278 4538 29330
rect 35014 29278 35066 29330
rect 35078 29278 35130 29330
rect 35142 29278 35194 29330
rect 35206 29278 35258 29330
rect 9046 29167 9098 29219
rect 14134 29167 14186 29219
rect 8374 29093 8426 29145
rect 22678 29167 22730 29219
rect 50614 29167 50666 29219
rect 55510 29167 55562 29219
rect 41302 28945 41354 28997
rect 15286 28914 15338 28923
rect 15286 28880 15295 28914
rect 15295 28880 15329 28914
rect 15329 28880 15338 28914
rect 15286 28871 15338 28880
rect 44854 28871 44906 28923
rect 8758 28723 8810 28775
rect 19654 28612 19706 28664
rect 19718 28612 19770 28664
rect 19782 28612 19834 28664
rect 19846 28612 19898 28664
rect 50374 28612 50426 28664
rect 50438 28612 50490 28664
rect 50502 28612 50554 28664
rect 50566 28612 50618 28664
rect 2902 28131 2954 28183
rect 20470 28057 20522 28109
rect 41782 28100 41834 28109
rect 41782 28066 41791 28100
rect 41791 28066 41825 28100
rect 41825 28066 41834 28100
rect 41782 28057 41834 28066
rect 4294 27946 4346 27998
rect 4358 27946 4410 27998
rect 4422 27946 4474 27998
rect 4486 27946 4538 27998
rect 35014 27946 35066 27998
rect 35078 27946 35130 27998
rect 35142 27946 35194 27998
rect 35206 27946 35258 27998
rect 7126 27835 7178 27887
rect 26422 27835 26474 27887
rect 41782 27835 41834 27887
rect 8374 27687 8426 27739
rect 14326 27582 14378 27591
rect 14326 27548 14335 27582
rect 14335 27548 14369 27582
rect 14369 27548 14378 27582
rect 14326 27539 14378 27548
rect 25078 27539 25130 27591
rect 8854 27391 8906 27443
rect 19654 27280 19706 27332
rect 19718 27280 19770 27332
rect 19782 27280 19834 27332
rect 19846 27280 19898 27332
rect 50374 27280 50426 27332
rect 50438 27280 50490 27332
rect 50502 27280 50554 27332
rect 50566 27280 50618 27332
rect 24310 26799 24362 26851
rect 7702 26725 7754 26777
rect 28630 26768 28682 26777
rect 28630 26734 28639 26768
rect 28639 26734 28673 26768
rect 28673 26734 28682 26768
rect 28630 26725 28682 26734
rect 4294 26614 4346 26666
rect 4358 26614 4410 26666
rect 4422 26614 4474 26666
rect 4486 26614 4538 26666
rect 35014 26614 35066 26666
rect 35078 26614 35130 26666
rect 35142 26614 35194 26666
rect 35206 26614 35258 26666
rect 8086 26355 8138 26407
rect 7942 26281 7994 26333
rect 24214 26250 24266 26259
rect 24214 26216 24223 26250
rect 24223 26216 24257 26250
rect 24257 26216 24266 26250
rect 24214 26207 24266 26216
rect 36118 26207 36170 26259
rect 16246 26133 16298 26185
rect 9238 26059 9290 26111
rect 19654 25948 19706 26000
rect 19718 25948 19770 26000
rect 19782 25948 19834 26000
rect 19846 25948 19898 26000
rect 50374 25948 50426 26000
rect 50438 25948 50490 26000
rect 50502 25948 50554 26000
rect 50566 25948 50618 26000
rect 55126 25837 55178 25889
rect 14710 25689 14762 25741
rect 5686 25393 5738 25445
rect 37654 25393 37706 25445
rect 4294 25282 4346 25334
rect 4358 25282 4410 25334
rect 4422 25282 4474 25334
rect 4486 25282 4538 25334
rect 35014 25282 35066 25334
rect 35078 25282 35130 25334
rect 35142 25282 35194 25334
rect 35206 25282 35258 25334
rect 9622 25171 9674 25223
rect 8374 24949 8426 25001
rect 9142 24949 9194 25001
rect 7942 24875 7994 24927
rect 8230 24875 8282 24927
rect 14614 24918 14666 24927
rect 14614 24884 14623 24918
rect 14623 24884 14657 24918
rect 14657 24884 14666 24918
rect 14614 24875 14666 24884
rect 49846 24918 49898 24927
rect 49846 24884 49855 24918
rect 49855 24884 49889 24918
rect 49889 24884 49898 24918
rect 49846 24875 49898 24884
rect 52534 24918 52586 24927
rect 52534 24884 52543 24918
rect 52543 24884 52577 24918
rect 52577 24884 52586 24918
rect 52534 24875 52586 24884
rect 19654 24616 19706 24668
rect 19718 24616 19770 24668
rect 19782 24616 19834 24668
rect 19846 24616 19898 24668
rect 50374 24616 50426 24668
rect 50438 24616 50490 24668
rect 50502 24616 50554 24668
rect 50566 24616 50618 24668
rect 8182 24505 8234 24557
rect 8566 24505 8618 24557
rect 5206 24135 5258 24187
rect 34870 24135 34922 24187
rect 8374 24061 8426 24113
rect 8566 24061 8618 24113
rect 11638 24104 11690 24113
rect 11638 24070 11647 24104
rect 11647 24070 11681 24104
rect 11681 24070 11690 24104
rect 11638 24061 11690 24070
rect 30166 24061 30218 24113
rect 4294 23950 4346 24002
rect 4358 23950 4410 24002
rect 4422 23950 4474 24002
rect 4486 23950 4538 24002
rect 35014 23950 35066 24002
rect 35078 23950 35130 24002
rect 35142 23950 35194 24002
rect 35206 23950 35258 24002
rect 7414 23839 7466 23891
rect 7798 23839 7850 23891
rect 15862 23839 15914 23891
rect 34870 23839 34922 23891
rect 8086 23617 8138 23669
rect 8374 23543 8426 23595
rect 12406 23586 12458 23595
rect 12406 23552 12415 23586
rect 12415 23552 12449 23586
rect 12449 23552 12458 23586
rect 12406 23543 12458 23552
rect 36886 23543 36938 23595
rect 42742 23543 42794 23595
rect 7942 23469 7994 23521
rect 19654 23284 19706 23336
rect 19718 23284 19770 23336
rect 19782 23284 19834 23336
rect 19846 23284 19898 23336
rect 50374 23284 50426 23336
rect 50438 23284 50490 23336
rect 50502 23284 50554 23336
rect 50566 23284 50618 23336
rect 7318 23173 7370 23225
rect 8374 23173 8426 23225
rect 7894 22729 7946 22781
rect 8086 22729 8138 22781
rect 12310 22729 12362 22781
rect 42838 22772 42890 22781
rect 42838 22738 42847 22772
rect 42847 22738 42881 22772
rect 42881 22738 42890 22772
rect 42838 22729 42890 22738
rect 4294 22618 4346 22670
rect 4358 22618 4410 22670
rect 4422 22618 4474 22670
rect 4486 22618 4538 22670
rect 35014 22618 35066 22670
rect 35078 22618 35130 22670
rect 35142 22618 35194 22670
rect 35206 22618 35258 22670
rect 7510 22507 7562 22559
rect 7702 22507 7754 22559
rect 8278 22507 8330 22559
rect 8470 22507 8522 22559
rect 7126 22433 7178 22485
rect 7606 22433 7658 22485
rect 7894 22433 7946 22485
rect 7702 22359 7754 22411
rect 28726 22211 28778 22263
rect 34870 22211 34922 22263
rect 36982 22211 37034 22263
rect 8278 22063 8330 22115
rect 19654 21952 19706 22004
rect 19718 21952 19770 22004
rect 19782 21952 19834 22004
rect 19846 21952 19898 22004
rect 50374 21952 50426 22004
rect 50438 21952 50490 22004
rect 50502 21952 50554 22004
rect 50566 21952 50618 22004
rect 8278 21841 8330 21893
rect 14710 21841 14762 21893
rect 22870 21693 22922 21745
rect 8278 21545 8330 21597
rect 43894 21545 43946 21597
rect 10006 21397 10058 21449
rect 4294 21286 4346 21338
rect 4358 21286 4410 21338
rect 4422 21286 4474 21338
rect 4486 21286 4538 21338
rect 35014 21286 35066 21338
rect 35078 21286 35130 21338
rect 35142 21286 35194 21338
rect 35206 21286 35258 21338
rect 57718 21101 57770 21153
rect 8230 20953 8282 21005
rect 15574 20879 15626 20931
rect 28342 20879 28394 20931
rect 10774 20805 10826 20857
rect 8278 20731 8330 20783
rect 9334 20731 9386 20783
rect 16630 20731 16682 20783
rect 19654 20620 19706 20672
rect 19718 20620 19770 20672
rect 19782 20620 19834 20672
rect 19846 20620 19898 20672
rect 50374 20620 50426 20672
rect 50438 20620 50490 20672
rect 50502 20620 50554 20672
rect 50566 20620 50618 20672
rect 8278 20509 8330 20561
rect 9334 20509 9386 20561
rect 10774 20509 10826 20561
rect 53974 20509 54026 20561
rect 30934 20435 30986 20487
rect 27094 20108 27146 20117
rect 27094 20074 27103 20108
rect 27103 20074 27137 20108
rect 27137 20074 27146 20108
rect 27094 20065 27146 20074
rect 53014 20108 53066 20117
rect 53014 20074 53023 20108
rect 53023 20074 53057 20108
rect 53057 20074 53066 20108
rect 53014 20065 53066 20074
rect 4294 19954 4346 20006
rect 4358 19954 4410 20006
rect 4422 19954 4474 20006
rect 4486 19954 4538 20006
rect 35014 19954 35066 20006
rect 35078 19954 35130 20006
rect 35142 19954 35194 20006
rect 35206 19954 35258 20006
rect 53686 19769 53738 19821
rect 27190 19547 27242 19599
rect 8086 19473 8138 19525
rect 16534 19473 16586 19525
rect 19654 19288 19706 19340
rect 19718 19288 19770 19340
rect 19782 19288 19834 19340
rect 19846 19288 19898 19340
rect 50374 19288 50426 19340
rect 50438 19288 50490 19340
rect 50502 19288 50554 19340
rect 50566 19288 50618 19340
rect 8086 19177 8138 19229
rect 50806 19177 50858 19229
rect 7030 18881 7082 18933
rect 7798 18881 7850 18933
rect 7510 18733 7562 18785
rect 7798 18733 7850 18785
rect 22966 18733 23018 18785
rect 4294 18622 4346 18674
rect 4358 18622 4410 18674
rect 4422 18622 4474 18674
rect 4486 18622 4538 18674
rect 35014 18622 35066 18674
rect 35078 18622 35130 18674
rect 35142 18622 35194 18674
rect 35206 18622 35258 18674
rect 8662 18511 8714 18563
rect 8230 18235 8282 18287
rect 34390 18437 34442 18489
rect 20662 18332 20714 18341
rect 20662 18298 20671 18332
rect 20671 18298 20705 18332
rect 20705 18298 20714 18332
rect 20662 18289 20714 18298
rect 48886 18289 48938 18341
rect 46102 18215 46154 18267
rect 50134 18215 50186 18267
rect 44758 18141 44810 18193
rect 7126 18067 7178 18119
rect 7318 18067 7370 18119
rect 8662 18067 8714 18119
rect 19654 17956 19706 18008
rect 19718 17956 19770 18008
rect 19782 17956 19834 18008
rect 19846 17956 19898 18008
rect 50374 17956 50426 18008
rect 50438 17956 50490 18008
rect 50502 17956 50554 18008
rect 50566 17956 50618 18008
rect 8662 17845 8714 17897
rect 9046 17845 9098 17897
rect 8182 17771 8234 17823
rect 42934 17771 42986 17823
rect 48886 17401 48938 17453
rect 4294 17290 4346 17342
rect 4358 17290 4410 17342
rect 4422 17290 4474 17342
rect 4486 17290 4538 17342
rect 35014 17290 35066 17342
rect 35078 17290 35130 17342
rect 35142 17290 35194 17342
rect 35206 17290 35258 17342
rect 7414 17179 7466 17231
rect 9046 17179 9098 17231
rect 42646 17179 42698 17231
rect 39766 17031 39818 17083
rect 24502 16883 24554 16935
rect 19654 16624 19706 16676
rect 19718 16624 19770 16676
rect 19782 16624 19834 16676
rect 19846 16624 19898 16676
rect 50374 16624 50426 16676
rect 50438 16624 50490 16676
rect 50502 16624 50554 16676
rect 50566 16624 50618 16676
rect 7414 16069 7466 16121
rect 8182 16069 8234 16121
rect 4294 15958 4346 16010
rect 4358 15958 4410 16010
rect 4422 15958 4474 16010
rect 4486 15958 4538 16010
rect 35014 15958 35066 16010
rect 35078 15958 35130 16010
rect 35142 15958 35194 16010
rect 35206 15958 35258 16010
rect 7414 15847 7466 15899
rect 8182 15847 8234 15899
rect 20374 15847 20426 15899
rect 38902 15773 38954 15825
rect 27670 15551 27722 15603
rect 8182 15477 8234 15529
rect 19654 15292 19706 15344
rect 19718 15292 19770 15344
rect 19782 15292 19834 15344
rect 19846 15292 19898 15344
rect 50374 15292 50426 15344
rect 50438 15292 50490 15344
rect 50502 15292 50554 15344
rect 50566 15292 50618 15344
rect 8182 15181 8234 15233
rect 36694 15181 36746 15233
rect 7894 15107 7946 15159
rect 8278 15107 8330 15159
rect 18454 14811 18506 14863
rect 24694 14737 24746 14789
rect 4294 14626 4346 14678
rect 4358 14626 4410 14678
rect 4422 14626 4474 14678
rect 4486 14626 4538 14678
rect 35014 14626 35066 14678
rect 35078 14626 35130 14678
rect 35142 14626 35194 14678
rect 35206 14626 35258 14678
rect 53398 14441 53450 14493
rect 51190 14262 51242 14271
rect 51190 14228 51199 14262
rect 51199 14228 51233 14262
rect 51233 14228 51242 14262
rect 51190 14219 51242 14228
rect 25558 14145 25610 14197
rect 36598 14071 36650 14123
rect 19654 13960 19706 14012
rect 19718 13960 19770 14012
rect 19782 13960 19834 14012
rect 19846 13960 19898 14012
rect 50374 13960 50426 14012
rect 50438 13960 50490 14012
rect 50502 13960 50554 14012
rect 50566 13960 50618 14012
rect 15958 13892 16010 13901
rect 15958 13858 15967 13892
rect 15967 13858 16001 13892
rect 16001 13858 16010 13892
rect 15958 13849 16010 13858
rect 3286 13405 3338 13457
rect 8182 13405 8234 13457
rect 11446 13448 11498 13457
rect 11446 13414 11455 13448
rect 11455 13414 11489 13448
rect 11489 13414 11498 13448
rect 11446 13405 11498 13414
rect 45142 13448 45194 13457
rect 45142 13414 45151 13448
rect 45151 13414 45185 13448
rect 45185 13414 45194 13448
rect 45142 13405 45194 13414
rect 4294 13294 4346 13346
rect 4358 13294 4410 13346
rect 4422 13294 4474 13346
rect 4486 13294 4538 13346
rect 35014 13294 35066 13346
rect 35078 13294 35130 13346
rect 35142 13294 35194 13346
rect 35206 13294 35258 13346
rect 7510 13183 7562 13235
rect 8182 13183 8234 13235
rect 45142 13183 45194 13235
rect 56950 13183 57002 13235
rect 7222 12961 7274 13013
rect 33046 13109 33098 13161
rect 56278 12961 56330 13013
rect 30070 12813 30122 12865
rect 19654 12628 19706 12680
rect 19718 12628 19770 12680
rect 19782 12628 19834 12680
rect 19846 12628 19898 12680
rect 50374 12628 50426 12680
rect 50438 12628 50490 12680
rect 50502 12628 50554 12680
rect 50566 12628 50618 12680
rect 7606 12517 7658 12569
rect 7798 12517 7850 12569
rect 57334 12560 57386 12569
rect 57334 12526 57343 12560
rect 57343 12526 57377 12560
rect 57377 12526 57386 12560
rect 57334 12517 57386 12526
rect 10006 12295 10058 12347
rect 17974 12295 18026 12347
rect 57430 12221 57482 12273
rect 10006 12147 10058 12199
rect 6550 12116 6602 12125
rect 6550 12082 6559 12116
rect 6559 12082 6593 12116
rect 6593 12082 6602 12116
rect 6550 12073 6602 12082
rect 13654 12073 13706 12125
rect 57526 12147 57578 12199
rect 4294 11962 4346 12014
rect 4358 11962 4410 12014
rect 4422 11962 4474 12014
rect 4486 11962 4538 12014
rect 35014 11962 35066 12014
rect 35078 11962 35130 12014
rect 35142 11962 35194 12014
rect 35206 11962 35258 12014
rect 7030 11851 7082 11903
rect 7318 11851 7370 11903
rect 29302 11777 29354 11829
rect 17974 11703 18026 11755
rect 25174 11629 25226 11681
rect 27094 11629 27146 11681
rect 24406 11555 24458 11607
rect 54742 11555 54794 11607
rect 58198 11555 58250 11607
rect 57142 11407 57194 11459
rect 19654 11296 19706 11348
rect 19718 11296 19770 11348
rect 19782 11296 19834 11348
rect 19846 11296 19898 11348
rect 50374 11296 50426 11348
rect 50438 11296 50490 11348
rect 50502 11296 50554 11348
rect 50566 11296 50618 11348
rect 7798 11185 7850 11237
rect 8086 11185 8138 11237
rect 8086 11037 8138 11089
rect 22294 11037 22346 11089
rect 28150 11037 28202 11089
rect 17782 10963 17834 11015
rect 9622 10889 9674 10941
rect 26518 10889 26570 10941
rect 29782 10889 29834 10941
rect 56758 10889 56810 10941
rect 4726 10815 4778 10867
rect 34294 10815 34346 10867
rect 56566 10815 56618 10867
rect 7990 10741 8042 10793
rect 11158 10741 11210 10793
rect 31702 10741 31754 10793
rect 48214 10741 48266 10793
rect 4294 10630 4346 10682
rect 4358 10630 4410 10682
rect 4422 10630 4474 10682
rect 4486 10630 4538 10682
rect 35014 10630 35066 10682
rect 35078 10630 35130 10682
rect 35142 10630 35194 10682
rect 35206 10630 35258 10682
rect 8182 10519 8234 10571
rect 8470 10519 8522 10571
rect 33814 10519 33866 10571
rect 48214 10519 48266 10571
rect 56470 10519 56522 10571
rect 9622 10445 9674 10497
rect 8086 10371 8138 10423
rect 55894 10414 55946 10423
rect 55894 10380 55903 10414
rect 55903 10380 55937 10414
rect 55937 10380 55946 10414
rect 55894 10371 55946 10380
rect 11638 10297 11690 10349
rect 55702 10297 55754 10349
rect 9142 10223 9194 10275
rect 9334 10223 9386 10275
rect 41494 10223 41546 10275
rect 56470 10223 56522 10275
rect 8758 10075 8810 10127
rect 9142 10075 9194 10127
rect 58582 10149 58634 10201
rect 55702 10075 55754 10127
rect 56086 10075 56138 10127
rect 19654 9964 19706 10016
rect 19718 9964 19770 10016
rect 19782 9964 19834 10016
rect 19846 9964 19898 10016
rect 50374 9964 50426 10016
rect 50438 9964 50490 10016
rect 50502 9964 50554 10016
rect 50566 9964 50618 10016
rect 7030 9853 7082 9905
rect 8758 9853 8810 9905
rect 23446 9853 23498 9905
rect 54934 9853 54986 9905
rect 55318 9853 55370 9905
rect 7990 9779 8042 9831
rect 9622 9779 9674 9831
rect 41590 9779 41642 9831
rect 49078 9779 49130 9831
rect 55606 9822 55658 9831
rect 55606 9788 55615 9822
rect 55615 9788 55649 9822
rect 55649 9788 55658 9822
rect 55606 9779 55658 9788
rect 8278 9705 8330 9757
rect 16150 9705 16202 9757
rect 41782 9705 41834 9757
rect 49942 9705 49994 9757
rect 3382 9631 3434 9683
rect 39574 9631 39626 9683
rect 8374 9557 8426 9609
rect 8566 9557 8618 9609
rect 28630 9557 28682 9609
rect 57622 9674 57674 9683
rect 57622 9640 57631 9674
rect 57631 9640 57665 9674
rect 57665 9640 57674 9674
rect 57622 9631 57674 9640
rect 54262 9557 54314 9609
rect 54454 9600 54506 9609
rect 54454 9566 54463 9600
rect 54463 9566 54497 9600
rect 54497 9566 54506 9600
rect 54454 9557 54506 9566
rect 8086 9483 8138 9535
rect 17878 9483 17930 9535
rect 57814 9483 57866 9535
rect 8566 9409 8618 9461
rect 19318 9409 19370 9461
rect 47542 9409 47594 9461
rect 52630 9452 52682 9461
rect 52630 9418 52639 9452
rect 52639 9418 52673 9452
rect 52673 9418 52682 9452
rect 52630 9409 52682 9418
rect 4294 9298 4346 9350
rect 4358 9298 4410 9350
rect 4422 9298 4474 9350
rect 4486 9298 4538 9350
rect 35014 9298 35066 9350
rect 35078 9298 35130 9350
rect 35142 9298 35194 9350
rect 35206 9298 35258 9350
rect 7030 9187 7082 9239
rect 8278 9187 8330 9239
rect 20950 9187 21002 9239
rect 52630 9187 52682 9239
rect 8566 9113 8618 9165
rect 8758 9113 8810 9165
rect 39574 9156 39626 9165
rect 39574 9122 39583 9156
rect 39583 9122 39617 9156
rect 39617 9122 39626 9156
rect 39574 9113 39626 9122
rect 40630 9113 40682 9165
rect 49846 9113 49898 9165
rect 54454 9113 54506 9165
rect 12598 9039 12650 9091
rect 15670 9039 15722 9091
rect 54646 9082 54698 9091
rect 8086 8965 8138 9017
rect 9046 8965 9098 9017
rect 20854 8965 20906 9017
rect 40054 8965 40106 9017
rect 53398 9008 53450 9017
rect 53398 8974 53407 9008
rect 53407 8974 53441 9008
rect 53441 8974 53450 9008
rect 53398 8965 53450 8974
rect 5206 8891 5258 8943
rect 8662 8891 8714 8943
rect 11254 8891 11306 8943
rect 11446 8891 11498 8943
rect 13174 8891 13226 8943
rect 32278 8891 32330 8943
rect 42934 8891 42986 8943
rect 44662 8891 44714 8943
rect 54646 9048 54655 9082
rect 54655 9048 54689 9082
rect 54689 9048 54698 9082
rect 54646 9039 54698 9048
rect 54550 8965 54602 9017
rect 57238 9008 57290 9017
rect 57238 8974 57247 9008
rect 57247 8974 57281 9008
rect 57281 8974 57290 9008
rect 57238 8965 57290 8974
rect 9046 8817 9098 8869
rect 10966 8817 11018 8869
rect 11350 8817 11402 8869
rect 13942 8817 13994 8869
rect 16150 8817 16202 8869
rect 17014 8817 17066 8869
rect 57334 8891 57386 8943
rect 9430 8743 9482 8795
rect 14998 8743 15050 8795
rect 23062 8743 23114 8795
rect 29014 8743 29066 8795
rect 36214 8743 36266 8795
rect 46390 8743 46442 8795
rect 55990 8817 56042 8869
rect 53878 8743 53930 8795
rect 19654 8632 19706 8684
rect 19718 8632 19770 8684
rect 19782 8632 19834 8684
rect 19846 8632 19898 8684
rect 50374 8632 50426 8684
rect 50438 8632 50490 8684
rect 50502 8632 50554 8684
rect 50566 8632 50618 8684
rect 3766 8521 3818 8573
rect 9622 8521 9674 8573
rect 10870 8521 10922 8573
rect 11542 8521 11594 8573
rect 12502 8521 12554 8573
rect 29206 8521 29258 8573
rect 31222 8521 31274 8573
rect 42646 8521 42698 8573
rect 46486 8521 46538 8573
rect 47926 8521 47978 8573
rect 52342 8521 52394 8573
rect 58966 8521 59018 8573
rect 7606 8447 7658 8499
rect 3286 8416 3338 8425
rect 3286 8382 3295 8416
rect 3295 8382 3329 8416
rect 3329 8382 3338 8416
rect 3286 8373 3338 8382
rect 1654 8268 1706 8277
rect 1654 8234 1663 8268
rect 1663 8234 1697 8268
rect 1697 8234 1706 8268
rect 1654 8225 1706 8234
rect 2134 8225 2186 8277
rect 3286 8225 3338 8277
rect 12214 8373 12266 8425
rect 7606 8225 7658 8277
rect 7702 8225 7754 8277
rect 8566 8225 8618 8277
rect 4822 8151 4874 8203
rect 5590 8151 5642 8203
rect 9430 8151 9482 8203
rect 9526 8151 9578 8203
rect 12502 8299 12554 8351
rect 12598 8342 12650 8351
rect 12598 8308 12607 8342
rect 12607 8308 12641 8342
rect 12641 8308 12650 8342
rect 12598 8299 12650 8308
rect 10294 8225 10346 8277
rect 10678 8225 10730 8277
rect 11446 8225 11498 8277
rect 12118 8268 12170 8277
rect 12118 8234 12127 8268
rect 12127 8234 12161 8268
rect 12161 8234 12170 8268
rect 12118 8225 12170 8234
rect 12982 8151 13034 8203
rect 13174 8447 13226 8499
rect 13654 8416 13706 8425
rect 13654 8382 13663 8416
rect 13663 8382 13697 8416
rect 13697 8382 13706 8416
rect 13654 8373 13706 8382
rect 16342 8373 16394 8425
rect 20566 8373 20618 8425
rect 16054 8299 16106 8351
rect 16438 8299 16490 8351
rect 38038 8299 38090 8351
rect 13174 8225 13226 8277
rect 14806 8225 14858 8277
rect 15958 8225 16010 8277
rect 16246 8268 16298 8277
rect 16246 8234 16255 8268
rect 16255 8234 16289 8268
rect 16289 8234 16298 8268
rect 16246 8225 16298 8234
rect 16342 8225 16394 8277
rect 17014 8268 17066 8277
rect 17014 8234 17023 8268
rect 17023 8234 17057 8268
rect 17057 8234 17066 8268
rect 17014 8225 17066 8234
rect 18838 8225 18890 8277
rect 46102 8373 46154 8425
rect 38230 8299 38282 8351
rect 48886 8416 48938 8425
rect 48886 8382 48895 8416
rect 48895 8382 48929 8416
rect 48929 8382 48938 8416
rect 48886 8373 48938 8382
rect 46390 8299 46442 8351
rect 38806 8225 38858 8277
rect 47542 8225 47594 8277
rect 48022 8225 48074 8277
rect 48694 8225 48746 8277
rect 49462 8225 49514 8277
rect 25654 8151 25706 8203
rect 29782 8194 29834 8203
rect 4918 8077 4970 8129
rect 24214 8077 24266 8129
rect 24406 8077 24458 8129
rect 29302 8077 29354 8129
rect 29782 8160 29791 8194
rect 29791 8160 29825 8194
rect 29825 8160 29834 8194
rect 29782 8151 29834 8160
rect 29974 8077 30026 8129
rect 32950 8077 33002 8129
rect 33238 8077 33290 8129
rect 39574 8077 39626 8129
rect 41110 8077 41162 8129
rect 46006 8077 46058 8129
rect 52918 8342 52970 8351
rect 52918 8308 52927 8342
rect 52927 8308 52961 8342
rect 52961 8308 52970 8342
rect 52918 8299 52970 8308
rect 53110 8151 53162 8203
rect 53494 8225 53546 8277
rect 54070 8268 54122 8277
rect 54070 8234 54079 8268
rect 54079 8234 54113 8268
rect 54113 8234 54122 8268
rect 54070 8225 54122 8234
rect 56950 8299 57002 8351
rect 58390 8225 58442 8277
rect 59830 8151 59882 8203
rect 54742 8077 54794 8129
rect 4294 7966 4346 8018
rect 4358 7966 4410 8018
rect 4422 7966 4474 8018
rect 4486 7966 4538 8018
rect 35014 7966 35066 8018
rect 35078 7966 35130 8018
rect 35142 7966 35194 8018
rect 35206 7966 35258 8018
rect 3670 7898 3722 7907
rect 3670 7864 3679 7898
rect 3679 7864 3713 7898
rect 3713 7864 3722 7898
rect 3670 7855 3722 7864
rect 3382 7707 3434 7759
rect 7894 7855 7946 7907
rect 4918 7707 4970 7759
rect 5590 7750 5642 7759
rect 5590 7716 5599 7750
rect 5599 7716 5633 7750
rect 5633 7716 5642 7750
rect 5590 7707 5642 7716
rect 9718 7855 9770 7907
rect 9910 7855 9962 7907
rect 10006 7781 10058 7833
rect 11446 7781 11498 7833
rect 9430 7750 9482 7759
rect 9430 7716 9439 7750
rect 9439 7716 9473 7750
rect 9473 7716 9482 7750
rect 9430 7707 9482 7716
rect 10198 7750 10250 7759
rect 10198 7716 10207 7750
rect 10207 7716 10241 7750
rect 10241 7716 10250 7750
rect 10198 7707 10250 7716
rect 1462 7633 1514 7685
rect 8518 7633 8570 7685
rect 8758 7633 8810 7685
rect 11926 7707 11978 7759
rect 12118 7855 12170 7907
rect 11062 7633 11114 7685
rect 15958 7855 16010 7907
rect 25942 7898 25994 7907
rect 25654 7781 25706 7833
rect 13270 7707 13322 7759
rect 15382 7707 15434 7759
rect 15766 7750 15818 7759
rect 15766 7716 15775 7750
rect 15775 7716 15809 7750
rect 15809 7716 15818 7750
rect 15766 7707 15818 7716
rect 16150 7707 16202 7759
rect 20950 7750 21002 7759
rect 20950 7716 20959 7750
rect 20959 7716 20993 7750
rect 20993 7716 21002 7750
rect 20950 7707 21002 7716
rect 24022 7707 24074 7759
rect 24694 7750 24746 7759
rect 24694 7716 24703 7750
rect 24703 7716 24737 7750
rect 24737 7716 24746 7750
rect 24694 7707 24746 7716
rect 25462 7750 25514 7759
rect 25462 7716 25471 7750
rect 25471 7716 25505 7750
rect 25505 7716 25514 7750
rect 25462 7707 25514 7716
rect 15478 7633 15530 7685
rect 15670 7633 15722 7685
rect 21046 7633 21098 7685
rect 25270 7633 25322 7685
rect 25654 7633 25706 7685
rect 25942 7864 25951 7898
rect 25951 7864 25985 7898
rect 25985 7864 25994 7898
rect 29110 7898 29162 7907
rect 25942 7855 25994 7864
rect 29110 7864 29119 7898
rect 29119 7864 29153 7898
rect 29153 7864 29162 7898
rect 29110 7855 29162 7864
rect 29206 7855 29258 7907
rect 34870 7855 34922 7907
rect 26230 7781 26282 7833
rect 29302 7781 29354 7833
rect 30166 7750 30218 7759
rect 30166 7716 30175 7750
rect 30175 7716 30209 7750
rect 30209 7716 30218 7750
rect 30166 7707 30218 7716
rect 30838 7750 30890 7759
rect 30838 7716 30847 7750
rect 30847 7716 30881 7750
rect 30881 7716 30890 7750
rect 30838 7707 30890 7716
rect 28534 7633 28586 7685
rect 34582 7750 34634 7759
rect 34582 7716 34591 7750
rect 34591 7716 34625 7750
rect 34625 7716 34634 7750
rect 34582 7707 34634 7716
rect 36118 7750 36170 7759
rect 36118 7716 36127 7750
rect 36127 7716 36161 7750
rect 36161 7716 36170 7750
rect 36118 7707 36170 7716
rect 36886 7750 36938 7759
rect 36886 7716 36895 7750
rect 36895 7716 36929 7750
rect 36929 7716 36938 7750
rect 36886 7707 36938 7716
rect 38806 7750 38858 7759
rect 38806 7716 38815 7750
rect 38815 7716 38849 7750
rect 38849 7716 38858 7750
rect 38806 7707 38858 7716
rect 39574 7750 39626 7759
rect 39574 7716 39583 7750
rect 39583 7716 39617 7750
rect 39617 7716 39626 7750
rect 39574 7707 39626 7716
rect 41110 7750 41162 7759
rect 41110 7716 41119 7750
rect 41119 7716 41153 7750
rect 41153 7716 41162 7750
rect 41110 7707 41162 7716
rect 44182 7781 44234 7833
rect 44374 7855 44426 7907
rect 45238 7898 45290 7907
rect 44662 7781 44714 7833
rect 42646 7750 42698 7759
rect 42646 7716 42655 7750
rect 42655 7716 42689 7750
rect 42689 7716 42698 7750
rect 42646 7707 42698 7716
rect 45238 7864 45247 7898
rect 45247 7864 45281 7898
rect 45281 7864 45290 7898
rect 45238 7855 45290 7864
rect 46006 7781 46058 7833
rect 51190 7855 51242 7907
rect 51862 7855 51914 7907
rect 53014 7855 53066 7907
rect 46486 7781 46538 7833
rect 47254 7707 47306 7759
rect 48406 7707 48458 7759
rect 2518 7602 2570 7611
rect 2518 7568 2527 7602
rect 2527 7568 2561 7602
rect 2561 7568 2570 7602
rect 2518 7559 2570 7568
rect 13942 7602 13994 7611
rect 13942 7568 13951 7602
rect 13951 7568 13985 7602
rect 13985 7568 13994 7602
rect 13942 7559 13994 7568
rect 14614 7559 14666 7611
rect 18838 7559 18890 7611
rect 27094 7559 27146 7611
rect 29686 7559 29738 7611
rect 33814 7602 33866 7611
rect 33814 7568 33823 7602
rect 33823 7568 33857 7602
rect 33857 7568 33866 7602
rect 33814 7559 33866 7568
rect 35254 7633 35306 7685
rect 35446 7633 35498 7685
rect 35158 7559 35210 7611
rect 8758 7485 8810 7537
rect 9910 7485 9962 7537
rect 2326 7411 2378 7463
rect 2998 7411 3050 7463
rect 3958 7454 4010 7463
rect 3958 7420 3967 7454
rect 3967 7420 4001 7454
rect 4001 7420 4010 7454
rect 3958 7411 4010 7420
rect 4054 7411 4106 7463
rect 5302 7411 5354 7463
rect 7606 7454 7658 7463
rect 7606 7420 7615 7454
rect 7615 7420 7649 7454
rect 7649 7420 7658 7454
rect 7606 7411 7658 7420
rect 8566 7411 8618 7463
rect 9142 7411 9194 7463
rect 11734 7485 11786 7537
rect 11062 7411 11114 7463
rect 12598 7485 12650 7537
rect 15286 7485 15338 7537
rect 28534 7485 28586 7537
rect 35542 7559 35594 7611
rect 40054 7485 40106 7537
rect 46006 7602 46058 7611
rect 46006 7568 46015 7602
rect 46015 7568 46049 7602
rect 46049 7568 46058 7602
rect 46006 7559 46058 7568
rect 47638 7559 47690 7611
rect 50134 7750 50186 7759
rect 50134 7716 50143 7750
rect 50143 7716 50177 7750
rect 50177 7716 50186 7750
rect 50134 7707 50186 7716
rect 59350 7781 59402 7833
rect 51766 7750 51818 7759
rect 51766 7716 51775 7750
rect 51775 7716 51809 7750
rect 51809 7716 51818 7750
rect 51766 7707 51818 7716
rect 52822 7707 52874 7759
rect 51862 7559 51914 7611
rect 53206 7633 53258 7685
rect 58774 7707 58826 7759
rect 55798 7676 55850 7685
rect 55798 7642 55807 7676
rect 55807 7642 55841 7676
rect 55841 7642 55850 7676
rect 55798 7633 55850 7642
rect 56182 7633 56234 7685
rect 56854 7633 56906 7685
rect 56278 7559 56330 7611
rect 13174 7411 13226 7463
rect 15574 7411 15626 7463
rect 15670 7411 15722 7463
rect 20758 7411 20810 7463
rect 23734 7411 23786 7463
rect 24118 7411 24170 7463
rect 24790 7411 24842 7463
rect 25942 7411 25994 7463
rect 26710 7411 26762 7463
rect 28150 7411 28202 7463
rect 29206 7411 29258 7463
rect 29590 7411 29642 7463
rect 31126 7411 31178 7463
rect 33622 7411 33674 7463
rect 34390 7411 34442 7463
rect 34870 7411 34922 7463
rect 35830 7411 35882 7463
rect 36598 7411 36650 7463
rect 38038 7411 38090 7463
rect 38806 7411 38858 7463
rect 39574 7411 39626 7463
rect 41398 7411 41450 7463
rect 42454 7411 42506 7463
rect 43894 7411 43946 7463
rect 44662 7411 44714 7463
rect 45046 7411 45098 7463
rect 45814 7411 45866 7463
rect 46486 7411 46538 7463
rect 47638 7454 47690 7463
rect 47638 7420 47647 7454
rect 47647 7420 47681 7454
rect 47681 7420 47690 7454
rect 47638 7411 47690 7420
rect 50038 7454 50090 7463
rect 50038 7420 50047 7454
rect 50047 7420 50081 7454
rect 50081 7420 50090 7454
rect 50038 7411 50090 7420
rect 51766 7411 51818 7463
rect 52342 7411 52394 7463
rect 19654 7300 19706 7352
rect 19718 7300 19770 7352
rect 19782 7300 19834 7352
rect 19846 7300 19898 7352
rect 50374 7300 50426 7352
rect 50438 7300 50490 7352
rect 50502 7300 50554 7352
rect 50566 7300 50618 7352
rect 3670 7115 3722 7167
rect 6550 7189 6602 7241
rect 6934 7189 6986 7241
rect 7606 7189 7658 7241
rect 8566 7189 8618 7241
rect 12790 7189 12842 7241
rect 5398 7041 5450 7093
rect 8758 7041 8810 7093
rect 9526 7041 9578 7093
rect 10054 7115 10106 7167
rect 12310 7115 12362 7167
rect 29302 7189 29354 7241
rect 29494 7189 29546 7241
rect 54070 7189 54122 7241
rect 1654 7010 1706 7019
rect 1654 6976 1663 7010
rect 1663 6976 1697 7010
rect 1697 6976 1706 7010
rect 1654 6967 1706 6976
rect 2518 7010 2570 7019
rect 2518 6976 2527 7010
rect 2527 6976 2561 7010
rect 2561 6976 2570 7010
rect 2518 6967 2570 6976
rect 7606 7010 7658 7019
rect 7606 6976 7615 7010
rect 7615 6976 7649 7010
rect 7649 6976 7658 7010
rect 7606 6967 7658 6976
rect 9814 7010 9866 7019
rect 9814 6976 9823 7010
rect 9823 6976 9857 7010
rect 9857 6976 9866 7010
rect 9814 6967 9866 6976
rect 10870 6967 10922 7019
rect 11254 7010 11306 7019
rect 11254 6976 11263 7010
rect 11263 6976 11297 7010
rect 11297 6976 11306 7010
rect 11254 6967 11306 6976
rect 12214 7084 12266 7093
rect 12214 7050 12223 7084
rect 12223 7050 12257 7084
rect 12257 7050 12266 7084
rect 12214 7041 12266 7050
rect 13174 7115 13226 7167
rect 14230 7115 14282 7167
rect 15286 7115 15338 7167
rect 19030 7115 19082 7167
rect 13078 7041 13130 7093
rect 20182 7041 20234 7093
rect 20470 7115 20522 7167
rect 23062 7115 23114 7167
rect 23158 7115 23210 7167
rect 25174 7115 25226 7167
rect 25366 7158 25418 7167
rect 25366 7124 25375 7158
rect 25375 7124 25409 7158
rect 25409 7124 25418 7158
rect 25366 7115 25418 7124
rect 25654 7115 25706 7167
rect 21910 7084 21962 7093
rect 21910 7050 21919 7084
rect 21919 7050 21953 7084
rect 21953 7050 21962 7084
rect 21910 7041 21962 7050
rect 22678 7084 22730 7093
rect 22678 7050 22687 7084
rect 22687 7050 22721 7084
rect 22721 7050 22730 7084
rect 22678 7041 22730 7050
rect 23926 7041 23978 7093
rect 26422 7084 26474 7093
rect 26422 7050 26431 7084
rect 26431 7050 26465 7084
rect 26465 7050 26474 7084
rect 26422 7041 26474 7050
rect 26902 7041 26954 7093
rect 27286 7115 27338 7167
rect 30742 7115 30794 7167
rect 31318 7158 31370 7167
rect 27190 7084 27242 7093
rect 27190 7050 27199 7084
rect 27199 7050 27233 7084
rect 27233 7050 27242 7084
rect 27190 7041 27242 7050
rect 28726 7084 28778 7093
rect 28726 7050 28735 7084
rect 28735 7050 28769 7084
rect 28769 7050 28778 7084
rect 28726 7041 28778 7050
rect 29782 7041 29834 7093
rect 29878 7041 29930 7093
rect 31030 7041 31082 7093
rect 31318 7124 31327 7158
rect 31327 7124 31361 7158
rect 31361 7124 31370 7158
rect 31318 7115 31370 7124
rect 31510 7041 31562 7093
rect 32854 7115 32906 7167
rect 39382 7115 39434 7167
rect 39862 7115 39914 7167
rect 41686 7115 41738 7167
rect 51670 7158 51722 7167
rect 51670 7124 51679 7158
rect 51679 7124 51713 7158
rect 51713 7124 51722 7158
rect 51670 7115 51722 7124
rect 32662 7041 32714 7093
rect 34774 7084 34826 7093
rect 12694 7010 12746 7019
rect 12694 6976 12703 7010
rect 12703 6976 12737 7010
rect 12737 6976 12746 7010
rect 12694 6967 12746 6976
rect 12982 6967 13034 7019
rect 27094 6967 27146 7019
rect 29686 6967 29738 7019
rect 34486 6967 34538 7019
rect 34774 7050 34783 7084
rect 34783 7050 34817 7084
rect 34817 7050 34826 7084
rect 34774 7041 34826 7050
rect 36982 7084 37034 7093
rect 36694 6967 36746 7019
rect 36982 7050 36991 7084
rect 36991 7050 37025 7084
rect 37025 7050 37034 7084
rect 36982 7041 37034 7050
rect 41782 7041 41834 7093
rect 42262 7084 42314 7093
rect 42262 7050 42271 7084
rect 42271 7050 42305 7084
rect 42305 7050 42314 7084
rect 42262 7041 42314 7050
rect 44470 7084 44522 7093
rect 44470 7050 44479 7084
rect 44479 7050 44513 7084
rect 44513 7050 44522 7084
rect 44470 7041 44522 7050
rect 48310 7084 48362 7093
rect 48310 7050 48319 7084
rect 48319 7050 48353 7084
rect 48353 7050 48362 7084
rect 48310 7041 48362 7050
rect 50230 7084 50282 7093
rect 50230 7050 50239 7084
rect 50239 7050 50273 7084
rect 50273 7050 50282 7084
rect 50230 7041 50282 7050
rect 38326 6967 38378 7019
rect 38614 6967 38666 7019
rect 4534 6936 4586 6945
rect 4534 6902 4543 6936
rect 4543 6902 4577 6936
rect 4577 6902 4586 6936
rect 4534 6893 4586 6902
rect 5878 6893 5930 6945
rect 6166 6893 6218 6945
rect 6550 6893 6602 6945
rect 5014 6819 5066 6871
rect 7318 6819 7370 6871
rect 9526 6893 9578 6945
rect 9718 6936 9770 6945
rect 9718 6902 9727 6936
rect 9727 6902 9761 6936
rect 9761 6902 9770 6936
rect 9718 6893 9770 6902
rect 9910 6893 9962 6945
rect 10582 6936 10634 6945
rect 10582 6902 10591 6936
rect 10591 6902 10625 6936
rect 10625 6902 10634 6936
rect 10582 6893 10634 6902
rect 13462 6893 13514 6945
rect 14518 6893 14570 6945
rect 14614 6893 14666 6945
rect 15286 6893 15338 6945
rect 15382 6893 15434 6945
rect 15862 6936 15914 6945
rect 15862 6902 15871 6936
rect 15871 6902 15905 6936
rect 15905 6902 15914 6936
rect 15862 6893 15914 6902
rect 17110 6893 17162 6945
rect 17302 6936 17354 6945
rect 17302 6902 17311 6936
rect 17311 6902 17345 6936
rect 17345 6902 17354 6936
rect 17782 6936 17834 6945
rect 17302 6893 17354 6902
rect 17782 6902 17791 6936
rect 17791 6902 17825 6936
rect 17825 6902 17834 6936
rect 17782 6893 17834 6902
rect 17878 6893 17930 6945
rect 18166 6893 18218 6945
rect 18550 6893 18602 6945
rect 10006 6862 10058 6871
rect 10006 6828 10015 6862
rect 10015 6828 10049 6862
rect 10049 6828 10058 6862
rect 10006 6819 10058 6828
rect 19222 6893 19274 6945
rect 20086 6893 20138 6945
rect 20278 6936 20330 6945
rect 20278 6902 20287 6936
rect 20287 6902 20321 6936
rect 20321 6902 20330 6936
rect 20278 6893 20330 6902
rect 20470 6893 20522 6945
rect 20854 6893 20906 6945
rect 21814 6936 21866 6945
rect 21814 6902 21823 6936
rect 21823 6902 21857 6936
rect 21857 6902 21866 6936
rect 21814 6893 21866 6902
rect 21910 6893 21962 6945
rect 22678 6893 22730 6945
rect 23542 6893 23594 6945
rect 17494 6745 17546 6797
rect 18934 6819 18986 6871
rect 23830 6819 23882 6871
rect 22870 6745 22922 6797
rect 23350 6745 23402 6797
rect 24598 6893 24650 6945
rect 25654 6936 25706 6945
rect 25654 6902 25663 6936
rect 25663 6902 25697 6936
rect 25697 6902 25706 6936
rect 26326 6936 26378 6945
rect 25654 6893 25706 6902
rect 26326 6902 26335 6936
rect 26335 6902 26369 6936
rect 26369 6902 26378 6936
rect 26326 6893 26378 6902
rect 26998 6819 27050 6871
rect 27958 6936 28010 6945
rect 27958 6902 27967 6936
rect 27967 6902 28001 6936
rect 28001 6902 28010 6936
rect 28630 6936 28682 6945
rect 27958 6893 28010 6902
rect 28630 6902 28639 6936
rect 28639 6902 28673 6936
rect 28673 6902 28682 6936
rect 28630 6893 28682 6902
rect 28534 6745 28586 6797
rect 29974 6893 30026 6945
rect 31990 6893 32042 6945
rect 32374 6936 32426 6945
rect 32374 6902 32383 6936
rect 32383 6902 32417 6936
rect 32417 6902 32426 6936
rect 32374 6893 32426 6902
rect 32470 6893 32522 6945
rect 33910 6936 33962 6945
rect 33910 6902 33919 6936
rect 33919 6902 33953 6936
rect 33953 6902 33962 6936
rect 33910 6893 33962 6902
rect 34102 6893 34154 6945
rect 34198 6893 34250 6945
rect 35542 6893 35594 6945
rect 36406 6893 36458 6945
rect 36982 6893 37034 6945
rect 37750 6936 37802 6945
rect 37750 6902 37759 6936
rect 37759 6902 37793 6936
rect 37793 6902 37802 6936
rect 37750 6893 37802 6902
rect 30070 6819 30122 6871
rect 33814 6819 33866 6871
rect 34582 6819 34634 6871
rect 37270 6819 37322 6871
rect 37366 6819 37418 6871
rect 38518 6936 38570 6945
rect 38518 6902 38527 6936
rect 38527 6902 38561 6936
rect 38561 6902 38570 6936
rect 41590 6967 41642 7019
rect 38518 6893 38570 6902
rect 29782 6745 29834 6797
rect 33238 6745 33290 6797
rect 34102 6745 34154 6797
rect 35446 6745 35498 6797
rect 37654 6745 37706 6797
rect 40630 6893 40682 6945
rect 39286 6819 39338 6871
rect 42070 6893 42122 6945
rect 41590 6819 41642 6871
rect 39382 6745 39434 6797
rect 42358 6745 42410 6797
rect 42646 6745 42698 6797
rect 43222 6967 43274 7019
rect 46870 6967 46922 7019
rect 43126 6819 43178 6871
rect 44278 6893 44330 6945
rect 44374 6893 44426 6945
rect 45334 6936 45386 6945
rect 45334 6902 45343 6936
rect 45343 6902 45377 6936
rect 45377 6902 45386 6936
rect 45334 6893 45386 6902
rect 46390 6893 46442 6945
rect 45622 6819 45674 6871
rect 47158 6893 47210 6945
rect 48502 6967 48554 7019
rect 54742 7010 54794 7019
rect 47062 6819 47114 6871
rect 48310 6893 48362 6945
rect 50134 6819 50186 6871
rect 51478 6893 51530 6945
rect 52726 6936 52778 6945
rect 52726 6902 52735 6936
rect 52735 6902 52769 6936
rect 52769 6902 52778 6936
rect 52726 6893 52778 6902
rect 54742 6976 54751 7010
rect 54751 6976 54785 7010
rect 54785 6976 54794 7010
rect 54742 6967 54794 6976
rect 55414 6967 55466 7019
rect 58486 6967 58538 7019
rect 50422 6819 50474 6871
rect 56278 6893 56330 6945
rect 46390 6788 46442 6797
rect 46390 6754 46399 6788
rect 46399 6754 46433 6788
rect 46433 6754 46442 6788
rect 46390 6745 46442 6754
rect 47158 6788 47210 6797
rect 47158 6754 47167 6788
rect 47167 6754 47201 6788
rect 47201 6754 47210 6788
rect 47158 6745 47210 6754
rect 4294 6634 4346 6686
rect 4358 6634 4410 6686
rect 4422 6634 4474 6686
rect 4486 6634 4538 6686
rect 35014 6634 35066 6686
rect 35078 6634 35130 6686
rect 35142 6634 35194 6686
rect 35206 6634 35258 6686
rect 6838 6566 6890 6575
rect 6838 6532 6847 6566
rect 6847 6532 6881 6566
rect 6881 6532 6890 6566
rect 6838 6523 6890 6532
rect 5686 6418 5738 6427
rect 5686 6384 5695 6418
rect 5695 6384 5729 6418
rect 5729 6384 5738 6418
rect 5686 6375 5738 6384
rect 8854 6523 8906 6575
rect 10582 6523 10634 6575
rect 10966 6523 11018 6575
rect 13846 6523 13898 6575
rect 14518 6523 14570 6575
rect 8950 6449 9002 6501
rect 11158 6449 11210 6501
rect 17494 6523 17546 6575
rect 24022 6523 24074 6575
rect 1558 6344 1610 6353
rect 1558 6310 1567 6344
rect 1567 6310 1601 6344
rect 1601 6310 1610 6344
rect 1558 6301 1610 6310
rect 2038 6301 2090 6353
rect 3190 6344 3242 6353
rect 3190 6310 3199 6344
rect 3199 6310 3233 6344
rect 3233 6310 3242 6344
rect 3190 6301 3242 6310
rect 3862 6301 3914 6353
rect 4630 6301 4682 6353
rect 5110 6301 5162 6353
rect 8374 6375 8426 6427
rect 9622 6375 9674 6427
rect 9430 6344 9482 6353
rect 9430 6310 9439 6344
rect 9439 6310 9473 6344
rect 9473 6310 9482 6344
rect 9430 6301 9482 6310
rect 10102 6301 10154 6353
rect 10870 6301 10922 6353
rect 11638 6301 11690 6353
rect 12310 6301 12362 6353
rect 13846 6418 13898 6427
rect 13846 6384 13855 6418
rect 13855 6384 13889 6418
rect 13889 6384 13898 6418
rect 14710 6418 14762 6427
rect 13846 6375 13898 6384
rect 14710 6384 14719 6418
rect 14719 6384 14753 6418
rect 14753 6384 14762 6418
rect 14710 6375 14762 6384
rect 15094 6418 15146 6427
rect 15094 6384 15103 6418
rect 15103 6384 15137 6418
rect 15137 6384 15146 6418
rect 15094 6375 15146 6384
rect 16726 6375 16778 6427
rect 17686 6375 17738 6427
rect 18454 6418 18506 6427
rect 18454 6384 18463 6418
rect 18463 6384 18497 6418
rect 18497 6384 18506 6418
rect 18454 6375 18506 6384
rect 19030 6449 19082 6501
rect 25174 6449 25226 6501
rect 27670 6449 27722 6501
rect 27958 6523 28010 6575
rect 28630 6523 28682 6575
rect 28822 6523 28874 6575
rect 29110 6523 29162 6575
rect 32278 6523 32330 6575
rect 33526 6523 33578 6575
rect 19606 6375 19658 6427
rect 19990 6418 20042 6427
rect 19990 6384 19999 6418
rect 19999 6384 20033 6418
rect 20033 6384 20042 6418
rect 19990 6375 20042 6384
rect 20086 6375 20138 6427
rect 24502 6418 24554 6427
rect 17302 6301 17354 6353
rect 9046 6227 9098 6279
rect 12982 6227 13034 6279
rect 19318 6301 19370 6353
rect 24502 6384 24511 6418
rect 24511 6384 24545 6418
rect 24545 6384 24554 6418
rect 24502 6375 24554 6384
rect 28246 6418 28298 6427
rect 28246 6384 28255 6418
rect 28255 6384 28289 6418
rect 28289 6384 28298 6418
rect 28246 6375 28298 6384
rect 29014 6418 29066 6427
rect 29014 6384 29023 6418
rect 29023 6384 29057 6418
rect 29057 6384 29066 6418
rect 29014 6375 29066 6384
rect 30646 6418 30698 6427
rect 30646 6384 30655 6418
rect 30655 6384 30689 6418
rect 30689 6384 30698 6418
rect 30646 6375 30698 6384
rect 30742 6375 30794 6427
rect 25654 6344 25706 6353
rect 8758 6153 8810 6205
rect 13078 6153 13130 6205
rect 5494 6079 5546 6131
rect 6262 6079 6314 6131
rect 9238 6079 9290 6131
rect 14902 6153 14954 6205
rect 13270 6079 13322 6131
rect 14518 6079 14570 6131
rect 14710 6079 14762 6131
rect 20470 6227 20522 6279
rect 20566 6227 20618 6279
rect 22774 6227 22826 6279
rect 22966 6270 23018 6279
rect 22966 6236 22975 6270
rect 22975 6236 23009 6270
rect 23009 6236 23018 6270
rect 22966 6227 23018 6236
rect 24406 6227 24458 6279
rect 25654 6310 25663 6344
rect 25663 6310 25697 6344
rect 25697 6310 25706 6344
rect 25654 6301 25706 6310
rect 26806 6344 26858 6353
rect 26806 6310 26815 6344
rect 26815 6310 26849 6344
rect 26849 6310 26858 6344
rect 26806 6301 26858 6310
rect 29686 6344 29738 6353
rect 29686 6310 29695 6344
rect 29695 6310 29729 6344
rect 29729 6310 29738 6344
rect 29686 6301 29738 6310
rect 31222 6344 31274 6353
rect 31222 6310 31231 6344
rect 31231 6310 31265 6344
rect 31265 6310 31274 6344
rect 31222 6301 31274 6310
rect 32086 6418 32138 6427
rect 32086 6384 32095 6418
rect 32095 6384 32129 6418
rect 32129 6384 32138 6418
rect 32086 6375 32138 6384
rect 34294 6418 34346 6427
rect 34294 6384 34303 6418
rect 34303 6384 34337 6418
rect 34337 6384 34346 6418
rect 34294 6375 34346 6384
rect 34678 6418 34730 6427
rect 34678 6384 34687 6418
rect 34687 6384 34721 6418
rect 34721 6384 34730 6418
rect 38518 6523 38570 6575
rect 41206 6523 41258 6575
rect 37270 6449 37322 6501
rect 43222 6523 43274 6575
rect 44566 6566 44618 6575
rect 44566 6532 44575 6566
rect 44575 6532 44609 6566
rect 44609 6532 44618 6566
rect 44566 6523 44618 6532
rect 42262 6449 42314 6501
rect 46582 6523 46634 6575
rect 51286 6566 51338 6575
rect 51286 6532 51295 6566
rect 51295 6532 51329 6566
rect 51329 6532 51338 6566
rect 51286 6523 51338 6532
rect 44950 6449 45002 6501
rect 34678 6375 34730 6384
rect 36310 6344 36362 6353
rect 17494 6079 17546 6131
rect 18454 6079 18506 6131
rect 19510 6079 19562 6131
rect 21430 6122 21482 6131
rect 21430 6088 21439 6122
rect 21439 6088 21473 6122
rect 21473 6088 21482 6122
rect 21430 6079 21482 6088
rect 21526 6079 21578 6131
rect 22966 6079 23018 6131
rect 24310 6079 24362 6131
rect 27574 6079 27626 6131
rect 28438 6079 28490 6131
rect 33142 6153 33194 6205
rect 29782 6079 29834 6131
rect 30646 6079 30698 6131
rect 33334 6153 33386 6205
rect 34486 6153 34538 6205
rect 35926 6153 35978 6205
rect 36310 6310 36319 6344
rect 36319 6310 36353 6344
rect 36353 6310 36362 6344
rect 36310 6301 36362 6310
rect 39478 6375 39530 6427
rect 41302 6418 41354 6427
rect 41302 6384 41311 6418
rect 41311 6384 41345 6418
rect 41345 6384 41354 6418
rect 41302 6375 41354 6384
rect 38902 6344 38954 6353
rect 38902 6310 38911 6344
rect 38911 6310 38945 6344
rect 38945 6310 38954 6344
rect 38902 6301 38954 6310
rect 40342 6344 40394 6353
rect 40342 6310 40351 6344
rect 40351 6310 40385 6344
rect 40385 6310 40394 6344
rect 40342 6301 40394 6310
rect 42646 6375 42698 6427
rect 44182 6375 44234 6427
rect 44566 6375 44618 6427
rect 41878 6344 41930 6353
rect 41878 6310 41887 6344
rect 41887 6310 41921 6344
rect 41921 6310 41930 6344
rect 41878 6301 41930 6310
rect 50422 6375 50474 6427
rect 52246 6375 52298 6427
rect 45526 6344 45578 6353
rect 40630 6227 40682 6279
rect 41302 6227 41354 6279
rect 41494 6227 41546 6279
rect 45526 6310 45535 6344
rect 45535 6310 45569 6344
rect 45569 6310 45578 6344
rect 45526 6301 45578 6310
rect 46966 6344 47018 6353
rect 46966 6310 46975 6344
rect 46975 6310 47009 6344
rect 47009 6310 47018 6344
rect 46966 6301 47018 6310
rect 47734 6344 47786 6353
rect 47734 6310 47743 6344
rect 47743 6310 47777 6344
rect 47777 6310 47786 6344
rect 47734 6301 47786 6310
rect 48790 6301 48842 6353
rect 49558 6301 49610 6353
rect 56374 6375 56426 6427
rect 53974 6301 54026 6353
rect 42358 6227 42410 6279
rect 43702 6270 43754 6279
rect 43702 6236 43711 6270
rect 43711 6236 43745 6270
rect 43745 6236 43754 6270
rect 43702 6227 43754 6236
rect 33430 6079 33482 6131
rect 33718 6079 33770 6131
rect 34294 6079 34346 6131
rect 35446 6079 35498 6131
rect 46582 6153 46634 6205
rect 52246 6227 52298 6279
rect 54358 6227 54410 6279
rect 51574 6153 51626 6205
rect 39190 6079 39242 6131
rect 41302 6079 41354 6131
rect 43990 6079 44042 6131
rect 49846 6079 49898 6131
rect 51094 6079 51146 6131
rect 55126 6153 55178 6205
rect 58102 6301 58154 6353
rect 58870 6227 58922 6279
rect 19654 5968 19706 6020
rect 19718 5968 19770 6020
rect 19782 5968 19834 6020
rect 19846 5968 19898 6020
rect 50374 5968 50426 6020
rect 50438 5968 50490 6020
rect 50502 5968 50554 6020
rect 50566 5968 50618 6020
rect 5206 5857 5258 5909
rect 42742 5857 42794 5909
rect 43318 5857 43370 5909
rect 47158 5857 47210 5909
rect 55030 5900 55082 5909
rect 55030 5866 55039 5900
rect 55039 5866 55073 5900
rect 55073 5866 55082 5900
rect 55030 5857 55082 5866
rect 7606 5783 7658 5835
rect 12022 5709 12074 5761
rect 14230 5709 14282 5761
rect 1078 5635 1130 5687
rect 2902 5678 2954 5687
rect 2902 5644 2911 5678
rect 2911 5644 2945 5678
rect 2945 5644 2954 5678
rect 2902 5635 2954 5644
rect 4918 5635 4970 5687
rect 5206 5678 5258 5687
rect 5206 5644 5215 5678
rect 5215 5644 5249 5678
rect 5249 5644 5258 5678
rect 5206 5635 5258 5644
rect 6838 5678 6890 5687
rect 6838 5644 6847 5678
rect 6847 5644 6881 5678
rect 6881 5644 6890 5678
rect 6838 5635 6890 5644
rect 7222 5635 7274 5687
rect 5782 5561 5834 5613
rect 7606 5487 7658 5539
rect 8758 5635 8810 5687
rect 10198 5635 10250 5687
rect 10486 5635 10538 5687
rect 12598 5678 12650 5687
rect 12598 5644 12607 5678
rect 12607 5644 12641 5678
rect 12641 5644 12650 5678
rect 12598 5635 12650 5644
rect 13366 5678 13418 5687
rect 13366 5644 13375 5678
rect 13375 5644 13409 5678
rect 13409 5644 13418 5678
rect 13366 5635 13418 5644
rect 10582 5561 10634 5613
rect 20566 5783 20618 5835
rect 22870 5709 22922 5761
rect 33142 5783 33194 5835
rect 23542 5709 23594 5761
rect 29878 5709 29930 5761
rect 32950 5709 33002 5761
rect 37750 5783 37802 5835
rect 35926 5709 35978 5761
rect 41974 5709 42026 5761
rect 14998 5678 15050 5687
rect 14998 5644 15007 5678
rect 15007 5644 15041 5678
rect 15041 5644 15050 5678
rect 14998 5635 15050 5644
rect 15862 5678 15914 5687
rect 15862 5644 15871 5678
rect 15871 5644 15905 5678
rect 15905 5644 15914 5678
rect 15862 5635 15914 5644
rect 16150 5635 16202 5687
rect 17398 5678 17450 5687
rect 17398 5644 17407 5678
rect 17407 5644 17441 5678
rect 17441 5644 17450 5678
rect 17398 5635 17450 5644
rect 18742 5678 18794 5687
rect 18742 5644 18751 5678
rect 18751 5644 18785 5678
rect 18785 5644 18794 5678
rect 18742 5635 18794 5644
rect 20182 5678 20234 5687
rect 20182 5644 20191 5678
rect 20191 5644 20225 5678
rect 20225 5644 20234 5678
rect 20182 5635 20234 5644
rect 20566 5635 20618 5687
rect 21718 5678 21770 5687
rect 21718 5644 21727 5678
rect 21727 5644 21761 5678
rect 21761 5644 21770 5678
rect 21718 5635 21770 5644
rect 21622 5561 21674 5613
rect 23062 5635 23114 5687
rect 23446 5635 23498 5687
rect 24598 5635 24650 5687
rect 26230 5678 26282 5687
rect 26230 5644 26239 5678
rect 26239 5644 26273 5678
rect 26273 5644 26282 5678
rect 26230 5635 26282 5644
rect 26038 5561 26090 5613
rect 27382 5635 27434 5687
rect 27862 5635 27914 5687
rect 28822 5635 28874 5687
rect 30262 5635 30314 5687
rect 30838 5635 30890 5687
rect 31702 5635 31754 5687
rect 33142 5678 33194 5687
rect 33142 5644 33151 5678
rect 33151 5644 33185 5678
rect 33185 5644 33194 5678
rect 33142 5635 33194 5644
rect 34678 5678 34730 5687
rect 33238 5561 33290 5613
rect 34678 5644 34687 5678
rect 34687 5644 34721 5678
rect 34721 5644 34730 5678
rect 34678 5635 34730 5644
rect 36022 5678 36074 5687
rect 36022 5644 36031 5678
rect 36031 5644 36065 5678
rect 36065 5644 36074 5678
rect 36022 5635 36074 5644
rect 36214 5635 36266 5687
rect 37558 5678 37610 5687
rect 37558 5644 37567 5678
rect 37567 5644 37601 5678
rect 37601 5644 37610 5678
rect 37558 5635 37610 5644
rect 39094 5678 39146 5687
rect 37462 5561 37514 5613
rect 39094 5644 39103 5678
rect 39103 5644 39137 5678
rect 39137 5644 39146 5678
rect 39094 5635 39146 5644
rect 39286 5635 39338 5687
rect 40726 5635 40778 5687
rect 41782 5635 41834 5687
rect 42262 5635 42314 5687
rect 43222 5635 43274 5687
rect 43702 5635 43754 5687
rect 45142 5678 45194 5687
rect 45142 5644 45151 5678
rect 45151 5644 45185 5678
rect 45185 5644 45194 5678
rect 45142 5635 45194 5644
rect 46102 5635 46154 5687
rect 46678 5635 46730 5687
rect 47542 5635 47594 5687
rect 48982 5678 49034 5687
rect 48982 5644 48991 5678
rect 48991 5644 49025 5678
rect 49025 5644 49034 5678
rect 48982 5635 49034 5644
rect 49654 5678 49706 5687
rect 49654 5644 49663 5678
rect 49663 5644 49697 5678
rect 49697 5644 49706 5678
rect 49654 5635 49706 5644
rect 50710 5635 50762 5687
rect 52150 5678 52202 5687
rect 52150 5644 52159 5678
rect 52159 5644 52193 5678
rect 52193 5644 52202 5678
rect 52150 5635 52202 5644
rect 52534 5635 52586 5687
rect 53686 5678 53738 5687
rect 53686 5644 53695 5678
rect 53695 5644 53729 5678
rect 53729 5644 53738 5678
rect 53686 5635 53738 5644
rect 57430 5678 57482 5687
rect 42742 5561 42794 5613
rect 43318 5561 43370 5613
rect 53590 5561 53642 5613
rect 57430 5644 57439 5678
rect 57439 5644 57473 5678
rect 57473 5644 57482 5678
rect 57430 5635 57482 5644
rect 59638 5561 59690 5613
rect 20470 5487 20522 5539
rect 29110 5487 29162 5539
rect 7126 5413 7178 5465
rect 11542 5413 11594 5465
rect 47638 5413 47690 5465
rect 4294 5302 4346 5354
rect 4358 5302 4410 5354
rect 4422 5302 4474 5354
rect 4486 5302 4538 5354
rect 35014 5302 35066 5354
rect 35078 5302 35130 5354
rect 35142 5302 35194 5354
rect 35206 5302 35258 5354
rect 4726 5191 4778 5243
rect 1846 5117 1898 5169
rect 3574 5117 3626 5169
rect 310 4969 362 5021
rect 1846 4969 1898 5021
rect 3094 5012 3146 5021
rect 3094 4978 3103 5012
rect 3103 4978 3137 5012
rect 3137 4978 3146 5012
rect 3094 4969 3146 4978
rect 4150 5012 4202 5021
rect 4150 4978 4159 5012
rect 4159 4978 4193 5012
rect 4193 4978 4202 5012
rect 4150 4969 4202 4978
rect 5398 5012 5450 5021
rect 5398 4978 5407 5012
rect 5407 4978 5441 5012
rect 5441 4978 5450 5012
rect 5398 4969 5450 4978
rect 6070 4969 6122 5021
rect 9238 5012 9290 5021
rect 9238 4978 9247 5012
rect 9247 4978 9281 5012
rect 9281 4978 9290 5012
rect 9238 4969 9290 4978
rect 10582 4969 10634 5021
rect 10966 4969 11018 5021
rect 11830 4969 11882 5021
rect 13942 5012 13994 5021
rect 12214 4821 12266 4873
rect 13942 4978 13951 5012
rect 13951 4978 13985 5012
rect 13985 4978 13994 5012
rect 13942 4969 13994 4978
rect 14422 4969 14474 5021
rect 14806 4969 14858 5021
rect 16438 4969 16490 5021
rect 17302 4969 17354 5021
rect 17974 4969 18026 5021
rect 19030 5012 19082 5021
rect 19030 4978 19039 5012
rect 19039 4978 19073 5012
rect 19073 4978 19082 5012
rect 19030 4969 19082 4978
rect 19126 4969 19178 5021
rect 20470 4969 20522 5021
rect 20950 4969 21002 5021
rect 22102 4969 22154 5021
rect 23542 5012 23594 5021
rect 23542 4978 23551 5012
rect 23551 4978 23585 5012
rect 23585 4978 23594 5012
rect 23542 4969 23594 4978
rect 25078 5012 25130 5021
rect 23158 4895 23210 4947
rect 25078 4978 25087 5012
rect 25087 4978 25121 5012
rect 25121 4978 25130 5012
rect 25078 4969 25130 4978
rect 25846 5012 25898 5021
rect 25846 4978 25855 5012
rect 25855 4978 25889 5012
rect 25889 4978 25898 5012
rect 25846 4969 25898 4978
rect 26614 5012 26666 5021
rect 26614 4978 26623 5012
rect 26623 4978 26657 5012
rect 26657 4978 26666 5012
rect 26614 4969 26666 4978
rect 28054 5012 28106 5021
rect 28054 4978 28063 5012
rect 28063 4978 28097 5012
rect 28097 4978 28106 5012
rect 28054 4969 28106 4978
rect 28918 5012 28970 5021
rect 28918 4978 28927 5012
rect 28927 4978 28961 5012
rect 28961 4978 28970 5012
rect 28918 4969 28970 4978
rect 29014 4969 29066 5021
rect 30358 5012 30410 5021
rect 30358 4978 30367 5012
rect 30367 4978 30401 5012
rect 30401 4978 30410 5012
rect 30358 4969 30410 4978
rect 30454 4969 30506 5021
rect 31894 5012 31946 5021
rect 31894 4978 31903 5012
rect 31903 4978 31937 5012
rect 31937 4978 31946 5012
rect 31894 4969 31946 4978
rect 33334 5012 33386 5021
rect 33334 4978 33343 5012
rect 33343 4978 33377 5012
rect 33377 4978 33386 5012
rect 33334 4969 33386 4978
rect 34102 5012 34154 5021
rect 34102 4978 34111 5012
rect 34111 4978 34145 5012
rect 34145 4978 34154 5012
rect 34102 4969 34154 4978
rect 34774 4969 34826 5021
rect 34582 4895 34634 4947
rect 36502 4969 36554 5021
rect 38614 5012 38666 5021
rect 38614 4978 38623 5012
rect 38623 4978 38657 5012
rect 38657 4978 38666 5012
rect 38614 4969 38666 4978
rect 39382 5012 39434 5021
rect 39382 4978 39391 5012
rect 39391 4978 39425 5012
rect 39425 4978 39434 5012
rect 39382 4969 39434 4978
rect 40150 5012 40202 5021
rect 40150 4978 40159 5012
rect 40159 4978 40193 5012
rect 40193 4978 40202 5012
rect 40150 4969 40202 4978
rect 40918 5012 40970 5021
rect 40918 4978 40927 5012
rect 40927 4978 40961 5012
rect 40961 4978 40970 5012
rect 40918 4969 40970 4978
rect 41014 4969 41066 5021
rect 42070 4969 42122 5021
rect 43510 4969 43562 5021
rect 44758 5012 44810 5021
rect 44758 4978 44767 5012
rect 44767 4978 44801 5012
rect 44801 4978 44810 5012
rect 44758 4969 44810 4978
rect 45430 5012 45482 5021
rect 45430 4978 45439 5012
rect 45439 4978 45473 5012
rect 45473 4978 45482 5012
rect 45430 4969 45482 4978
rect 46198 5012 46250 5021
rect 46198 4978 46207 5012
rect 46207 4978 46241 5012
rect 46241 4978 46250 5012
rect 46198 4969 46250 4978
rect 46390 4969 46442 5021
rect 47638 4969 47690 5021
rect 49366 5012 49418 5021
rect 49366 4978 49375 5012
rect 49375 4978 49409 5012
rect 49409 4978 49418 5012
rect 49366 4969 49418 4978
rect 50422 5012 50474 5021
rect 50422 4978 50431 5012
rect 50431 4978 50465 5012
rect 50465 4978 50474 5012
rect 50422 4969 50474 4978
rect 50902 4969 50954 5021
rect 51862 5012 51914 5021
rect 51862 4978 51871 5012
rect 51871 4978 51905 5012
rect 51905 4978 51914 5012
rect 51862 4969 51914 4978
rect 51958 4969 52010 5021
rect 53302 4969 53354 5021
rect 57046 5012 57098 5021
rect 36886 4895 36938 4947
rect 57046 4978 57055 5012
rect 57055 4978 57089 5012
rect 57089 4978 57098 5012
rect 57046 4969 57098 4978
rect 57814 4895 57866 4947
rect 59254 4821 59306 4873
rect 8854 4747 8906 4799
rect 9910 4747 9962 4799
rect 39958 4747 40010 4799
rect 19654 4636 19706 4688
rect 19718 4636 19770 4688
rect 19782 4636 19834 4688
rect 19846 4636 19898 4688
rect 50374 4636 50426 4688
rect 50438 4636 50490 4688
rect 50502 4636 50554 4688
rect 50566 4636 50618 4688
rect 7414 4525 7466 4577
rect 43798 4525 43850 4577
rect 8086 4451 8138 4503
rect 8950 4451 9002 4503
rect 10774 4451 10826 4503
rect 11446 4451 11498 4503
rect 11542 4451 11594 4503
rect 790 4377 842 4429
rect 1174 4303 1226 4355
rect 8278 4377 8330 4429
rect 32950 4451 33002 4503
rect 33910 4451 33962 4503
rect 17590 4377 17642 4429
rect 1366 4229 1418 4281
rect 3766 4229 3818 4281
rect 4726 4303 4778 4355
rect 3478 4155 3530 4207
rect 4918 4155 4970 4207
rect 5110 4155 5162 4207
rect 7414 4346 7466 4355
rect 5686 4229 5738 4281
rect 7414 4312 7423 4346
rect 7423 4312 7457 4346
rect 7457 4312 7466 4346
rect 7414 4303 7466 4312
rect 6454 4155 6506 4207
rect 9622 4346 9674 4355
rect 9622 4312 9631 4346
rect 9631 4312 9665 4346
rect 9665 4312 9674 4346
rect 9622 4303 9674 4312
rect 10390 4346 10442 4355
rect 10390 4312 10399 4346
rect 10399 4312 10433 4346
rect 10433 4312 10442 4346
rect 10390 4303 10442 4312
rect 10774 4303 10826 4355
rect 7894 4229 7946 4281
rect 9814 4229 9866 4281
rect 9334 4155 9386 4207
rect 982 4081 1034 4133
rect 2326 4081 2378 4133
rect 2422 4081 2474 4133
rect 5014 4081 5066 4133
rect 9046 4081 9098 4133
rect 10966 4081 11018 4133
rect 11158 4155 11210 4207
rect 13558 4346 13610 4355
rect 11446 4229 11498 4281
rect 13558 4312 13567 4346
rect 13567 4312 13601 4346
rect 13601 4312 13610 4346
rect 13558 4303 13610 4312
rect 15478 4346 15530 4355
rect 15478 4312 15487 4346
rect 15487 4312 15521 4346
rect 15521 4312 15530 4346
rect 15478 4303 15530 4312
rect 15958 4303 16010 4355
rect 24406 4377 24458 4429
rect 56758 4451 56810 4503
rect 57334 4451 57386 4503
rect 20278 4346 20330 4355
rect 13846 4229 13898 4281
rect 14518 4229 14570 4281
rect 11926 4081 11978 4133
rect 13078 4081 13130 4133
rect 14134 4155 14186 4207
rect 14710 4155 14762 4207
rect 16246 4155 16298 4207
rect 16822 4081 16874 4133
rect 16918 4081 16970 4133
rect 20278 4312 20287 4346
rect 20287 4312 20321 4346
rect 20321 4312 20330 4346
rect 20278 4303 20330 4312
rect 21046 4346 21098 4355
rect 21046 4312 21055 4346
rect 21055 4312 21089 4346
rect 21089 4312 21098 4346
rect 21046 4303 21098 4312
rect 21814 4346 21866 4355
rect 21814 4312 21823 4346
rect 21823 4312 21857 4346
rect 21857 4312 21866 4346
rect 21814 4303 21866 4312
rect 23254 4346 23306 4355
rect 23254 4312 23263 4346
rect 23263 4312 23297 4346
rect 23297 4312 23306 4346
rect 23254 4303 23306 4312
rect 24022 4346 24074 4355
rect 24022 4312 24031 4346
rect 24031 4312 24065 4346
rect 24065 4312 24074 4346
rect 24022 4303 24074 4312
rect 25462 4346 25514 4355
rect 25462 4312 25471 4346
rect 25471 4312 25505 4346
rect 25505 4312 25514 4346
rect 25462 4303 25514 4312
rect 21238 4229 21290 4281
rect 22006 4229 22058 4281
rect 22774 4272 22826 4281
rect 22774 4238 22783 4272
rect 22783 4238 22817 4272
rect 22817 4238 22826 4272
rect 22774 4229 22826 4238
rect 24214 4229 24266 4281
rect 25846 4229 25898 4281
rect 26134 4303 26186 4355
rect 26518 4303 26570 4355
rect 28342 4346 28394 4355
rect 28342 4312 28351 4346
rect 28351 4312 28385 4346
rect 28385 4312 28394 4346
rect 28342 4303 28394 4312
rect 29110 4346 29162 4355
rect 29110 4312 29119 4346
rect 29119 4312 29153 4346
rect 29153 4312 29162 4346
rect 29110 4303 29162 4312
rect 30934 4346 30986 4355
rect 30934 4312 30943 4346
rect 30943 4312 30977 4346
rect 30977 4312 30986 4346
rect 30934 4303 30986 4312
rect 22294 4155 22346 4207
rect 22966 4155 23018 4207
rect 25366 4155 25418 4207
rect 26230 4155 26282 4207
rect 31702 4346 31754 4355
rect 31702 4312 31711 4346
rect 31711 4312 31745 4346
rect 31745 4312 31754 4346
rect 31702 4303 31754 4312
rect 32758 4346 32810 4355
rect 32758 4312 32767 4346
rect 32767 4312 32801 4346
rect 32801 4312 32810 4346
rect 32758 4303 32810 4312
rect 33910 4346 33962 4355
rect 33910 4312 33919 4346
rect 33919 4312 33953 4346
rect 33953 4312 33962 4346
rect 33910 4303 33962 4312
rect 34582 4303 34634 4355
rect 31414 4155 31466 4207
rect 32374 4155 32426 4207
rect 34198 4229 34250 4281
rect 36790 4346 36842 4355
rect 36790 4312 36799 4346
rect 36799 4312 36833 4346
rect 36833 4312 36842 4346
rect 36790 4303 36842 4312
rect 38998 4346 39050 4355
rect 37174 4229 37226 4281
rect 38998 4312 39007 4346
rect 39007 4312 39041 4346
rect 39041 4312 39050 4346
rect 38998 4303 39050 4312
rect 39766 4346 39818 4355
rect 39766 4312 39775 4346
rect 39775 4312 39809 4346
rect 39809 4312 39818 4346
rect 39766 4303 39818 4312
rect 41974 4346 42026 4355
rect 41974 4312 41983 4346
rect 41983 4312 42017 4346
rect 42017 4312 42026 4346
rect 41974 4303 42026 4312
rect 42358 4303 42410 4355
rect 43414 4303 43466 4355
rect 44950 4346 45002 4355
rect 44950 4312 44959 4346
rect 44959 4312 44993 4346
rect 44993 4312 45002 4346
rect 44950 4303 45002 4312
rect 46774 4346 46826 4355
rect 46774 4312 46783 4346
rect 46783 4312 46817 4346
rect 46817 4312 46826 4346
rect 46774 4303 46826 4312
rect 38134 4229 38186 4281
rect 39094 4229 39146 4281
rect 41494 4229 41546 4281
rect 41782 4229 41834 4281
rect 43606 4229 43658 4281
rect 44374 4229 44426 4281
rect 44470 4229 44522 4281
rect 45142 4229 45194 4281
rect 47446 4229 47498 4281
rect 47830 4303 47882 4355
rect 48598 4229 48650 4281
rect 49174 4303 49226 4355
rect 52630 4346 52682 4355
rect 49942 4229 49994 4281
rect 50998 4229 51050 4281
rect 52630 4312 52639 4346
rect 52639 4312 52673 4346
rect 52673 4312 52682 4346
rect 52630 4303 52682 4312
rect 53014 4229 53066 4281
rect 54070 4303 54122 4355
rect 55606 4346 55658 4355
rect 55606 4312 55615 4346
rect 55615 4312 55649 4346
rect 55649 4312 55658 4346
rect 55606 4303 55658 4312
rect 57334 4303 57386 4355
rect 56566 4229 56618 4281
rect 58294 4229 58346 4281
rect 55990 4155 56042 4207
rect 57910 4155 57962 4207
rect 25558 4081 25610 4133
rect 25942 4081 25994 4133
rect 26422 4081 26474 4133
rect 28054 4081 28106 4133
rect 28246 4081 28298 4133
rect 29014 4081 29066 4133
rect 29302 4081 29354 4133
rect 30454 4081 30506 4133
rect 31798 4081 31850 4133
rect 33046 4081 33098 4133
rect 33814 4081 33866 4133
rect 34678 4081 34730 4133
rect 38518 4081 38570 4133
rect 40150 4081 40202 4133
rect 48118 4081 48170 4133
rect 48982 4081 49034 4133
rect 49270 4081 49322 4133
rect 50710 4081 50762 4133
rect 4294 3970 4346 4022
rect 4358 3970 4410 4022
rect 4422 3970 4474 4022
rect 4486 3970 4538 4022
rect 35014 3970 35066 4022
rect 35078 3970 35130 4022
rect 35142 3970 35194 4022
rect 35206 3970 35258 4022
rect 1942 3859 1994 3911
rect 2998 3859 3050 3911
rect 7894 3859 7946 3911
rect 9238 3859 9290 3911
rect 9814 3859 9866 3911
rect 502 3785 554 3837
rect 1654 3785 1706 3837
rect 2326 3785 2378 3837
rect 3094 3785 3146 3837
rect 8278 3785 8330 3837
rect 10582 3785 10634 3837
rect 11542 3859 11594 3911
rect 16534 3859 16586 3911
rect 17398 3859 17450 3911
rect 18358 3859 18410 3911
rect 19030 3859 19082 3911
rect 19222 3859 19274 3911
rect 19414 3859 19466 3911
rect 20470 3859 20522 3911
rect 21334 3859 21386 3911
rect 22102 3859 22154 3911
rect 23830 3859 23882 3911
rect 25078 3859 25130 3911
rect 25942 3859 25994 3911
rect 26902 3859 26954 3911
rect 27478 3859 27530 3911
rect 28918 3859 28970 3911
rect 29014 3859 29066 3911
rect 30358 3859 30410 3911
rect 30742 3859 30794 3911
rect 31990 3859 32042 3911
rect 33430 3859 33482 3911
rect 34774 3859 34826 3911
rect 37078 3859 37130 3911
rect 38614 3859 38666 3911
rect 39670 3859 39722 3911
rect 40918 3859 40970 3911
rect 41110 3859 41162 3911
rect 42070 3859 42122 3911
rect 43318 3859 43370 3911
rect 44758 3859 44810 3911
rect 44854 3859 44906 3911
rect 46198 3859 46250 3911
rect 46294 3859 46346 3911
rect 47638 3859 47690 3911
rect 48502 3859 48554 3911
rect 49654 3859 49706 3911
rect 51382 3859 51434 3911
rect 51862 3859 51914 3911
rect 56278 3859 56330 3911
rect 2998 3711 3050 3763
rect 3286 3711 3338 3763
rect 3382 3711 3434 3763
rect 118 3637 170 3689
rect 1654 3637 1706 3689
rect 2710 3637 2762 3689
rect 18934 3785 18986 3837
rect 5590 3680 5642 3689
rect 214 3563 266 3615
rect 1750 3563 1802 3615
rect 598 3489 650 3541
rect 1462 3489 1514 3541
rect 3094 3489 3146 3541
rect 5590 3646 5599 3680
rect 5599 3646 5633 3680
rect 5633 3646 5642 3680
rect 5590 3637 5642 3646
rect 6358 3637 6410 3689
rect 7030 3637 7082 3689
rect 7798 3637 7850 3689
rect 8566 3637 8618 3689
rect 9334 3637 9386 3689
rect 7990 3563 8042 3615
rect 20470 3711 20522 3763
rect 20854 3711 20906 3763
rect 25174 3711 25226 3763
rect 26326 3711 26378 3763
rect 27382 3711 27434 3763
rect 28438 3711 28490 3763
rect 28726 3711 28778 3763
rect 34678 3785 34730 3837
rect 35446 3785 35498 3837
rect 35638 3785 35690 3837
rect 36502 3785 36554 3837
rect 37846 3785 37898 3837
rect 39382 3785 39434 3837
rect 39958 3785 40010 3837
rect 41014 3785 41066 3837
rect 44086 3785 44138 3837
rect 45430 3785 45482 3837
rect 56758 3785 56810 3837
rect 59446 3785 59498 3837
rect 10582 3637 10634 3689
rect 13174 3637 13226 3689
rect 13654 3680 13706 3689
rect 13654 3646 13663 3680
rect 13663 3646 13697 3680
rect 13697 3646 13706 3680
rect 13654 3637 13706 3646
rect 14038 3637 14090 3689
rect 14806 3637 14858 3689
rect 15286 3637 15338 3689
rect 17398 3637 17450 3689
rect 18070 3637 18122 3689
rect 18454 3637 18506 3689
rect 19222 3637 19274 3689
rect 19990 3637 20042 3689
rect 20662 3637 20714 3689
rect 22102 3637 22154 3689
rect 22870 3637 22922 3689
rect 23638 3637 23690 3689
rect 24406 3637 24458 3689
rect 10006 3489 10058 3541
rect 10582 3489 10634 3541
rect 24694 3563 24746 3615
rect 19030 3489 19082 3541
rect 19510 3489 19562 3541
rect 25846 3489 25898 3541
rect 27286 3637 27338 3689
rect 36694 3711 36746 3763
rect 41302 3711 41354 3763
rect 41590 3711 41642 3763
rect 45238 3711 45290 3763
rect 28054 3489 28106 3541
rect 29494 3563 29546 3615
rect 30454 3637 30506 3689
rect 31318 3637 31370 3689
rect 32470 3637 32522 3689
rect 33526 3637 33578 3689
rect 34294 3637 34346 3689
rect 35350 3637 35402 3689
rect 35734 3637 35786 3689
rect 36502 3637 36554 3689
rect 37942 3637 37994 3689
rect 38710 3637 38762 3689
rect 39478 3637 39530 3689
rect 40246 3637 40298 3689
rect 41014 3637 41066 3689
rect 36694 3563 36746 3615
rect 37558 3563 37610 3615
rect 41590 3563 41642 3615
rect 42742 3637 42794 3689
rect 47542 3711 47594 3763
rect 48310 3711 48362 3763
rect 55894 3711 55946 3763
rect 43798 3563 43850 3615
rect 30454 3489 30506 3541
rect 31894 3489 31946 3541
rect 44566 3489 44618 3541
rect 46006 3563 46058 3615
rect 47158 3637 47210 3689
rect 48214 3637 48266 3689
rect 50710 3637 50762 3689
rect 50806 3637 50858 3689
rect 51286 3637 51338 3689
rect 52054 3637 52106 3689
rect 53398 3637 53450 3689
rect 59158 3711 59210 3763
rect 45718 3489 45770 3541
rect 46390 3489 46442 3541
rect 49078 3489 49130 3541
rect 50038 3489 50090 3541
rect 51286 3489 51338 3541
rect 51478 3489 51530 3541
rect 52054 3489 52106 3541
rect 52726 3489 52778 3541
rect 54454 3489 54506 3541
rect 3286 3415 3338 3467
rect 3958 3415 4010 3467
rect 7510 3415 7562 3467
rect 11926 3415 11978 3467
rect 12022 3415 12074 3467
rect 13366 3415 13418 3467
rect 14230 3415 14282 3467
rect 20854 3458 20906 3467
rect 20854 3424 20863 3458
rect 20863 3424 20897 3458
rect 20897 3424 20906 3458
rect 20854 3415 20906 3424
rect 26326 3415 26378 3467
rect 27574 3415 27626 3467
rect 28918 3415 28970 3467
rect 29782 3415 29834 3467
rect 32566 3415 32618 3467
rect 33718 3415 33770 3467
rect 45430 3415 45482 3467
rect 45622 3415 45674 3467
rect 55222 3415 55274 3467
rect 56566 3563 56618 3615
rect 56854 3563 56906 3615
rect 56278 3489 56330 3541
rect 58198 3637 58250 3689
rect 59734 3637 59786 3689
rect 19654 3304 19706 3356
rect 19718 3304 19770 3356
rect 19782 3304 19834 3356
rect 19846 3304 19898 3356
rect 50374 3304 50426 3356
rect 50438 3304 50490 3356
rect 50502 3304 50554 3356
rect 50566 3304 50618 3356
rect 1462 3193 1514 3245
rect 2134 3193 2186 3245
rect 3958 3193 4010 3245
rect 5206 3193 5258 3245
rect 8182 3193 8234 3245
rect 7126 3119 7178 3171
rect 13078 3119 13130 3171
rect 13750 3193 13802 3245
rect 16822 3236 16874 3245
rect 16822 3202 16831 3236
rect 16831 3202 16865 3236
rect 16865 3202 16874 3236
rect 16822 3193 16874 3202
rect 18934 3193 18986 3245
rect 19702 3193 19754 3245
rect 20374 3193 20426 3245
rect 20950 3193 21002 3245
rect 21718 3193 21770 3245
rect 22006 3193 22058 3245
rect 24022 3193 24074 3245
rect 24982 3193 25034 3245
rect 26614 3193 26666 3245
rect 32662 3193 32714 3245
rect 34102 3193 34154 3245
rect 40054 3193 40106 3245
rect 40246 3193 40298 3245
rect 41206 3193 41258 3245
rect 56374 3193 56426 3245
rect 58006 3193 58058 3245
rect 8950 3045 9002 3097
rect 22 2971 74 3023
rect 694 2897 746 2949
rect 2134 2897 2186 2949
rect 4918 3014 4970 3023
rect 4918 2980 4927 3014
rect 4927 2980 4961 3014
rect 4961 2980 4970 3014
rect 4918 2971 4970 2980
rect 5206 2971 5258 3023
rect 5974 2971 6026 3023
rect 5110 2749 5162 2801
rect 5782 2897 5834 2949
rect 6742 2897 6794 2949
rect 8182 2971 8234 3023
rect 8950 2897 9002 2949
rect 19798 3119 19850 3171
rect 20182 3119 20234 3171
rect 21142 3119 21194 3171
rect 21430 3119 21482 3171
rect 22966 3119 23018 3171
rect 24310 3119 24362 3171
rect 40822 3119 40874 3171
rect 42070 3119 42122 3171
rect 44182 3119 44234 3171
rect 15382 3045 15434 3097
rect 16438 3045 16490 3097
rect 19510 3045 19562 3097
rect 22390 3045 22442 3097
rect 23542 3045 23594 3097
rect 31894 3045 31946 3097
rect 33334 3045 33386 3097
rect 42550 3045 42602 3097
rect 43510 3045 43562 3097
rect 46390 3045 46442 3097
rect 12982 3014 13034 3023
rect 12982 2980 12991 3014
rect 12991 2980 13025 3014
rect 13025 2980 13034 3014
rect 12982 2971 13034 2980
rect 13366 2971 13418 3023
rect 14518 2971 14570 3023
rect 16630 3014 16682 3023
rect 16630 2980 16639 3014
rect 16639 2980 16673 3014
rect 16673 2980 16682 3014
rect 16630 2971 16682 2980
rect 17014 2971 17066 3023
rect 14230 2897 14282 2949
rect 17686 2897 17738 2949
rect 18934 2971 18986 3023
rect 19606 2897 19658 2949
rect 21430 2971 21482 3023
rect 21142 2897 21194 2949
rect 22486 2897 22538 2949
rect 24022 2971 24074 3023
rect 25078 2897 25130 2949
rect 26902 2971 26954 3023
rect 27574 2897 27626 2949
rect 29878 2971 29930 3023
rect 30550 2897 30602 2949
rect 32086 2971 32138 3023
rect 32278 2897 32330 2949
rect 33142 2897 33194 2949
rect 33334 2897 33386 2949
rect 35446 2971 35498 3023
rect 36118 2897 36170 2949
rect 37558 2971 37610 3023
rect 38326 2897 38378 2949
rect 40534 2971 40586 3023
rect 41206 2897 41258 2949
rect 43030 2971 43082 3023
rect 44182 2897 44234 2949
rect 45622 2971 45674 3023
rect 52246 3045 52298 3097
rect 56374 3045 56426 3097
rect 49654 2971 49706 3023
rect 51478 2971 51530 3023
rect 52246 2897 52298 2949
rect 53782 2971 53834 3023
rect 52918 2897 52970 2949
rect 53686 2897 53738 2949
rect 54838 2897 54890 2949
rect 56662 2971 56714 3023
rect 57334 2971 57386 3023
rect 6166 2823 6218 2875
rect 19510 2749 19562 2801
rect 20086 2749 20138 2801
rect 23926 2749 23978 2801
rect 27766 2749 27818 2801
rect 27958 2749 28010 2801
rect 50038 2823 50090 2875
rect 45334 2749 45386 2801
rect 46102 2749 46154 2801
rect 47062 2749 47114 2801
rect 4294 2638 4346 2690
rect 4358 2638 4410 2690
rect 4422 2638 4474 2690
rect 4486 2638 4538 2690
rect 35014 2638 35066 2690
rect 35078 2638 35130 2690
rect 35142 2638 35194 2690
rect 35206 2638 35258 2690
rect 3958 2527 4010 2579
rect 4246 2527 4298 2579
rect 4342 2527 4394 2579
rect 4822 2527 4874 2579
rect 9814 2527 9866 2579
rect 10198 2527 10250 2579
rect 13078 2527 13130 2579
rect 13270 2527 13322 2579
rect 20182 2527 20234 2579
rect 20854 2527 20906 2579
rect 43222 2527 43274 2579
rect 43990 2527 44042 2579
rect 45142 2527 45194 2579
rect 45718 2527 45770 2579
rect 4726 2009 4778 2061
rect 5302 2009 5354 2061
rect 4534 1861 4586 1913
rect 4822 1861 4874 1913
rect 30358 1713 30410 1765
rect 30646 1713 30698 1765
rect 50518 1713 50570 1765
rect 51094 1713 51146 1765
rect 36118 1639 36170 1691
rect 50710 1639 50762 1691
rect 50902 1639 50954 1691
rect 35158 1417 35210 1469
rect 35542 1417 35594 1469
rect 36310 1491 36362 1543
rect 50902 1491 50954 1543
rect 51574 1491 51626 1543
rect 33238 1269 33290 1321
rect 33718 1269 33770 1321
rect 36118 1269 36170 1321
rect 41014 1269 41066 1321
rect 41302 1269 41354 1321
rect 34678 1121 34730 1173
rect 35446 1121 35498 1173
rect 36310 1121 36362 1173
rect 34870 1047 34922 1099
rect 36886 1047 36938 1099
rect 35254 973 35306 1025
rect 35926 973 35978 1025
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 226 56975 254 59200
rect 214 56969 266 56975
rect 214 56911 266 56917
rect 706 56531 734 59200
rect 694 56525 746 56531
rect 694 56467 746 56473
rect 1186 55717 1214 59200
rect 1762 57049 1790 59200
rect 1750 57043 1802 57049
rect 1750 56985 1802 56991
rect 1750 56895 1802 56901
rect 1750 56837 1802 56843
rect 1174 55711 1226 55717
rect 1174 55653 1226 55659
rect 1762 17294 1790 56837
rect 2242 56531 2270 59200
rect 2818 56531 2846 59200
rect 3298 57049 3326 59200
rect 3286 57043 3338 57049
rect 3286 56985 3338 56991
rect 3574 56895 3626 56901
rect 3574 56837 3626 56843
rect 2230 56525 2282 56531
rect 2230 56467 2282 56473
rect 2806 56525 2858 56531
rect 2806 56467 2858 56473
rect 1942 56229 1994 56235
rect 1942 56171 1994 56177
rect 2518 56229 2570 56235
rect 2518 56171 2570 56177
rect 2902 56229 2954 56235
rect 2902 56171 2954 56177
rect 1846 55563 1898 55569
rect 1846 55505 1898 55511
rect 1858 33665 1886 55505
rect 1846 33659 1898 33665
rect 1846 33601 1898 33607
rect 1954 29595 1982 56171
rect 2230 53417 2282 53423
rect 2230 53359 2282 53365
rect 1942 29589 1994 29595
rect 1942 29531 1994 29537
rect 1762 17266 1886 17294
rect 1654 8277 1706 8283
rect 1654 8219 1706 8225
rect 1462 7685 1514 7691
rect 1462 7627 1514 7633
rect 1078 5687 1130 5693
rect 1078 5629 1130 5635
rect 310 5021 362 5027
rect 310 4963 362 4969
rect 118 3689 170 3695
rect 118 3631 170 3637
rect 22 3023 74 3029
rect 22 2965 74 2971
rect 34 800 62 2965
rect 130 800 158 3631
rect 214 3615 266 3621
rect 214 3557 266 3563
rect 226 800 254 3557
rect 322 800 350 4963
rect 790 4429 842 4435
rect 790 4371 842 4377
rect 502 3837 554 3843
rect 502 3779 554 3785
rect 514 800 542 3779
rect 598 3541 650 3547
rect 598 3483 650 3489
rect 610 800 638 3483
rect 694 2949 746 2955
rect 694 2891 746 2897
rect 706 800 734 2891
rect 802 800 830 4371
rect 982 4133 1034 4139
rect 982 4075 1034 4081
rect 994 800 1022 4075
rect 1090 800 1118 5629
rect 1174 4355 1226 4361
rect 1174 4297 1226 4303
rect 1186 800 1214 4297
rect 1366 4281 1418 4287
rect 1366 4223 1418 4229
rect 1378 800 1406 4223
rect 1474 3547 1502 7627
rect 1666 7214 1694 8219
rect 1666 7186 1790 7214
rect 1654 7019 1706 7025
rect 1654 6961 1706 6967
rect 1558 6353 1610 6359
rect 1558 6295 1610 6301
rect 1462 3541 1514 3547
rect 1462 3483 1514 3489
rect 1462 3245 1514 3251
rect 1462 3187 1514 3193
rect 1474 800 1502 3187
rect 1570 800 1598 6295
rect 1666 3843 1694 6961
rect 1654 3837 1706 3843
rect 1654 3779 1706 3785
rect 1654 3689 1706 3695
rect 1654 3631 1706 3637
rect 1666 800 1694 3631
rect 1762 3621 1790 7186
rect 1858 5175 1886 17266
rect 2134 8277 2186 8283
rect 2242 8251 2270 53359
rect 2530 46097 2558 56171
rect 2518 46091 2570 46097
rect 2518 46033 2570 46039
rect 2914 28189 2942 56171
rect 2902 28183 2954 28189
rect 2902 28125 2954 28131
rect 3286 13457 3338 13463
rect 3286 13399 3338 13405
rect 3298 8431 3326 13399
rect 3382 9683 3434 9689
rect 3382 9625 3434 9631
rect 3286 8425 3338 8431
rect 3286 8367 3338 8373
rect 3286 8277 3338 8283
rect 2134 8219 2186 8225
rect 2228 8242 2284 8251
rect 2038 6353 2090 6359
rect 2038 6295 2090 6301
rect 1846 5169 1898 5175
rect 1846 5111 1898 5117
rect 1846 5021 1898 5027
rect 1846 4963 1898 4969
rect 1750 3615 1802 3621
rect 1750 3557 1802 3563
rect 1858 800 1886 4963
rect 1942 3911 1994 3917
rect 1942 3853 1994 3859
rect 1954 800 1982 3853
rect 2050 800 2078 6295
rect 2146 3251 2174 8219
rect 3286 8219 3338 8225
rect 2228 8177 2284 8186
rect 2516 7650 2572 7659
rect 2516 7585 2518 7594
rect 2570 7585 2572 7594
rect 2518 7553 2570 7559
rect 2326 7463 2378 7469
rect 2326 7405 2378 7411
rect 2998 7463 3050 7469
rect 2998 7405 3050 7411
rect 2338 4139 2366 7405
rect 2518 7019 2570 7025
rect 2518 6961 2570 6967
rect 2326 4133 2378 4139
rect 2326 4075 2378 4081
rect 2422 4133 2474 4139
rect 2422 4075 2474 4081
rect 2326 3837 2378 3843
rect 2326 3779 2378 3785
rect 2134 3245 2186 3251
rect 2134 3187 2186 3193
rect 2134 2949 2186 2955
rect 2134 2891 2186 2897
rect 2146 800 2174 2891
rect 2338 800 2366 3779
rect 2434 800 2462 4075
rect 2530 800 2558 6961
rect 2902 5687 2954 5693
rect 2902 5629 2954 5635
rect 2710 3689 2762 3695
rect 2710 3631 2762 3637
rect 2722 800 2750 3631
rect 2914 2900 2942 5629
rect 3010 3917 3038 7405
rect 3190 6353 3242 6359
rect 3190 6295 3242 6301
rect 3094 5021 3146 5027
rect 3094 4963 3146 4969
rect 2998 3911 3050 3917
rect 2998 3853 3050 3859
rect 3106 3843 3134 4963
rect 3094 3837 3146 3843
rect 3094 3779 3146 3785
rect 2998 3763 3050 3769
rect 2998 3705 3050 3711
rect 2818 2872 2942 2900
rect 2818 800 2846 2872
rect 3010 2752 3038 3705
rect 3094 3541 3146 3547
rect 3094 3483 3146 3489
rect 2914 2724 3038 2752
rect 2914 800 2942 2724
rect 3106 1864 3134 3483
rect 3010 1836 3134 1864
rect 3010 800 3038 1836
rect 3202 800 3230 6295
rect 3298 3769 3326 8219
rect 3394 7765 3422 9625
rect 3382 7759 3434 7765
rect 3382 7701 3434 7707
rect 3586 5175 3614 56837
rect 3874 56531 3902 59200
rect 4354 57614 4382 59200
rect 4354 57586 4670 57614
rect 4268 57304 4564 57324
rect 4324 57302 4348 57304
rect 4404 57302 4428 57304
rect 4484 57302 4508 57304
rect 4346 57250 4348 57302
rect 4410 57250 4422 57302
rect 4484 57250 4486 57302
rect 4324 57248 4348 57250
rect 4404 57248 4428 57250
rect 4484 57248 4508 57250
rect 4268 57228 4564 57248
rect 3862 56525 3914 56531
rect 3862 56467 3914 56473
rect 4268 55972 4564 55992
rect 4324 55970 4348 55972
rect 4404 55970 4428 55972
rect 4484 55970 4508 55972
rect 4346 55918 4348 55970
rect 4410 55918 4422 55970
rect 4484 55918 4486 55970
rect 4324 55916 4348 55918
rect 4404 55916 4428 55918
rect 4484 55916 4508 55918
rect 4268 55896 4564 55916
rect 4642 55717 4670 57586
rect 4930 56975 4958 59200
rect 4918 56969 4970 56975
rect 4918 56911 4970 56917
rect 5110 56895 5162 56901
rect 5110 56837 5162 56843
rect 4726 56229 4778 56235
rect 4726 56171 4778 56177
rect 4630 55711 4682 55717
rect 4630 55653 4682 55659
rect 4630 55563 4682 55569
rect 4630 55505 4682 55511
rect 4268 54640 4564 54660
rect 4324 54638 4348 54640
rect 4404 54638 4428 54640
rect 4484 54638 4508 54640
rect 4346 54586 4348 54638
rect 4410 54586 4422 54638
rect 4484 54586 4486 54638
rect 4324 54584 4348 54586
rect 4404 54584 4428 54586
rect 4484 54584 4508 54586
rect 4268 54564 4564 54584
rect 3670 53565 3722 53571
rect 3670 53507 3722 53513
rect 3682 7913 3710 53507
rect 4268 53308 4564 53328
rect 4324 53306 4348 53308
rect 4404 53306 4428 53308
rect 4484 53306 4508 53308
rect 4346 53254 4348 53306
rect 4410 53254 4422 53306
rect 4484 53254 4486 53306
rect 4324 53252 4348 53254
rect 4404 53252 4428 53254
rect 4484 53252 4508 53254
rect 4268 53232 4564 53252
rect 4268 51976 4564 51996
rect 4324 51974 4348 51976
rect 4404 51974 4428 51976
rect 4484 51974 4508 51976
rect 4346 51922 4348 51974
rect 4410 51922 4422 51974
rect 4484 51922 4486 51974
rect 4324 51920 4348 51922
rect 4404 51920 4428 51922
rect 4484 51920 4508 51922
rect 4268 51900 4564 51920
rect 4268 50644 4564 50664
rect 4324 50642 4348 50644
rect 4404 50642 4428 50644
rect 4484 50642 4508 50644
rect 4346 50590 4348 50642
rect 4410 50590 4422 50642
rect 4484 50590 4486 50642
rect 4324 50588 4348 50590
rect 4404 50588 4428 50590
rect 4484 50588 4508 50590
rect 4268 50568 4564 50588
rect 4268 49312 4564 49332
rect 4324 49310 4348 49312
rect 4404 49310 4428 49312
rect 4484 49310 4508 49312
rect 4346 49258 4348 49310
rect 4410 49258 4422 49310
rect 4484 49258 4486 49310
rect 4324 49256 4348 49258
rect 4404 49256 4428 49258
rect 4484 49256 4508 49258
rect 4268 49236 4564 49256
rect 3766 48089 3818 48095
rect 3766 48031 3818 48037
rect 3778 8579 3806 48031
rect 4268 47980 4564 48000
rect 4324 47978 4348 47980
rect 4404 47978 4428 47980
rect 4484 47978 4508 47980
rect 4346 47926 4348 47978
rect 4410 47926 4422 47978
rect 4484 47926 4486 47978
rect 4324 47924 4348 47926
rect 4404 47924 4428 47926
rect 4484 47924 4508 47926
rect 4268 47904 4564 47924
rect 4268 46648 4564 46668
rect 4324 46646 4348 46648
rect 4404 46646 4428 46648
rect 4484 46646 4508 46648
rect 4346 46594 4348 46646
rect 4410 46594 4422 46646
rect 4484 46594 4486 46646
rect 4324 46592 4348 46594
rect 4404 46592 4428 46594
rect 4484 46592 4508 46594
rect 4268 46572 4564 46592
rect 4268 45316 4564 45336
rect 4324 45314 4348 45316
rect 4404 45314 4428 45316
rect 4484 45314 4508 45316
rect 4346 45262 4348 45314
rect 4410 45262 4422 45314
rect 4484 45262 4486 45314
rect 4324 45260 4348 45262
rect 4404 45260 4428 45262
rect 4484 45260 4508 45262
rect 4268 45240 4564 45260
rect 4268 43984 4564 44004
rect 4324 43982 4348 43984
rect 4404 43982 4428 43984
rect 4484 43982 4508 43984
rect 4346 43930 4348 43982
rect 4410 43930 4422 43982
rect 4484 43930 4486 43982
rect 4324 43928 4348 43930
rect 4404 43928 4428 43930
rect 4484 43928 4508 43930
rect 4268 43908 4564 43928
rect 4268 42652 4564 42672
rect 4324 42650 4348 42652
rect 4404 42650 4428 42652
rect 4484 42650 4508 42652
rect 4346 42598 4348 42650
rect 4410 42598 4422 42650
rect 4484 42598 4486 42650
rect 4324 42596 4348 42598
rect 4404 42596 4428 42598
rect 4484 42596 4508 42598
rect 4268 42576 4564 42596
rect 4268 41320 4564 41340
rect 4324 41318 4348 41320
rect 4404 41318 4428 41320
rect 4484 41318 4508 41320
rect 4346 41266 4348 41318
rect 4410 41266 4422 41318
rect 4484 41266 4486 41318
rect 4324 41264 4348 41266
rect 4404 41264 4428 41266
rect 4484 41264 4508 41266
rect 4268 41244 4564 41264
rect 4268 39988 4564 40008
rect 4324 39986 4348 39988
rect 4404 39986 4428 39988
rect 4484 39986 4508 39988
rect 4346 39934 4348 39986
rect 4410 39934 4422 39986
rect 4484 39934 4486 39986
rect 4324 39932 4348 39934
rect 4404 39932 4428 39934
rect 4484 39932 4508 39934
rect 4268 39912 4564 39932
rect 4268 38656 4564 38676
rect 4324 38654 4348 38656
rect 4404 38654 4428 38656
rect 4484 38654 4508 38656
rect 4346 38602 4348 38654
rect 4410 38602 4422 38654
rect 4484 38602 4486 38654
rect 4324 38600 4348 38602
rect 4404 38600 4428 38602
rect 4484 38600 4508 38602
rect 4268 38580 4564 38600
rect 4268 37324 4564 37344
rect 4324 37322 4348 37324
rect 4404 37322 4428 37324
rect 4484 37322 4508 37324
rect 4346 37270 4348 37322
rect 4410 37270 4422 37322
rect 4484 37270 4486 37322
rect 4324 37268 4348 37270
rect 4404 37268 4428 37270
rect 4484 37268 4508 37270
rect 4268 37248 4564 37268
rect 4268 35992 4564 36012
rect 4324 35990 4348 35992
rect 4404 35990 4428 35992
rect 4484 35990 4508 35992
rect 4346 35938 4348 35990
rect 4410 35938 4422 35990
rect 4484 35938 4486 35990
rect 4324 35936 4348 35938
rect 4404 35936 4428 35938
rect 4484 35936 4508 35938
rect 4268 35916 4564 35936
rect 4268 34660 4564 34680
rect 4324 34658 4348 34660
rect 4404 34658 4428 34660
rect 4484 34658 4508 34660
rect 4346 34606 4348 34658
rect 4410 34606 4422 34658
rect 4484 34606 4486 34658
rect 4324 34604 4348 34606
rect 4404 34604 4428 34606
rect 4484 34604 4508 34606
rect 4268 34584 4564 34604
rect 4268 33328 4564 33348
rect 4324 33326 4348 33328
rect 4404 33326 4428 33328
rect 4484 33326 4508 33328
rect 4346 33274 4348 33326
rect 4410 33274 4422 33326
rect 4484 33274 4486 33326
rect 4324 33272 4348 33274
rect 4404 33272 4428 33274
rect 4484 33272 4508 33274
rect 4268 33252 4564 33272
rect 4268 31996 4564 32016
rect 4324 31994 4348 31996
rect 4404 31994 4428 31996
rect 4484 31994 4508 31996
rect 4346 31942 4348 31994
rect 4410 31942 4422 31994
rect 4484 31942 4486 31994
rect 4324 31940 4348 31942
rect 4404 31940 4428 31942
rect 4484 31940 4508 31942
rect 4268 31920 4564 31940
rect 4268 30664 4564 30684
rect 4324 30662 4348 30664
rect 4404 30662 4428 30664
rect 4484 30662 4508 30664
rect 4346 30610 4348 30662
rect 4410 30610 4422 30662
rect 4484 30610 4486 30662
rect 4324 30608 4348 30610
rect 4404 30608 4428 30610
rect 4484 30608 4508 30610
rect 4268 30588 4564 30608
rect 4268 29332 4564 29352
rect 4324 29330 4348 29332
rect 4404 29330 4428 29332
rect 4484 29330 4508 29332
rect 4346 29278 4348 29330
rect 4410 29278 4422 29330
rect 4484 29278 4486 29330
rect 4324 29276 4348 29278
rect 4404 29276 4428 29278
rect 4484 29276 4508 29278
rect 4268 29256 4564 29276
rect 4268 28000 4564 28020
rect 4324 27998 4348 28000
rect 4404 27998 4428 28000
rect 4484 27998 4508 28000
rect 4346 27946 4348 27998
rect 4410 27946 4422 27998
rect 4484 27946 4486 27998
rect 4324 27944 4348 27946
rect 4404 27944 4428 27946
rect 4484 27944 4508 27946
rect 4268 27924 4564 27944
rect 4268 26668 4564 26688
rect 4324 26666 4348 26668
rect 4404 26666 4428 26668
rect 4484 26666 4508 26668
rect 4346 26614 4348 26666
rect 4410 26614 4422 26666
rect 4484 26614 4486 26666
rect 4324 26612 4348 26614
rect 4404 26612 4428 26614
rect 4484 26612 4508 26614
rect 4268 26592 4564 26612
rect 4268 25336 4564 25356
rect 4324 25334 4348 25336
rect 4404 25334 4428 25336
rect 4484 25334 4508 25336
rect 4346 25282 4348 25334
rect 4410 25282 4422 25334
rect 4484 25282 4486 25334
rect 4324 25280 4348 25282
rect 4404 25280 4428 25282
rect 4484 25280 4508 25282
rect 4268 25260 4564 25280
rect 4268 24004 4564 24024
rect 4324 24002 4348 24004
rect 4404 24002 4428 24004
rect 4484 24002 4508 24004
rect 4346 23950 4348 24002
rect 4410 23950 4422 24002
rect 4484 23950 4486 24002
rect 4324 23948 4348 23950
rect 4404 23948 4428 23950
rect 4484 23948 4508 23950
rect 4268 23928 4564 23948
rect 4268 22672 4564 22692
rect 4324 22670 4348 22672
rect 4404 22670 4428 22672
rect 4484 22670 4508 22672
rect 4346 22618 4348 22670
rect 4410 22618 4422 22670
rect 4484 22618 4486 22670
rect 4324 22616 4348 22618
rect 4404 22616 4428 22618
rect 4484 22616 4508 22618
rect 4268 22596 4564 22616
rect 4268 21340 4564 21360
rect 4324 21338 4348 21340
rect 4404 21338 4428 21340
rect 4484 21338 4508 21340
rect 4346 21286 4348 21338
rect 4410 21286 4422 21338
rect 4484 21286 4486 21338
rect 4324 21284 4348 21286
rect 4404 21284 4428 21286
rect 4484 21284 4508 21286
rect 4268 21264 4564 21284
rect 4268 20008 4564 20028
rect 4324 20006 4348 20008
rect 4404 20006 4428 20008
rect 4484 20006 4508 20008
rect 4346 19954 4348 20006
rect 4410 19954 4422 20006
rect 4484 19954 4486 20006
rect 4324 19952 4348 19954
rect 4404 19952 4428 19954
rect 4484 19952 4508 19954
rect 4268 19932 4564 19952
rect 4268 18676 4564 18696
rect 4324 18674 4348 18676
rect 4404 18674 4428 18676
rect 4484 18674 4508 18676
rect 4346 18622 4348 18674
rect 4410 18622 4422 18674
rect 4484 18622 4486 18674
rect 4324 18620 4348 18622
rect 4404 18620 4428 18622
rect 4484 18620 4508 18622
rect 4268 18600 4564 18620
rect 4268 17344 4564 17364
rect 4324 17342 4348 17344
rect 4404 17342 4428 17344
rect 4484 17342 4508 17344
rect 4346 17290 4348 17342
rect 4410 17290 4422 17342
rect 4484 17290 4486 17342
rect 4324 17288 4348 17290
rect 4404 17288 4428 17290
rect 4484 17288 4508 17290
rect 4268 17268 4564 17288
rect 4268 16012 4564 16032
rect 4324 16010 4348 16012
rect 4404 16010 4428 16012
rect 4484 16010 4508 16012
rect 4346 15958 4348 16010
rect 4410 15958 4422 16010
rect 4484 15958 4486 16010
rect 4324 15956 4348 15958
rect 4404 15956 4428 15958
rect 4484 15956 4508 15958
rect 4268 15936 4564 15956
rect 4268 14680 4564 14700
rect 4324 14678 4348 14680
rect 4404 14678 4428 14680
rect 4484 14678 4508 14680
rect 4346 14626 4348 14678
rect 4410 14626 4422 14678
rect 4484 14626 4486 14678
rect 4324 14624 4348 14626
rect 4404 14624 4428 14626
rect 4484 14624 4508 14626
rect 4268 14604 4564 14624
rect 4268 13348 4564 13368
rect 4324 13346 4348 13348
rect 4404 13346 4428 13348
rect 4484 13346 4508 13348
rect 4346 13294 4348 13346
rect 4410 13294 4422 13346
rect 4484 13294 4486 13346
rect 4324 13292 4348 13294
rect 4404 13292 4428 13294
rect 4484 13292 4508 13294
rect 4268 13272 4564 13292
rect 4268 12016 4564 12036
rect 4324 12014 4348 12016
rect 4404 12014 4428 12016
rect 4484 12014 4508 12016
rect 4346 11962 4348 12014
rect 4410 11962 4422 12014
rect 4484 11962 4486 12014
rect 4324 11960 4348 11962
rect 4404 11960 4428 11962
rect 4484 11960 4508 11962
rect 4268 11940 4564 11960
rect 4268 10684 4564 10704
rect 4324 10682 4348 10684
rect 4404 10682 4428 10684
rect 4484 10682 4508 10684
rect 4346 10630 4348 10682
rect 4410 10630 4422 10682
rect 4484 10630 4486 10682
rect 4324 10628 4348 10630
rect 4404 10628 4428 10630
rect 4484 10628 4508 10630
rect 4268 10608 4564 10628
rect 4268 9352 4564 9372
rect 4324 9350 4348 9352
rect 4404 9350 4428 9352
rect 4484 9350 4508 9352
rect 4346 9298 4348 9350
rect 4410 9298 4422 9350
rect 4484 9298 4486 9350
rect 4324 9296 4348 9298
rect 4404 9296 4428 9298
rect 4484 9296 4508 9298
rect 4268 9276 4564 9296
rect 3766 8573 3818 8579
rect 3766 8515 3818 8521
rect 4268 8020 4564 8040
rect 4324 8018 4348 8020
rect 4404 8018 4428 8020
rect 4484 8018 4508 8020
rect 4346 7966 4348 8018
rect 4410 7966 4422 8018
rect 4484 7966 4486 8018
rect 4324 7964 4348 7966
rect 4404 7964 4428 7966
rect 4484 7964 4508 7966
rect 4268 7944 4564 7964
rect 3670 7907 3722 7913
rect 3670 7849 3722 7855
rect 3958 7463 4010 7469
rect 3958 7405 4010 7411
rect 4054 7463 4106 7469
rect 4054 7405 4106 7411
rect 3670 7167 3722 7173
rect 3670 7109 3722 7115
rect 3574 5169 3626 5175
rect 3574 5111 3626 5117
rect 3478 4207 3530 4213
rect 3478 4149 3530 4155
rect 3286 3763 3338 3769
rect 3286 3705 3338 3711
rect 3382 3763 3434 3769
rect 3382 3705 3434 3711
rect 3286 3467 3338 3473
rect 3286 3409 3338 3415
rect 3298 800 3326 3409
rect 3394 800 3422 3705
rect 3490 800 3518 4149
rect 3682 800 3710 7109
rect 3862 6353 3914 6359
rect 3862 6295 3914 6301
rect 3766 4281 3818 4287
rect 3766 4223 3818 4229
rect 3778 800 3806 4223
rect 3874 800 3902 6295
rect 3970 3473 3998 7405
rect 3958 3467 4010 3473
rect 3958 3409 4010 3415
rect 3958 3245 4010 3251
rect 3958 3187 4010 3193
rect 3970 2585 3998 3187
rect 3958 2579 4010 2585
rect 3958 2521 4010 2527
rect 4066 800 4094 7405
rect 4534 6945 4586 6951
rect 4532 6910 4534 6919
rect 4586 6910 4588 6919
rect 4532 6845 4588 6854
rect 4268 6688 4564 6708
rect 4324 6686 4348 6688
rect 4404 6686 4428 6688
rect 4484 6686 4508 6688
rect 4346 6634 4348 6686
rect 4410 6634 4422 6686
rect 4484 6634 4486 6686
rect 4324 6632 4348 6634
rect 4404 6632 4428 6634
rect 4484 6632 4508 6634
rect 4268 6612 4564 6632
rect 4642 6452 4670 55505
rect 4738 10873 4766 56171
rect 4726 10867 4778 10873
rect 4726 10809 4778 10815
rect 4822 8203 4874 8209
rect 4822 8145 4874 8151
rect 4642 6424 4766 6452
rect 4630 6353 4682 6359
rect 4630 6295 4682 6301
rect 4268 5356 4564 5376
rect 4324 5354 4348 5356
rect 4404 5354 4428 5356
rect 4484 5354 4508 5356
rect 4346 5302 4348 5354
rect 4410 5302 4422 5354
rect 4484 5302 4486 5354
rect 4324 5300 4348 5302
rect 4404 5300 4428 5302
rect 4484 5300 4508 5302
rect 4268 5280 4564 5300
rect 4150 5021 4202 5027
rect 4150 4963 4202 4969
rect 4162 800 4190 4963
rect 4268 4024 4564 4044
rect 4324 4022 4348 4024
rect 4404 4022 4428 4024
rect 4484 4022 4508 4024
rect 4346 3970 4348 4022
rect 4410 3970 4422 4022
rect 4484 3970 4486 4022
rect 4324 3968 4348 3970
rect 4404 3968 4428 3970
rect 4484 3968 4508 3970
rect 4268 3948 4564 3968
rect 4268 2692 4564 2712
rect 4324 2690 4348 2692
rect 4404 2690 4428 2692
rect 4484 2690 4508 2692
rect 4346 2638 4348 2690
rect 4410 2638 4422 2690
rect 4484 2638 4486 2690
rect 4324 2636 4348 2638
rect 4404 2636 4428 2638
rect 4484 2636 4508 2638
rect 4268 2616 4564 2636
rect 4246 2579 4298 2585
rect 4246 2521 4298 2527
rect 4342 2579 4394 2585
rect 4342 2521 4394 2527
rect 4258 800 4286 2521
rect 4354 800 4382 2521
rect 4642 2456 4670 6295
rect 4738 5249 4766 6424
rect 4726 5243 4778 5249
rect 4726 5185 4778 5191
rect 4726 4355 4778 4361
rect 4726 4297 4778 4303
rect 4450 2428 4670 2456
rect 4450 2012 4478 2428
rect 4738 2160 4766 4297
rect 4834 2585 4862 8145
rect 4918 8129 4970 8135
rect 4918 8071 4970 8077
rect 4930 7765 4958 8071
rect 4918 7759 4970 7765
rect 4918 7701 4970 7707
rect 5014 6871 5066 6877
rect 5014 6813 5066 6819
rect 4918 5687 4970 5693
rect 4918 5629 4970 5635
rect 4930 4213 4958 5629
rect 4918 4207 4970 4213
rect 4918 4149 4970 4155
rect 5026 4139 5054 6813
rect 5122 6359 5150 56837
rect 5410 56531 5438 59200
rect 5986 56531 6014 59200
rect 6466 56975 6494 59200
rect 6454 56969 6506 56975
rect 6454 56911 6506 56917
rect 7042 56531 7070 59200
rect 5398 56525 5450 56531
rect 5398 56467 5450 56473
rect 5974 56525 6026 56531
rect 5974 56467 6026 56473
rect 7030 56525 7082 56531
rect 7030 56467 7082 56473
rect 6742 56303 6794 56309
rect 6742 56245 6794 56251
rect 5206 56229 5258 56235
rect 5206 56171 5258 56177
rect 6358 56229 6410 56235
rect 6358 56171 6410 56177
rect 5218 24193 5246 56171
rect 6370 29669 6398 56171
rect 6754 47059 6782 56245
rect 7222 56229 7274 56235
rect 7220 56194 7222 56203
rect 7274 56194 7276 56203
rect 7220 56129 7276 56138
rect 7522 55717 7550 59200
rect 8098 56975 8126 59200
rect 8086 56969 8138 56975
rect 8086 56911 8138 56917
rect 8278 56895 8330 56901
rect 8278 56837 8330 56843
rect 7510 55711 7562 55717
rect 7510 55653 7562 55659
rect 7702 55563 7754 55569
rect 7702 55505 7754 55511
rect 6742 47053 6794 47059
rect 6742 46995 6794 47001
rect 6742 39431 6794 39437
rect 6742 39373 6794 39379
rect 6358 29663 6410 29669
rect 6358 29605 6410 29611
rect 5686 25445 5738 25451
rect 5686 25387 5738 25393
rect 5206 24187 5258 24193
rect 5206 24129 5258 24135
rect 5206 8943 5258 8949
rect 5206 8885 5258 8891
rect 5110 6353 5162 6359
rect 5110 6295 5162 6301
rect 5218 5915 5246 8885
rect 5590 8203 5642 8209
rect 5590 8145 5642 8151
rect 5602 7765 5630 8145
rect 5590 7759 5642 7765
rect 5590 7701 5642 7707
rect 5302 7463 5354 7469
rect 5302 7405 5354 7411
rect 5206 5909 5258 5915
rect 5206 5851 5258 5857
rect 5206 5687 5258 5693
rect 5206 5629 5258 5635
rect 5110 4207 5162 4213
rect 5110 4149 5162 4155
rect 5014 4133 5066 4139
rect 5014 4075 5066 4081
rect 4918 3023 4970 3029
rect 4918 2965 4970 2971
rect 4822 2579 4874 2585
rect 4822 2521 4874 2527
rect 4738 2132 4862 2160
rect 4726 2061 4778 2067
rect 4450 1984 4670 2012
rect 4726 2003 4778 2009
rect 4534 1913 4586 1919
rect 4534 1855 4586 1861
rect 4546 800 4574 1855
rect 4642 800 4670 1984
rect 4738 800 4766 2003
rect 4834 1919 4862 2132
rect 4822 1913 4874 1919
rect 4822 1855 4874 1861
rect 4930 800 4958 2965
rect 5122 2894 5150 4149
rect 5218 3251 5246 5629
rect 5206 3245 5258 3251
rect 5206 3187 5258 3193
rect 5206 3023 5258 3029
rect 5206 2965 5258 2971
rect 5026 2866 5150 2894
rect 5026 800 5054 2866
rect 5110 2801 5162 2807
rect 5110 2743 5162 2749
rect 5122 800 5150 2743
rect 5218 800 5246 2965
rect 5314 2067 5342 7405
rect 5398 7093 5450 7099
rect 5396 7058 5398 7067
rect 5450 7058 5452 7067
rect 5396 6993 5452 7002
rect 5698 6433 5726 25387
rect 6550 12125 6602 12131
rect 6550 12067 6602 12073
rect 6562 7247 6590 12067
rect 6754 7363 6782 39373
rect 6838 37877 6890 37883
rect 6838 37819 6890 37825
rect 6740 7354 6796 7363
rect 6740 7289 6796 7298
rect 6550 7241 6602 7247
rect 6550 7183 6602 7189
rect 5878 6945 5930 6951
rect 5878 6887 5930 6893
rect 6166 6945 6218 6951
rect 6166 6887 6218 6893
rect 6550 6945 6602 6951
rect 6550 6887 6602 6893
rect 5686 6427 5738 6433
rect 5686 6369 5738 6375
rect 5494 6131 5546 6137
rect 5494 6073 5546 6079
rect 5398 5021 5450 5027
rect 5398 4963 5450 4969
rect 5302 2061 5354 2067
rect 5302 2003 5354 2009
rect 5410 800 5438 4963
rect 5506 800 5534 6073
rect 5782 5613 5834 5619
rect 5782 5555 5834 5561
rect 5686 4281 5738 4287
rect 5686 4223 5738 4229
rect 5590 3689 5642 3695
rect 5590 3631 5642 3637
rect 5602 800 5630 3631
rect 5698 800 5726 4223
rect 5794 2955 5822 5555
rect 5782 2949 5834 2955
rect 5782 2891 5834 2897
rect 5890 800 5918 6887
rect 6070 5021 6122 5027
rect 6070 4963 6122 4969
rect 5974 3023 6026 3029
rect 5974 2965 6026 2971
rect 5986 800 6014 2965
rect 6082 800 6110 4963
rect 6178 2881 6206 6887
rect 6262 6131 6314 6137
rect 6262 6073 6314 6079
rect 6166 2875 6218 2881
rect 6166 2817 6218 2823
rect 6274 800 6302 6073
rect 6454 4207 6506 4213
rect 6454 4149 6506 4155
rect 6358 3689 6410 3695
rect 6358 3631 6410 3637
rect 6370 800 6398 3631
rect 6466 800 6494 4149
rect 6562 800 6590 6887
rect 6850 6581 6878 37819
rect 7126 27887 7178 27893
rect 7126 27829 7178 27835
rect 7138 22491 7166 27829
rect 7714 26783 7742 55505
rect 8290 36014 8318 56837
rect 8578 56531 8606 59200
rect 8566 56525 8618 56531
rect 8566 56467 8618 56473
rect 8566 56229 8618 56235
rect 8566 56171 8618 56177
rect 8470 44907 8522 44913
rect 8470 44849 8522 44855
rect 8098 35986 8318 36014
rect 8098 33134 8126 35986
rect 8482 33134 8510 44849
rect 8578 35663 8606 56171
rect 9154 55717 9182 59200
rect 9634 57049 9662 59200
rect 9622 57043 9674 57049
rect 9622 56985 9674 56991
rect 9718 56747 9770 56753
rect 9718 56689 9770 56695
rect 9142 55711 9194 55717
rect 9142 55653 9194 55659
rect 8950 55415 9002 55421
rect 8950 55357 9002 55363
rect 8566 35657 8618 35663
rect 8566 35599 8618 35605
rect 8098 33106 8318 33134
rect 8482 33106 8606 33134
rect 8290 28814 8318 33106
rect 8374 29145 8426 29151
rect 8374 29087 8426 29093
rect 8386 28971 8414 29087
rect 8372 28962 8428 28971
rect 8372 28897 8428 28906
rect 8290 28786 8510 28814
rect 8374 27739 8426 27745
rect 8374 27681 8426 27687
rect 7702 26777 7754 26783
rect 7702 26719 7754 26725
rect 8086 26407 8138 26413
rect 8086 26349 8138 26355
rect 7942 26333 7994 26339
rect 7942 26275 7994 26281
rect 7954 26136 7982 26275
rect 7714 26108 7982 26136
rect 7220 24966 7276 24975
rect 7220 24901 7276 24910
rect 7126 22485 7178 22491
rect 7126 22427 7178 22433
rect 7030 18933 7082 18939
rect 7030 18875 7082 18881
rect 7042 11909 7070 18875
rect 7126 18119 7178 18125
rect 7126 18061 7178 18067
rect 7030 11903 7082 11909
rect 7030 11845 7082 11851
rect 7030 9905 7082 9911
rect 7030 9847 7082 9853
rect 7042 9245 7070 9847
rect 7030 9239 7082 9245
rect 7030 9181 7082 9187
rect 6934 7241 6986 7247
rect 6934 7183 6986 7189
rect 6838 6575 6890 6581
rect 6838 6517 6890 6523
rect 6838 5687 6890 5693
rect 6838 5629 6890 5635
rect 6742 2949 6794 2955
rect 6742 2891 6794 2897
rect 6754 800 6782 2891
rect 6850 800 6878 5629
rect 6946 800 6974 7183
rect 7138 6008 7166 18061
rect 7234 15184 7262 24901
rect 7414 23891 7466 23897
rect 7414 23833 7466 23839
rect 7318 23225 7370 23231
rect 7318 23167 7370 23173
rect 7330 18125 7358 23167
rect 7426 18144 7454 23833
rect 7714 22565 7742 26108
rect 7942 24927 7994 24933
rect 7942 24869 7994 24875
rect 7954 24656 7982 24869
rect 8098 24804 8126 26349
rect 8386 26159 8414 27681
rect 8372 26150 8428 26159
rect 8372 26085 8428 26094
rect 8374 25001 8426 25007
rect 8228 24966 8284 24975
rect 8374 24943 8426 24949
rect 8228 24901 8230 24910
rect 8282 24901 8284 24910
rect 8230 24869 8282 24875
rect 8098 24776 8318 24804
rect 7810 24628 7982 24656
rect 7810 23897 7838 24628
rect 8182 24557 8234 24563
rect 8182 24499 8234 24505
rect 7798 23891 7850 23897
rect 7798 23833 7850 23839
rect 8086 23669 8138 23675
rect 7810 23617 8086 23620
rect 7810 23611 8138 23617
rect 7810 23592 8126 23611
rect 7510 22559 7562 22565
rect 7510 22501 7562 22507
rect 7702 22559 7754 22565
rect 7702 22501 7754 22507
rect 7522 18791 7550 22501
rect 7606 22485 7658 22491
rect 7606 22427 7658 22433
rect 7510 18785 7562 18791
rect 7510 18727 7562 18733
rect 7318 18119 7370 18125
rect 7426 18116 7550 18144
rect 7318 18061 7370 18067
rect 7412 17270 7468 17279
rect 7412 17205 7414 17214
rect 7466 17205 7468 17214
rect 7414 17173 7466 17179
rect 7414 16121 7466 16127
rect 7414 16063 7466 16069
rect 7426 15905 7454 16063
rect 7414 15899 7466 15905
rect 7414 15841 7466 15847
rect 7234 15156 7454 15184
rect 7222 13013 7274 13019
rect 7222 12955 7274 12961
rect 7042 5980 7166 6008
rect 7042 4084 7070 5980
rect 7234 5860 7262 12955
rect 7318 11903 7370 11909
rect 7318 11845 7370 11851
rect 7330 7215 7358 11845
rect 7316 7206 7372 7215
rect 7316 7141 7372 7150
rect 7318 6871 7370 6877
rect 7318 6813 7370 6819
rect 7138 5832 7262 5860
rect 7138 5471 7166 5832
rect 7222 5687 7274 5693
rect 7222 5629 7274 5635
rect 7126 5465 7178 5471
rect 7126 5407 7178 5413
rect 7042 4056 7166 4084
rect 7030 3689 7082 3695
rect 7030 3631 7082 3637
rect 7042 800 7070 3631
rect 7138 3177 7166 4056
rect 7126 3171 7178 3177
rect 7126 3113 7178 3119
rect 7234 800 7262 5629
rect 7330 800 7358 6813
rect 7426 4583 7454 15156
rect 7522 13241 7550 18116
rect 7510 13235 7562 13241
rect 7510 13177 7562 13183
rect 7618 13112 7646 22427
rect 7702 22411 7754 22417
rect 7702 22353 7754 22359
rect 7522 13084 7646 13112
rect 7522 8547 7550 13084
rect 7606 12569 7658 12575
rect 7606 12511 7658 12517
rect 7508 8538 7564 8547
rect 7618 8505 7646 12511
rect 7508 8473 7564 8482
rect 7606 8499 7658 8505
rect 7606 8441 7658 8447
rect 7714 8376 7742 22353
rect 7810 18939 7838 23592
rect 7942 23521 7994 23527
rect 7906 23469 7942 23472
rect 7906 23463 7994 23469
rect 7906 23444 7982 23463
rect 7906 22787 7934 23444
rect 8194 23324 8222 24499
rect 8002 23296 8222 23324
rect 7894 22781 7946 22787
rect 7894 22723 7946 22729
rect 7894 22485 7946 22491
rect 7894 22427 7946 22433
rect 7798 18933 7850 18939
rect 7798 18875 7850 18881
rect 7798 18785 7850 18791
rect 7798 18727 7850 18733
rect 7810 13431 7838 18727
rect 7906 15165 7934 22427
rect 7894 15159 7946 15165
rect 7894 15101 7946 15107
rect 8002 13556 8030 23296
rect 8086 22781 8138 22787
rect 8086 22723 8138 22729
rect 8098 19624 8126 22723
rect 8290 22565 8318 24776
rect 8386 24119 8414 24943
rect 8374 24113 8426 24119
rect 8374 24055 8426 24061
rect 8374 23595 8426 23601
rect 8374 23537 8426 23543
rect 8386 23231 8414 23537
rect 8374 23225 8426 23231
rect 8374 23167 8426 23173
rect 8482 23054 8510 28786
rect 8578 24563 8606 33106
rect 8758 28775 8810 28781
rect 8758 28717 8810 28723
rect 8770 25988 8798 28717
rect 8854 27443 8906 27449
rect 8854 27385 8906 27391
rect 8674 25960 8798 25988
rect 8566 24557 8618 24563
rect 8566 24499 8618 24505
rect 8566 24113 8618 24119
rect 8566 24055 8618 24061
rect 8386 23026 8510 23054
rect 8278 22559 8330 22565
rect 8278 22501 8330 22507
rect 8278 22115 8330 22121
rect 8278 22057 8330 22063
rect 8290 21899 8318 22057
rect 8278 21893 8330 21899
rect 8278 21835 8330 21841
rect 8278 21597 8330 21603
rect 8278 21539 8330 21545
rect 8290 21252 8318 21539
rect 8242 21224 8318 21252
rect 8242 21011 8270 21224
rect 8230 21005 8282 21011
rect 8230 20947 8282 20953
rect 8278 20783 8330 20789
rect 8278 20725 8330 20731
rect 8290 20567 8318 20725
rect 8278 20561 8330 20567
rect 8278 20503 8330 20509
rect 8098 19596 8222 19624
rect 8086 19525 8138 19531
rect 8086 19467 8138 19473
rect 8098 19235 8126 19467
rect 8086 19229 8138 19235
rect 8086 19171 8138 19177
rect 8194 18736 8222 19596
rect 7906 13528 8030 13556
rect 8098 18708 8222 18736
rect 7796 13422 7852 13431
rect 7796 13357 7852 13366
rect 7906 13223 7934 13528
rect 7988 13422 8044 13431
rect 7988 13357 8044 13366
rect 7810 13195 7934 13223
rect 7810 12575 7838 13195
rect 8002 13112 8030 13357
rect 7906 13084 8030 13112
rect 7798 12569 7850 12575
rect 7798 12511 7850 12517
rect 7798 11237 7850 11243
rect 7798 11179 7850 11185
rect 7522 8348 7742 8376
rect 7414 4577 7466 4583
rect 7414 4519 7466 4525
rect 7414 4355 7466 4361
rect 7414 4297 7466 4303
rect 7426 800 7454 4297
rect 7522 3473 7550 8348
rect 7606 8277 7658 8283
rect 7606 8219 7658 8225
rect 7702 8277 7754 8283
rect 7702 8219 7754 8225
rect 7618 7807 7646 8219
rect 7604 7798 7660 7807
rect 7604 7733 7660 7742
rect 7606 7463 7658 7469
rect 7606 7405 7658 7411
rect 7618 7247 7646 7405
rect 7606 7241 7658 7247
rect 7606 7183 7658 7189
rect 7606 7019 7658 7025
rect 7606 6961 7658 6967
rect 7618 5841 7646 6961
rect 7606 5835 7658 5841
rect 7606 5777 7658 5783
rect 7606 5539 7658 5545
rect 7606 5481 7658 5487
rect 7510 3467 7562 3473
rect 7510 3409 7562 3415
rect 7618 800 7646 5481
rect 7714 800 7742 8219
rect 7810 4084 7838 11179
rect 7906 8672 7934 13084
rect 8098 11243 8126 18708
rect 8230 18287 8282 18293
rect 8230 18229 8282 18235
rect 8242 17996 8270 18229
rect 8194 17968 8270 17996
rect 8194 17829 8222 17968
rect 8182 17823 8234 17829
rect 8182 17765 8234 17771
rect 8182 16121 8234 16127
rect 8182 16063 8234 16069
rect 8194 15905 8222 16063
rect 8182 15899 8234 15905
rect 8182 15841 8234 15847
rect 8182 15529 8234 15535
rect 8182 15471 8234 15477
rect 8194 15239 8222 15471
rect 8182 15233 8234 15239
rect 8182 15175 8234 15181
rect 8278 15159 8330 15165
rect 8278 15101 8330 15107
rect 8182 13457 8234 13463
rect 8182 13399 8234 13405
rect 8194 13241 8222 13399
rect 8182 13235 8234 13241
rect 8182 13177 8234 13183
rect 8086 11237 8138 11243
rect 8086 11179 8138 11185
rect 8086 11089 8138 11095
rect 8086 11031 8138 11037
rect 7990 10793 8042 10799
rect 7990 10735 8042 10741
rect 8002 9837 8030 10735
rect 8098 10429 8126 11031
rect 8182 10571 8234 10577
rect 8182 10513 8234 10519
rect 8086 10423 8138 10429
rect 8086 10365 8138 10371
rect 7990 9831 8042 9837
rect 7990 9773 8042 9779
rect 8086 9535 8138 9541
rect 8086 9477 8138 9483
rect 8098 9023 8126 9477
rect 8086 9017 8138 9023
rect 8086 8959 8138 8965
rect 7906 8644 8126 8672
rect 7892 8538 7948 8547
rect 7892 8473 7948 8482
rect 7906 7913 7934 8473
rect 7988 8390 8044 8399
rect 7988 8325 8044 8334
rect 7894 7907 7946 7913
rect 7894 7849 7946 7855
rect 7892 7206 7948 7215
rect 7892 7141 7948 7150
rect 7906 4287 7934 7141
rect 7894 4281 7946 4287
rect 8002 4255 8030 8325
rect 8098 4509 8126 8644
rect 8086 4503 8138 4509
rect 8086 4445 8138 4451
rect 8084 4394 8140 4403
rect 8084 4329 8140 4338
rect 7894 4223 7946 4229
rect 7988 4246 8044 4255
rect 7988 4181 8044 4190
rect 7810 4056 8030 4084
rect 7894 3911 7946 3917
rect 7894 3853 7946 3859
rect 7798 3689 7850 3695
rect 7798 3631 7850 3637
rect 7810 800 7838 3631
rect 7906 800 7934 3853
rect 8002 3621 8030 4056
rect 7990 3615 8042 3621
rect 7990 3557 8042 3563
rect 8098 800 8126 4329
rect 8194 3251 8222 10513
rect 8290 9856 8318 15101
rect 8386 10004 8414 23026
rect 8470 22559 8522 22565
rect 8470 22501 8522 22507
rect 8482 10577 8510 22501
rect 8470 10571 8522 10577
rect 8470 10513 8522 10519
rect 8386 9976 8510 10004
rect 8290 9828 8414 9856
rect 8278 9757 8330 9763
rect 8386 9731 8414 9828
rect 8278 9699 8330 9705
rect 8372 9722 8428 9731
rect 8290 9245 8318 9699
rect 8372 9657 8428 9666
rect 8374 9609 8426 9615
rect 8374 9551 8426 9557
rect 8278 9239 8330 9245
rect 8278 9181 8330 9187
rect 8386 9153 8414 9551
rect 8290 9125 8414 9153
rect 8290 4435 8318 9125
rect 8482 7895 8510 9976
rect 8578 9615 8606 24055
rect 8674 23054 8702 25960
rect 8674 23026 8798 23054
rect 8662 18563 8714 18569
rect 8662 18505 8714 18511
rect 8674 18125 8702 18505
rect 8662 18119 8714 18125
rect 8662 18061 8714 18067
rect 8662 17897 8714 17903
rect 8662 17839 8714 17845
rect 8566 9609 8618 9615
rect 8566 9551 8618 9557
rect 8566 9461 8618 9467
rect 8566 9403 8618 9409
rect 8578 9171 8606 9403
rect 8566 9165 8618 9171
rect 8674 9139 8702 17839
rect 8770 10133 8798 23026
rect 8758 10127 8810 10133
rect 8758 10069 8810 10075
rect 8758 9905 8810 9911
rect 8758 9847 8810 9853
rect 8770 9171 8798 9847
rect 8758 9165 8810 9171
rect 8566 9107 8618 9113
rect 8660 9130 8716 9139
rect 8758 9107 8810 9113
rect 8660 9065 8716 9074
rect 8564 8982 8620 8991
rect 8756 8982 8812 8991
rect 8564 8917 8620 8926
rect 8662 8943 8714 8949
rect 8578 8376 8606 8917
rect 8714 8926 8756 8931
rect 8714 8917 8812 8926
rect 8714 8903 8798 8917
rect 8662 8885 8714 8891
rect 8578 8348 8702 8376
rect 8566 8277 8618 8283
rect 8564 8242 8566 8251
rect 8618 8242 8620 8251
rect 8564 8177 8620 8186
rect 8386 7867 8510 7895
rect 8564 7946 8620 7955
rect 8564 7881 8620 7890
rect 8386 6433 8414 7867
rect 8578 7747 8606 7881
rect 8530 7719 8606 7747
rect 8530 7691 8558 7719
rect 8518 7685 8570 7691
rect 8518 7627 8570 7633
rect 8468 7502 8524 7511
rect 8468 7437 8524 7446
rect 8566 7463 8618 7469
rect 8374 6427 8426 6433
rect 8374 6369 8426 6375
rect 8278 4429 8330 4435
rect 8278 4371 8330 4377
rect 8278 3837 8330 3843
rect 8278 3779 8330 3785
rect 8182 3245 8234 3251
rect 8182 3187 8234 3193
rect 8182 3023 8234 3029
rect 8182 2965 8234 2971
rect 8194 800 8222 2965
rect 8290 800 8318 3779
rect 8482 800 8510 7437
rect 8566 7405 8618 7411
rect 8578 7247 8606 7405
rect 8566 7241 8618 7247
rect 8566 7183 8618 7189
rect 8674 7155 8702 8348
rect 8756 7798 8812 7807
rect 8756 7733 8812 7742
rect 8770 7691 8798 7733
rect 8758 7685 8810 7691
rect 8758 7627 8810 7633
rect 8758 7537 8810 7543
rect 8756 7502 8758 7511
rect 8810 7502 8812 7511
rect 8756 7437 8812 7446
rect 8578 7127 8702 7155
rect 8578 3811 8606 7127
rect 8758 7093 8810 7099
rect 8758 7035 8810 7041
rect 8770 6211 8798 7035
rect 8866 6581 8894 27385
rect 8854 6575 8906 6581
rect 8854 6517 8906 6523
rect 8962 6507 8990 55357
rect 9046 29219 9098 29225
rect 9046 29161 9098 29167
rect 9058 17903 9086 29161
rect 9238 26111 9290 26117
rect 9238 26053 9290 26059
rect 9142 25001 9194 25007
rect 9142 24943 9194 24949
rect 9046 17897 9098 17903
rect 9046 17839 9098 17845
rect 9044 17270 9100 17279
rect 9044 17205 9046 17214
rect 9098 17205 9100 17214
rect 9046 17173 9098 17179
rect 9154 10281 9182 24943
rect 9142 10275 9194 10281
rect 9142 10217 9194 10223
rect 9142 10127 9194 10133
rect 9142 10069 9194 10075
rect 9046 9017 9098 9023
rect 9044 8982 9046 8991
rect 9098 8982 9100 8991
rect 9044 8917 9100 8926
rect 9046 8869 9098 8875
rect 9046 8811 9098 8817
rect 9058 7955 9086 8811
rect 9044 7946 9100 7955
rect 9044 7881 9100 7890
rect 9154 7599 9182 10069
rect 9058 7571 9182 7599
rect 8950 6501 9002 6507
rect 8950 6443 9002 6449
rect 9058 6285 9086 7571
rect 9142 7463 9194 7469
rect 9142 7405 9194 7411
rect 9046 6279 9098 6285
rect 9046 6221 9098 6227
rect 8758 6205 8810 6211
rect 8758 6147 8810 6153
rect 8758 5687 8810 5693
rect 8758 5629 8810 5635
rect 8770 4232 8798 5629
rect 8854 4799 8906 4805
rect 8854 4741 8906 4747
rect 8674 4204 8798 4232
rect 8564 3802 8620 3811
rect 8564 3737 8620 3746
rect 8566 3689 8618 3695
rect 8566 3631 8618 3637
rect 8578 800 8606 3631
rect 8674 800 8702 4204
rect 8866 3492 8894 4741
rect 8950 4503 9002 4509
rect 8950 4445 9002 4451
rect 8770 3464 8894 3492
rect 8770 800 8798 3464
rect 8962 3103 8990 4445
rect 9046 4133 9098 4139
rect 9046 4075 9098 4081
rect 8950 3097 9002 3103
rect 8950 3039 9002 3045
rect 8950 2949 9002 2955
rect 8950 2891 9002 2897
rect 8962 800 8990 2891
rect 9058 800 9086 4075
rect 9154 800 9182 7405
rect 9250 6137 9278 26053
rect 9622 25223 9674 25229
rect 9622 25165 9674 25171
rect 9334 20783 9386 20789
rect 9334 20725 9386 20731
rect 9346 20567 9374 20725
rect 9334 20561 9386 20567
rect 9334 20503 9386 20509
rect 9634 12974 9662 25165
rect 9538 12946 9662 12974
rect 9334 10275 9386 10281
rect 9334 10217 9386 10223
rect 9238 6131 9290 6137
rect 9238 6073 9290 6079
rect 9238 5021 9290 5027
rect 9238 4963 9290 4969
rect 9250 3917 9278 4963
rect 9346 4213 9374 10217
rect 9430 8795 9482 8801
rect 9430 8737 9482 8743
rect 9442 8209 9470 8737
rect 9538 8265 9566 12946
rect 9622 10941 9674 10947
rect 9622 10883 9674 10889
rect 9634 10503 9662 10883
rect 9622 10497 9674 10503
rect 9622 10439 9674 10445
rect 9622 9831 9674 9837
rect 9622 9773 9674 9779
rect 9634 8579 9662 9773
rect 9622 8573 9674 8579
rect 9622 8515 9674 8521
rect 9538 8237 9662 8265
rect 9430 8203 9482 8209
rect 9430 8145 9482 8151
rect 9526 8203 9578 8209
rect 9526 8145 9578 8151
rect 9428 7946 9484 7955
rect 9428 7881 9484 7890
rect 9442 7765 9470 7881
rect 9430 7759 9482 7765
rect 9430 7701 9482 7707
rect 9538 7099 9566 8145
rect 9526 7093 9578 7099
rect 9526 7035 9578 7041
rect 9526 6945 9578 6951
rect 9526 6887 9578 6893
rect 9430 6353 9482 6359
rect 9430 6295 9482 6301
rect 9334 4207 9386 4213
rect 9334 4149 9386 4155
rect 9238 3911 9290 3917
rect 9238 3853 9290 3859
rect 9334 3689 9386 3695
rect 9334 3631 9386 3637
rect 9346 2894 9374 3631
rect 9250 2866 9374 2894
rect 9250 800 9278 2866
rect 9442 800 9470 6295
rect 9538 800 9566 6887
rect 9634 6433 9662 8237
rect 9730 7913 9758 56689
rect 10210 56531 10238 59200
rect 10690 56531 10718 59200
rect 11266 57049 11294 59200
rect 11254 57043 11306 57049
rect 11254 56985 11306 56991
rect 11254 56895 11306 56901
rect 11254 56837 11306 56843
rect 10198 56525 10250 56531
rect 10198 56467 10250 56473
rect 10678 56525 10730 56531
rect 10678 56467 10730 56473
rect 10582 56229 10634 56235
rect 10582 56171 10634 56177
rect 11158 56229 11210 56235
rect 11158 56171 11210 56177
rect 9910 46239 9962 46245
rect 9910 46181 9962 46187
rect 9922 7913 9950 46181
rect 10594 36014 10622 56171
rect 11170 44987 11198 56171
rect 11158 44981 11210 44987
rect 11158 44923 11210 44929
rect 10594 35986 10718 36014
rect 10006 21449 10058 21455
rect 10006 21391 10058 21397
rect 10018 12353 10046 21391
rect 10690 12974 10718 35986
rect 10774 20857 10826 20863
rect 10774 20799 10826 20805
rect 10786 20567 10814 20799
rect 10774 20561 10826 20567
rect 10774 20503 10826 20509
rect 10690 12946 10814 12974
rect 10006 12347 10058 12353
rect 10006 12289 10058 12295
rect 10006 12199 10058 12205
rect 10006 12141 10058 12147
rect 9718 7907 9770 7913
rect 9718 7849 9770 7855
rect 9910 7907 9962 7913
rect 9910 7849 9962 7855
rect 10018 7839 10046 12141
rect 10294 8277 10346 8283
rect 10294 8219 10346 8225
rect 10678 8277 10730 8283
rect 10678 8219 10730 8225
rect 10006 7833 10058 7839
rect 10006 7775 10058 7781
rect 10196 7798 10252 7807
rect 10196 7733 10198 7742
rect 10250 7733 10252 7742
rect 10198 7701 10250 7707
rect 9910 7537 9962 7543
rect 9908 7502 9910 7511
rect 9962 7502 9964 7511
rect 9908 7437 9964 7446
rect 10054 7167 10106 7173
rect 9826 7127 10054 7155
rect 9826 7025 9854 7127
rect 10054 7109 10106 7115
rect 9814 7019 9866 7025
rect 9814 6961 9866 6967
rect 9718 6945 9770 6951
rect 9718 6887 9770 6893
rect 9910 6945 9962 6951
rect 9910 6887 9962 6893
rect 10004 6910 10060 6919
rect 9622 6427 9674 6433
rect 9622 6369 9674 6375
rect 9730 4551 9758 6887
rect 9922 4805 9950 6887
rect 10004 6845 10006 6854
rect 10058 6845 10060 6854
rect 10006 6813 10058 6819
rect 10102 6353 10154 6359
rect 10102 6295 10154 6301
rect 9910 4799 9962 4805
rect 9910 4741 9962 4747
rect 9716 4542 9772 4551
rect 9716 4477 9772 4486
rect 9622 4355 9674 4361
rect 9622 4297 9674 4303
rect 9634 800 9662 4297
rect 9814 4281 9866 4287
rect 9814 4223 9866 4229
rect 9826 3917 9854 4223
rect 9908 3950 9964 3959
rect 9814 3911 9866 3917
rect 9908 3885 9964 3894
rect 9814 3853 9866 3859
rect 9814 2579 9866 2585
rect 9814 2521 9866 2527
rect 9826 800 9854 2521
rect 9922 800 9950 3885
rect 10006 3541 10058 3547
rect 10006 3483 10058 3489
rect 10018 800 10046 3483
rect 10114 800 10142 6295
rect 10198 5687 10250 5693
rect 10198 5629 10250 5635
rect 10210 2585 10238 5629
rect 10198 2579 10250 2585
rect 10198 2521 10250 2527
rect 10306 800 10334 8219
rect 10582 6945 10634 6951
rect 10580 6910 10582 6919
rect 10634 6910 10636 6919
rect 10580 6845 10636 6854
rect 10582 6575 10634 6581
rect 10582 6517 10634 6523
rect 10486 5687 10538 5693
rect 10486 5629 10538 5635
rect 10390 4355 10442 4361
rect 10390 4297 10442 4303
rect 10402 800 10430 4297
rect 10498 800 10526 5629
rect 10594 5619 10622 6517
rect 10582 5613 10634 5619
rect 10582 5555 10634 5561
rect 10582 5021 10634 5027
rect 10582 4963 10634 4969
rect 10594 3843 10622 4963
rect 10582 3837 10634 3843
rect 10582 3779 10634 3785
rect 10582 3689 10634 3695
rect 10582 3631 10634 3637
rect 10594 3547 10622 3631
rect 10582 3541 10634 3547
rect 10582 3483 10634 3489
rect 10690 2894 10718 8219
rect 10786 4509 10814 12946
rect 11158 10793 11210 10799
rect 11158 10735 11210 10741
rect 10966 8869 11018 8875
rect 10868 8834 10924 8843
rect 10966 8811 11018 8817
rect 10868 8769 10924 8778
rect 10882 8579 10910 8769
rect 10870 8573 10922 8579
rect 10870 8515 10922 8521
rect 10870 7019 10922 7025
rect 10870 6961 10922 6967
rect 10882 6771 10910 6961
rect 10868 6762 10924 6771
rect 10868 6697 10924 6706
rect 10978 6581 11006 8811
rect 11060 8686 11116 8695
rect 11060 8621 11116 8630
rect 11074 7691 11102 8621
rect 11062 7685 11114 7691
rect 11062 7627 11114 7633
rect 11062 7463 11114 7469
rect 11062 7405 11114 7411
rect 10966 6575 11018 6581
rect 10966 6517 11018 6523
rect 10870 6353 10922 6359
rect 10870 6295 10922 6301
rect 10774 4503 10826 4509
rect 10774 4445 10826 4451
rect 10774 4355 10826 4361
rect 10774 4297 10826 4303
rect 10594 2866 10718 2894
rect 10594 800 10622 2866
rect 10786 800 10814 4297
rect 10882 800 10910 6295
rect 10966 5021 11018 5027
rect 10966 4963 11018 4969
rect 10978 4139 11006 4963
rect 10966 4133 11018 4139
rect 10966 4075 11018 4081
rect 11074 2894 11102 7405
rect 11170 6507 11198 10735
rect 11266 8949 11294 56837
rect 11746 56531 11774 59200
rect 12322 56531 12350 59200
rect 12802 56975 12830 59200
rect 12790 56969 12842 56975
rect 12790 56911 12842 56917
rect 12982 56895 13034 56901
rect 12982 56837 13034 56843
rect 11734 56525 11786 56531
rect 11734 56467 11786 56473
rect 12310 56525 12362 56531
rect 12310 56467 12362 56473
rect 11542 56229 11594 56235
rect 11542 56171 11594 56177
rect 12694 56229 12746 56235
rect 12694 56171 12746 56177
rect 11350 37433 11402 37439
rect 11350 37375 11402 37381
rect 11254 8943 11306 8949
rect 11254 8885 11306 8891
rect 11362 8875 11390 37375
rect 11554 29521 11582 56171
rect 11926 49421 11978 49427
rect 11926 49363 11978 49369
rect 11542 29515 11594 29521
rect 11542 29457 11594 29463
rect 11638 24113 11690 24119
rect 11638 24055 11690 24061
rect 11446 13457 11498 13463
rect 11446 13399 11498 13405
rect 11458 8949 11486 13399
rect 11650 10355 11678 24055
rect 11638 10349 11690 10355
rect 11638 10291 11690 10297
rect 11446 8943 11498 8949
rect 11446 8885 11498 8891
rect 11350 8869 11402 8875
rect 11350 8811 11402 8817
rect 11542 8573 11594 8579
rect 11362 8521 11542 8524
rect 11362 8515 11594 8521
rect 11362 8496 11582 8515
rect 11254 7019 11306 7025
rect 11254 6961 11306 6967
rect 11158 6501 11210 6507
rect 11158 6443 11210 6449
rect 11158 4207 11210 4213
rect 11158 4149 11210 4155
rect 10978 2866 11102 2894
rect 10978 800 11006 2866
rect 11170 800 11198 4149
rect 11266 800 11294 6961
rect 11362 800 11390 8496
rect 11446 8277 11498 8283
rect 11446 8219 11498 8225
rect 11458 7839 11486 8219
rect 11446 7833 11498 7839
rect 11446 7775 11498 7781
rect 11938 7765 11966 49363
rect 12214 40763 12266 40769
rect 12214 40705 12266 40711
rect 12226 12974 12254 40705
rect 12706 33443 12734 56171
rect 12694 33437 12746 33443
rect 12694 33379 12746 33385
rect 12406 23595 12458 23601
rect 12406 23537 12458 23543
rect 12310 22781 12362 22787
rect 12310 22723 12362 22729
rect 12034 12946 12254 12974
rect 11926 7759 11978 7765
rect 11926 7701 11978 7707
rect 11734 7537 11786 7543
rect 11734 7479 11786 7485
rect 11638 6353 11690 6359
rect 11638 6295 11690 6301
rect 11542 5465 11594 5471
rect 11542 5407 11594 5413
rect 11554 4509 11582 5407
rect 11446 4503 11498 4509
rect 11446 4445 11498 4451
rect 11542 4503 11594 4509
rect 11542 4445 11594 4451
rect 11458 4380 11486 4445
rect 11458 4352 11582 4380
rect 11446 4281 11498 4287
rect 11446 4223 11498 4229
rect 11458 800 11486 4223
rect 11554 3917 11582 4352
rect 11542 3911 11594 3917
rect 11542 3853 11594 3859
rect 11650 800 11678 6295
rect 11746 800 11774 7479
rect 12034 5767 12062 12946
rect 12214 8425 12266 8431
rect 12214 8367 12266 8373
rect 12118 8277 12170 8283
rect 12118 8219 12170 8225
rect 12130 7913 12158 8219
rect 12118 7907 12170 7913
rect 12118 7849 12170 7855
rect 12226 7340 12254 8367
rect 12130 7312 12254 7340
rect 12022 5761 12074 5767
rect 12022 5703 12074 5709
rect 11830 5021 11882 5027
rect 11830 4963 11882 4969
rect 11842 800 11870 4963
rect 11926 4133 11978 4139
rect 11926 4075 11978 4081
rect 11938 3473 11966 4075
rect 11926 3467 11978 3473
rect 11926 3409 11978 3415
rect 12022 3467 12074 3473
rect 12022 3409 12074 3415
rect 12034 800 12062 3409
rect 12130 800 12158 7312
rect 12212 7206 12268 7215
rect 12322 7173 12350 22723
rect 12418 8399 12446 23537
rect 12598 9091 12650 9097
rect 12598 9033 12650 9039
rect 12502 8573 12554 8579
rect 12502 8515 12554 8521
rect 12404 8390 12460 8399
rect 12514 8357 12542 8515
rect 12610 8357 12638 9033
rect 12994 8547 13022 56837
rect 13378 56531 13406 59200
rect 13366 56525 13418 56531
rect 13366 56467 13418 56473
rect 13558 56229 13610 56235
rect 13558 56171 13610 56177
rect 13570 38327 13598 56171
rect 13858 55717 13886 59200
rect 14434 56975 14462 59200
rect 14422 56969 14474 56975
rect 14422 56911 14474 56917
rect 14914 56531 14942 59200
rect 14902 56525 14954 56531
rect 14902 56467 14954 56473
rect 15286 56377 15338 56383
rect 15286 56319 15338 56325
rect 14710 56229 14762 56235
rect 14710 56171 14762 56177
rect 13846 55711 13898 55717
rect 13846 55653 13898 55659
rect 13654 55415 13706 55421
rect 13654 55357 13706 55363
rect 13558 38321 13610 38327
rect 13558 38263 13610 38269
rect 13666 12131 13694 55357
rect 14230 38099 14282 38105
rect 14230 38041 14282 38047
rect 13942 32105 13994 32111
rect 13942 32047 13994 32053
rect 13654 12125 13706 12131
rect 13654 12067 13706 12073
rect 13174 8943 13226 8949
rect 13174 8885 13226 8891
rect 12980 8538 13036 8547
rect 13186 8505 13214 8885
rect 13954 8875 13982 32047
rect 14134 29589 14186 29595
rect 14134 29531 14186 29537
rect 14146 29225 14174 29531
rect 14134 29219 14186 29225
rect 14134 29161 14186 29167
rect 13942 8869 13994 8875
rect 13942 8811 13994 8817
rect 13652 8538 13708 8547
rect 12980 8473 13036 8482
rect 13174 8499 13226 8505
rect 13652 8473 13708 8482
rect 13174 8441 13226 8447
rect 13666 8431 13694 8473
rect 13654 8425 13706 8431
rect 13654 8367 13706 8373
rect 12404 8325 12460 8334
rect 12502 8351 12554 8357
rect 12502 8293 12554 8299
rect 12598 8351 12650 8357
rect 12598 8293 12650 8299
rect 13174 8277 13226 8283
rect 12898 8237 13174 8265
rect 12598 7537 12650 7543
rect 12598 7479 12650 7485
rect 12610 7451 12638 7479
rect 12514 7423 12638 7451
rect 12212 7141 12268 7150
rect 12310 7167 12362 7173
rect 12226 7099 12254 7141
rect 12310 7109 12362 7115
rect 12214 7093 12266 7099
rect 12214 7035 12266 7041
rect 12310 6353 12362 6359
rect 12310 6295 12362 6301
rect 12214 4873 12266 4879
rect 12214 4815 12266 4821
rect 12226 800 12254 4815
rect 12322 800 12350 6295
rect 12514 800 12542 7423
rect 12788 7354 12844 7363
rect 12788 7289 12844 7298
rect 12802 7247 12830 7289
rect 12790 7241 12842 7247
rect 12790 7183 12842 7189
rect 12694 7019 12746 7025
rect 12694 6961 12746 6967
rect 12598 5687 12650 5693
rect 12598 5629 12650 5635
rect 12610 800 12638 5629
rect 12706 800 12734 6961
rect 12898 4195 12926 8237
rect 13174 8219 13226 8225
rect 12982 8203 13034 8209
rect 12982 8145 13034 8151
rect 12994 8080 13022 8145
rect 12994 8052 13214 8080
rect 13186 7469 13214 8052
rect 13270 7759 13322 7765
rect 13270 7701 13322 7707
rect 13174 7463 13226 7469
rect 13174 7405 13226 7411
rect 13282 7363 13310 7701
rect 13942 7611 13994 7617
rect 13942 7553 13994 7559
rect 13954 7511 13982 7553
rect 13940 7502 13996 7511
rect 13940 7437 13996 7446
rect 13268 7354 13324 7363
rect 13268 7289 13324 7298
rect 14242 7173 14270 38041
rect 14326 27591 14378 27597
rect 14326 27533 14378 27539
rect 13174 7167 13226 7173
rect 13174 7109 13226 7115
rect 14230 7167 14282 7173
rect 14230 7109 14282 7115
rect 13078 7093 13130 7099
rect 13078 7035 13130 7041
rect 12982 7019 13034 7025
rect 12982 6961 13034 6967
rect 12994 6771 13022 6961
rect 12980 6762 13036 6771
rect 12980 6697 13036 6706
rect 13090 6304 13118 7035
rect 12994 6285 13118 6304
rect 12982 6279 13118 6285
rect 13034 6276 13118 6279
rect 12982 6221 13034 6227
rect 13078 6205 13130 6211
rect 13186 6156 13214 7109
rect 13462 6945 13514 6951
rect 13462 6887 13514 6893
rect 13130 6153 13214 6156
rect 13078 6147 13214 6153
rect 13090 6128 13214 6147
rect 13270 6131 13322 6137
rect 13270 6073 13322 6079
rect 12802 4167 12926 4195
rect 12802 800 12830 4167
rect 13078 4133 13130 4139
rect 13078 4075 13130 4081
rect 13090 3177 13118 4075
rect 13174 3689 13226 3695
rect 13174 3631 13226 3637
rect 13078 3171 13130 3177
rect 13078 3113 13130 3119
rect 12982 3023 13034 3029
rect 12982 2965 13034 2971
rect 12994 800 13022 2965
rect 13078 2579 13130 2585
rect 13078 2521 13130 2527
rect 13090 800 13118 2521
rect 13186 800 13214 3631
rect 13282 2585 13310 6073
rect 13366 5687 13418 5693
rect 13366 5629 13418 5635
rect 13378 3473 13406 5629
rect 13366 3467 13418 3473
rect 13366 3409 13418 3415
rect 13366 3023 13418 3029
rect 13366 2965 13418 2971
rect 13270 2579 13322 2585
rect 13270 2521 13322 2527
rect 13378 800 13406 2965
rect 13474 800 13502 6887
rect 13846 6575 13898 6581
rect 13846 6517 13898 6523
rect 13858 6433 13886 6517
rect 13846 6427 13898 6433
rect 13846 6369 13898 6375
rect 14338 6304 14366 27533
rect 14722 25747 14750 56171
rect 15298 38845 15326 56319
rect 15394 56161 15422 59200
rect 15970 56975 15998 59200
rect 16450 57049 16478 59200
rect 16630 57191 16682 57197
rect 16630 57133 16682 57139
rect 16438 57043 16490 57049
rect 16438 56985 16490 56991
rect 15958 56969 16010 56975
rect 15958 56911 16010 56917
rect 15574 56895 15626 56901
rect 15574 56837 15626 56843
rect 16150 56895 16202 56901
rect 16150 56837 16202 56843
rect 15478 56229 15530 56235
rect 15478 56171 15530 56177
rect 15382 56155 15434 56161
rect 15382 56097 15434 56103
rect 15286 38839 15338 38845
rect 15286 38781 15338 38787
rect 15094 36915 15146 36921
rect 15094 36857 15146 36863
rect 14998 36101 15050 36107
rect 14998 36043 15050 36049
rect 14806 34769 14858 34775
rect 14806 34711 14858 34717
rect 14710 25741 14762 25747
rect 14710 25683 14762 25689
rect 14614 24927 14666 24933
rect 14614 24869 14666 24875
rect 14626 7617 14654 24869
rect 14710 21893 14762 21899
rect 14710 21835 14762 21841
rect 14614 7611 14666 7617
rect 14614 7553 14666 7559
rect 14518 6945 14570 6951
rect 14518 6887 14570 6893
rect 14614 6945 14666 6951
rect 14614 6887 14666 6893
rect 14530 6581 14558 6887
rect 14518 6575 14570 6581
rect 14518 6517 14570 6523
rect 14242 6276 14366 6304
rect 14242 5767 14270 6276
rect 14518 6131 14570 6137
rect 14518 6073 14570 6079
rect 14230 5761 14282 5767
rect 14230 5703 14282 5709
rect 13942 5021 13994 5027
rect 13942 4963 13994 4969
rect 14422 5021 14474 5027
rect 14422 4963 14474 4969
rect 13558 4355 13610 4361
rect 13558 4297 13610 4303
rect 13570 800 13598 4297
rect 13846 4281 13898 4287
rect 13846 4223 13898 4229
rect 13748 3802 13804 3811
rect 13748 3737 13804 3746
rect 13654 3689 13706 3695
rect 13654 3631 13706 3637
rect 13666 800 13694 3631
rect 13762 3251 13790 3737
rect 13750 3245 13802 3251
rect 13750 3187 13802 3193
rect 13858 800 13886 4223
rect 13954 800 13982 4963
rect 14134 4207 14186 4213
rect 14134 4149 14186 4155
rect 14038 3689 14090 3695
rect 14038 3631 14090 3637
rect 14050 800 14078 3631
rect 14146 800 14174 4149
rect 14230 3467 14282 3473
rect 14230 3409 14282 3415
rect 14242 2955 14270 3409
rect 14230 2949 14282 2955
rect 14230 2891 14282 2897
rect 14434 2894 14462 4963
rect 14530 4287 14558 6073
rect 14518 4281 14570 4287
rect 14518 4223 14570 4229
rect 14518 3023 14570 3029
rect 14518 2965 14570 2971
rect 14338 2866 14462 2894
rect 14338 800 14366 2866
rect 14530 1568 14558 2965
rect 14434 1540 14558 1568
rect 14434 800 14462 1540
rect 14626 1420 14654 6887
rect 14722 6433 14750 21835
rect 14818 8283 14846 34711
rect 15010 8801 15038 36043
rect 14998 8795 15050 8801
rect 14998 8737 15050 8743
rect 14806 8277 14858 8283
rect 14806 8219 14858 8225
rect 15106 6433 15134 36857
rect 15286 28923 15338 28929
rect 15286 28865 15338 28871
rect 15298 7543 15326 28865
rect 15490 17294 15518 56171
rect 15586 53053 15614 56837
rect 15958 56229 16010 56235
rect 15958 56171 16010 56177
rect 15574 53047 15626 53053
rect 15574 52989 15626 52995
rect 15670 49421 15722 49427
rect 15670 49363 15722 49369
rect 15574 20931 15626 20937
rect 15574 20873 15626 20879
rect 15394 17266 15518 17294
rect 15394 7765 15422 17266
rect 15586 12974 15614 20873
rect 15490 12946 15614 12974
rect 15382 7759 15434 7765
rect 15382 7701 15434 7707
rect 15490 7691 15518 12946
rect 15682 9097 15710 49363
rect 15766 43575 15818 43581
rect 15766 43517 15818 43523
rect 15670 9091 15722 9097
rect 15670 9033 15722 9039
rect 15778 7765 15806 43517
rect 15862 23891 15914 23897
rect 15862 23833 15914 23839
rect 15766 7759 15818 7765
rect 15766 7701 15818 7707
rect 15478 7685 15530 7691
rect 15670 7685 15722 7691
rect 15478 7627 15530 7633
rect 15586 7633 15670 7636
rect 15586 7627 15722 7633
rect 15586 7608 15710 7627
rect 15286 7537 15338 7543
rect 15286 7479 15338 7485
rect 15586 7469 15614 7608
rect 15574 7463 15626 7469
rect 15574 7405 15626 7411
rect 15670 7463 15722 7469
rect 15670 7405 15722 7411
rect 15286 7167 15338 7173
rect 15286 7109 15338 7115
rect 15298 6951 15326 7109
rect 15286 6945 15338 6951
rect 15286 6887 15338 6893
rect 15382 6945 15434 6951
rect 15382 6887 15434 6893
rect 14710 6427 14762 6433
rect 14710 6369 14762 6375
rect 15094 6427 15146 6433
rect 15094 6369 15146 6375
rect 14902 6205 14954 6211
rect 14902 6147 14954 6153
rect 14710 6131 14762 6137
rect 14710 6073 14762 6079
rect 14722 4213 14750 6073
rect 14806 5021 14858 5027
rect 14806 4963 14858 4969
rect 14710 4207 14762 4213
rect 14710 4149 14762 4155
rect 14818 3936 14846 4963
rect 14530 1392 14654 1420
rect 14722 3908 14846 3936
rect 14530 800 14558 1392
rect 14722 800 14750 3908
rect 14806 3689 14858 3695
rect 14806 3631 14858 3637
rect 14818 800 14846 3631
rect 14914 800 14942 6147
rect 14998 5687 15050 5693
rect 14998 5629 15050 5635
rect 15010 800 15038 5629
rect 15286 3689 15338 3695
rect 15286 3631 15338 3637
rect 15298 3344 15326 3631
rect 15202 3316 15326 3344
rect 15202 800 15230 3316
rect 15394 3196 15422 6887
rect 15478 4355 15530 4361
rect 15478 4297 15530 4303
rect 15298 3168 15422 3196
rect 15298 800 15326 3168
rect 15382 3097 15434 3103
rect 15382 3039 15434 3045
rect 15394 800 15422 3039
rect 15490 800 15518 4297
rect 15682 800 15710 7405
rect 15874 6951 15902 23833
rect 15970 13907 15998 56171
rect 15958 13901 16010 13907
rect 15958 13843 16010 13849
rect 16162 9763 16190 56837
rect 16534 56451 16586 56457
rect 16534 56393 16586 56399
rect 16246 26185 16298 26191
rect 16246 26127 16298 26133
rect 16150 9757 16202 9763
rect 16150 9699 16202 9705
rect 16150 8869 16202 8875
rect 16150 8811 16202 8817
rect 16054 8351 16106 8357
rect 16054 8293 16106 8299
rect 15958 8277 16010 8283
rect 15958 8219 16010 8225
rect 15970 7913 15998 8219
rect 15958 7907 16010 7913
rect 15958 7849 16010 7855
rect 15862 6945 15914 6951
rect 15862 6887 15914 6893
rect 15862 5687 15914 5693
rect 15862 5629 15914 5635
rect 15874 2894 15902 5629
rect 15958 4355 16010 4361
rect 15958 4297 16010 4303
rect 15778 2866 15902 2894
rect 15778 800 15806 2866
rect 15970 2160 15998 4297
rect 15874 2132 15998 2160
rect 15874 800 15902 2132
rect 16066 800 16094 8293
rect 16162 7765 16190 8811
rect 16258 8283 16286 26127
rect 16546 19531 16574 56393
rect 16642 20789 16670 57133
rect 17026 56531 17054 59200
rect 17506 56975 17534 59200
rect 17494 56969 17546 56975
rect 17494 56911 17546 56917
rect 17974 56895 18026 56901
rect 17974 56837 18026 56843
rect 17014 56525 17066 56531
rect 17014 56467 17066 56473
rect 17590 53417 17642 53423
rect 17590 53359 17642 53365
rect 16630 20783 16682 20789
rect 16630 20725 16682 20731
rect 16534 19525 16586 19531
rect 16534 19467 16586 19473
rect 17014 8869 17066 8875
rect 16436 8834 16492 8843
rect 17014 8811 17066 8817
rect 16436 8769 16492 8778
rect 16340 8686 16396 8695
rect 16340 8621 16396 8630
rect 16354 8431 16382 8621
rect 16342 8425 16394 8431
rect 16342 8367 16394 8373
rect 16450 8357 16478 8769
rect 16438 8351 16490 8357
rect 16438 8293 16490 8299
rect 17026 8283 17054 8811
rect 16246 8277 16298 8283
rect 16246 8219 16298 8225
rect 16342 8277 16394 8283
rect 16342 8219 16394 8225
rect 17014 8277 17066 8283
rect 17014 8219 17066 8225
rect 16150 7759 16202 7765
rect 16150 7701 16202 7707
rect 16150 5687 16202 5693
rect 16150 5629 16202 5635
rect 16162 800 16190 5629
rect 16246 4207 16298 4213
rect 16246 4149 16298 4155
rect 16258 800 16286 4149
rect 16354 800 16382 8219
rect 17110 6945 17162 6951
rect 17110 6887 17162 6893
rect 17302 6945 17354 6951
rect 17302 6887 17354 6893
rect 16726 6427 16778 6433
rect 16726 6369 16778 6375
rect 16438 5021 16490 5027
rect 16438 4963 16490 4969
rect 16450 3103 16478 4963
rect 16534 3911 16586 3917
rect 16534 3853 16586 3859
rect 16438 3097 16490 3103
rect 16438 3039 16490 3045
rect 16546 800 16574 3853
rect 16630 3023 16682 3029
rect 16630 2965 16682 2971
rect 16642 800 16670 2965
rect 16738 800 16766 6369
rect 16822 4133 16874 4139
rect 16822 4075 16874 4081
rect 16918 4133 16970 4139
rect 16918 4075 16970 4081
rect 16834 3251 16862 4075
rect 16822 3245 16874 3251
rect 16822 3187 16874 3193
rect 16930 800 16958 4075
rect 17014 3023 17066 3029
rect 17014 2965 17066 2971
rect 17026 800 17054 2965
rect 17122 800 17150 6887
rect 17314 6359 17342 6887
rect 17494 6797 17546 6803
rect 17494 6739 17546 6745
rect 17506 6581 17534 6739
rect 17494 6575 17546 6581
rect 17494 6517 17546 6523
rect 17302 6353 17354 6359
rect 17302 6295 17354 6301
rect 17602 6179 17630 53359
rect 17686 30773 17738 30779
rect 17686 30715 17738 30721
rect 17698 6433 17726 30715
rect 17782 29441 17834 29447
rect 17782 29383 17834 29389
rect 17794 11021 17822 29383
rect 17986 12974 18014 56837
rect 18082 56531 18110 59200
rect 18562 56531 18590 59200
rect 19138 56975 19166 59200
rect 19618 57614 19646 59200
rect 19618 57586 20030 57614
rect 19126 56969 19178 56975
rect 19126 56911 19178 56917
rect 19318 56895 19370 56901
rect 19318 56837 19370 56843
rect 18070 56525 18122 56531
rect 18070 56467 18122 56473
rect 18550 56525 18602 56531
rect 18550 56467 18602 56473
rect 18262 56229 18314 56235
rect 18262 56171 18314 56177
rect 19030 56229 19082 56235
rect 19030 56171 19082 56177
rect 18274 50093 18302 56171
rect 18358 52085 18410 52091
rect 18358 52027 18410 52033
rect 18262 50087 18314 50093
rect 18262 50029 18314 50035
rect 18070 38099 18122 38105
rect 18070 38041 18122 38047
rect 18082 37883 18110 38041
rect 18070 37877 18122 37883
rect 18070 37819 18122 37825
rect 17890 12946 18014 12974
rect 17782 11015 17834 11021
rect 17782 10957 17834 10963
rect 17890 9541 17918 12946
rect 17974 12347 18026 12353
rect 17974 12289 18026 12295
rect 17986 11761 18014 12289
rect 17974 11755 18026 11761
rect 17974 11697 18026 11703
rect 17878 9535 17930 9541
rect 17878 9477 17930 9483
rect 17794 6979 18206 7007
rect 17794 6951 17822 6979
rect 18178 6951 18206 6979
rect 17782 6945 17834 6951
rect 17782 6887 17834 6893
rect 17878 6945 17930 6951
rect 17878 6887 17930 6893
rect 18166 6945 18218 6951
rect 18166 6887 18218 6893
rect 17686 6427 17738 6433
rect 17686 6369 17738 6375
rect 17588 6170 17644 6179
rect 17494 6131 17546 6137
rect 17588 6105 17644 6114
rect 17494 6073 17546 6079
rect 17398 5687 17450 5693
rect 17398 5629 17450 5635
rect 17302 5021 17354 5027
rect 17302 4963 17354 4969
rect 17314 2894 17342 4963
rect 17410 3917 17438 5629
rect 17398 3911 17450 3917
rect 17398 3853 17450 3859
rect 17398 3689 17450 3695
rect 17398 3631 17450 3637
rect 17218 2866 17342 2894
rect 17218 800 17246 2866
rect 17410 800 17438 3631
rect 17506 800 17534 6073
rect 17794 5883 17822 6887
rect 17780 5874 17836 5883
rect 17780 5809 17836 5818
rect 17590 4429 17642 4435
rect 17590 4371 17642 4377
rect 17602 800 17630 4371
rect 17686 2949 17738 2955
rect 17686 2891 17738 2897
rect 17698 800 17726 2891
rect 17890 800 17918 6887
rect 18370 6623 18398 52027
rect 19042 34775 19070 56171
rect 19030 34769 19082 34775
rect 19030 34711 19082 34717
rect 19222 29441 19274 29447
rect 19222 29383 19274 29389
rect 18454 14863 18506 14869
rect 18454 14805 18506 14811
rect 18356 6614 18412 6623
rect 18356 6549 18412 6558
rect 18466 6433 18494 14805
rect 18838 8277 18890 8283
rect 18838 8219 18890 8225
rect 18850 7617 18878 8219
rect 18838 7611 18890 7617
rect 18838 7553 18890 7559
rect 18932 7354 18988 7363
rect 18932 7289 18988 7298
rect 18550 6945 18602 6951
rect 18550 6887 18602 6893
rect 18454 6427 18506 6433
rect 18454 6369 18506 6375
rect 18454 6131 18506 6137
rect 18454 6073 18506 6079
rect 17974 5021 18026 5027
rect 17974 4963 18026 4969
rect 17986 800 18014 4963
rect 18466 4528 18494 6073
rect 18274 4500 18494 4528
rect 18070 3689 18122 3695
rect 18070 3631 18122 3637
rect 18082 800 18110 3631
rect 18274 800 18302 4500
rect 18358 3911 18410 3917
rect 18358 3853 18410 3859
rect 18370 800 18398 3853
rect 18454 3689 18506 3695
rect 18454 3631 18506 3637
rect 18466 800 18494 3631
rect 18562 800 18590 6887
rect 18946 6877 18974 7289
rect 19030 7167 19082 7173
rect 19030 7109 19082 7115
rect 18934 6871 18986 6877
rect 18934 6813 18986 6819
rect 19042 6507 19070 7109
rect 19234 6951 19262 29383
rect 19330 9467 19358 56837
rect 19628 56638 19924 56658
rect 19684 56636 19708 56638
rect 19764 56636 19788 56638
rect 19844 56636 19868 56638
rect 19706 56584 19708 56636
rect 19770 56584 19782 56636
rect 19844 56584 19846 56636
rect 19684 56582 19708 56584
rect 19764 56582 19788 56584
rect 19844 56582 19868 56584
rect 19628 56562 19924 56582
rect 20002 56531 20030 57586
rect 19990 56525 20042 56531
rect 19990 56467 20042 56473
rect 20194 55717 20222 59200
rect 20674 56975 20702 59200
rect 20662 56969 20714 56975
rect 20662 56911 20714 56917
rect 20854 56895 20906 56901
rect 20854 56837 20906 56843
rect 20566 56229 20618 56235
rect 20566 56171 20618 56177
rect 20182 55711 20234 55717
rect 20182 55653 20234 55659
rect 20374 55563 20426 55569
rect 20374 55505 20426 55511
rect 19628 55306 19924 55326
rect 19684 55304 19708 55306
rect 19764 55304 19788 55306
rect 19844 55304 19868 55306
rect 19706 55252 19708 55304
rect 19770 55252 19782 55304
rect 19844 55252 19846 55304
rect 19684 55250 19708 55252
rect 19764 55250 19788 55252
rect 19844 55250 19868 55252
rect 19628 55230 19924 55250
rect 19628 53974 19924 53994
rect 19684 53972 19708 53974
rect 19764 53972 19788 53974
rect 19844 53972 19868 53974
rect 19706 53920 19708 53972
rect 19770 53920 19782 53972
rect 19844 53920 19846 53972
rect 19684 53918 19708 53920
rect 19764 53918 19788 53920
rect 19844 53918 19868 53920
rect 19628 53898 19924 53918
rect 19628 52642 19924 52662
rect 19684 52640 19708 52642
rect 19764 52640 19788 52642
rect 19844 52640 19868 52642
rect 19706 52588 19708 52640
rect 19770 52588 19782 52640
rect 19844 52588 19846 52640
rect 19684 52586 19708 52588
rect 19764 52586 19788 52588
rect 19844 52586 19868 52588
rect 19628 52566 19924 52586
rect 19628 51310 19924 51330
rect 19684 51308 19708 51310
rect 19764 51308 19788 51310
rect 19844 51308 19868 51310
rect 19706 51256 19708 51308
rect 19770 51256 19782 51308
rect 19844 51256 19846 51308
rect 19684 51254 19708 51256
rect 19764 51254 19788 51256
rect 19844 51254 19868 51256
rect 19628 51234 19924 51254
rect 19628 49978 19924 49998
rect 19684 49976 19708 49978
rect 19764 49976 19788 49978
rect 19844 49976 19868 49978
rect 19706 49924 19708 49976
rect 19770 49924 19782 49976
rect 19844 49924 19846 49976
rect 19684 49922 19708 49924
rect 19764 49922 19788 49924
rect 19844 49922 19868 49924
rect 19628 49902 19924 49922
rect 19628 48646 19924 48666
rect 19684 48644 19708 48646
rect 19764 48644 19788 48646
rect 19844 48644 19868 48646
rect 19706 48592 19708 48644
rect 19770 48592 19782 48644
rect 19844 48592 19846 48644
rect 19684 48590 19708 48592
rect 19764 48590 19788 48592
rect 19844 48590 19868 48592
rect 19628 48570 19924 48590
rect 19628 47314 19924 47334
rect 19684 47312 19708 47314
rect 19764 47312 19788 47314
rect 19844 47312 19868 47314
rect 19706 47260 19708 47312
rect 19770 47260 19782 47312
rect 19844 47260 19846 47312
rect 19684 47258 19708 47260
rect 19764 47258 19788 47260
rect 19844 47258 19868 47260
rect 19628 47238 19924 47258
rect 19628 45982 19924 46002
rect 19684 45980 19708 45982
rect 19764 45980 19788 45982
rect 19844 45980 19868 45982
rect 19706 45928 19708 45980
rect 19770 45928 19782 45980
rect 19844 45928 19846 45980
rect 19684 45926 19708 45928
rect 19764 45926 19788 45928
rect 19844 45926 19868 45928
rect 19628 45906 19924 45926
rect 19990 45203 20042 45209
rect 19990 45145 20042 45151
rect 19628 44650 19924 44670
rect 19684 44648 19708 44650
rect 19764 44648 19788 44650
rect 19844 44648 19868 44650
rect 19706 44596 19708 44648
rect 19770 44596 19782 44648
rect 19844 44596 19846 44648
rect 19684 44594 19708 44596
rect 19764 44594 19788 44596
rect 19844 44594 19868 44596
rect 19628 44574 19924 44594
rect 19628 43318 19924 43338
rect 19684 43316 19708 43318
rect 19764 43316 19788 43318
rect 19844 43316 19868 43318
rect 19706 43264 19708 43316
rect 19770 43264 19782 43316
rect 19844 43264 19846 43316
rect 19684 43262 19708 43264
rect 19764 43262 19788 43264
rect 19844 43262 19868 43264
rect 19628 43242 19924 43262
rect 19628 41986 19924 42006
rect 19684 41984 19708 41986
rect 19764 41984 19788 41986
rect 19844 41984 19868 41986
rect 19706 41932 19708 41984
rect 19770 41932 19782 41984
rect 19844 41932 19846 41984
rect 19684 41930 19708 41932
rect 19764 41930 19788 41932
rect 19844 41930 19868 41932
rect 19628 41910 19924 41930
rect 19628 40654 19924 40674
rect 19684 40652 19708 40654
rect 19764 40652 19788 40654
rect 19844 40652 19868 40654
rect 19706 40600 19708 40652
rect 19770 40600 19782 40652
rect 19844 40600 19846 40652
rect 19684 40598 19708 40600
rect 19764 40598 19788 40600
rect 19844 40598 19868 40600
rect 19628 40578 19924 40598
rect 19628 39322 19924 39342
rect 19684 39320 19708 39322
rect 19764 39320 19788 39322
rect 19844 39320 19868 39322
rect 19706 39268 19708 39320
rect 19770 39268 19782 39320
rect 19844 39268 19846 39320
rect 19684 39266 19708 39268
rect 19764 39266 19788 39268
rect 19844 39266 19868 39268
rect 19628 39246 19924 39266
rect 19628 37990 19924 38010
rect 19684 37988 19708 37990
rect 19764 37988 19788 37990
rect 19844 37988 19868 37990
rect 19706 37936 19708 37988
rect 19770 37936 19782 37988
rect 19844 37936 19846 37988
rect 19684 37934 19708 37936
rect 19764 37934 19788 37936
rect 19844 37934 19868 37936
rect 19628 37914 19924 37934
rect 19628 36658 19924 36678
rect 19684 36656 19708 36658
rect 19764 36656 19788 36658
rect 19844 36656 19868 36658
rect 19706 36604 19708 36656
rect 19770 36604 19782 36656
rect 19844 36604 19846 36656
rect 19684 36602 19708 36604
rect 19764 36602 19788 36604
rect 19844 36602 19868 36604
rect 19628 36582 19924 36602
rect 19628 35326 19924 35346
rect 19684 35324 19708 35326
rect 19764 35324 19788 35326
rect 19844 35324 19868 35326
rect 19706 35272 19708 35324
rect 19770 35272 19782 35324
rect 19844 35272 19846 35324
rect 19684 35270 19708 35272
rect 19764 35270 19788 35272
rect 19844 35270 19868 35272
rect 19628 35250 19924 35270
rect 19628 33994 19924 34014
rect 19684 33992 19708 33994
rect 19764 33992 19788 33994
rect 19844 33992 19868 33994
rect 19706 33940 19708 33992
rect 19770 33940 19782 33992
rect 19844 33940 19846 33992
rect 19684 33938 19708 33940
rect 19764 33938 19788 33940
rect 19844 33938 19868 33940
rect 19628 33918 19924 33938
rect 19628 32662 19924 32682
rect 19684 32660 19708 32662
rect 19764 32660 19788 32662
rect 19844 32660 19868 32662
rect 19706 32608 19708 32660
rect 19770 32608 19782 32660
rect 19844 32608 19846 32660
rect 19684 32606 19708 32608
rect 19764 32606 19788 32608
rect 19844 32606 19868 32608
rect 19628 32586 19924 32606
rect 19628 31330 19924 31350
rect 19684 31328 19708 31330
rect 19764 31328 19788 31330
rect 19844 31328 19868 31330
rect 19706 31276 19708 31328
rect 19770 31276 19782 31328
rect 19844 31276 19846 31328
rect 19684 31274 19708 31276
rect 19764 31274 19788 31276
rect 19844 31274 19868 31276
rect 19628 31254 19924 31274
rect 19628 29998 19924 30018
rect 19684 29996 19708 29998
rect 19764 29996 19788 29998
rect 19844 29996 19868 29998
rect 19706 29944 19708 29996
rect 19770 29944 19782 29996
rect 19844 29944 19846 29996
rect 19684 29942 19708 29944
rect 19764 29942 19788 29944
rect 19844 29942 19868 29944
rect 19628 29922 19924 29942
rect 19628 28666 19924 28686
rect 19684 28664 19708 28666
rect 19764 28664 19788 28666
rect 19844 28664 19868 28666
rect 19706 28612 19708 28664
rect 19770 28612 19782 28664
rect 19844 28612 19846 28664
rect 19684 28610 19708 28612
rect 19764 28610 19788 28612
rect 19844 28610 19868 28612
rect 19628 28590 19924 28610
rect 19628 27334 19924 27354
rect 19684 27332 19708 27334
rect 19764 27332 19788 27334
rect 19844 27332 19868 27334
rect 19706 27280 19708 27332
rect 19770 27280 19782 27332
rect 19844 27280 19846 27332
rect 19684 27278 19708 27280
rect 19764 27278 19788 27280
rect 19844 27278 19868 27280
rect 19628 27258 19924 27278
rect 19628 26002 19924 26022
rect 19684 26000 19708 26002
rect 19764 26000 19788 26002
rect 19844 26000 19868 26002
rect 19706 25948 19708 26000
rect 19770 25948 19782 26000
rect 19844 25948 19846 26000
rect 19684 25946 19708 25948
rect 19764 25946 19788 25948
rect 19844 25946 19868 25948
rect 19628 25926 19924 25946
rect 19628 24670 19924 24690
rect 19684 24668 19708 24670
rect 19764 24668 19788 24670
rect 19844 24668 19868 24670
rect 19706 24616 19708 24668
rect 19770 24616 19782 24668
rect 19844 24616 19846 24668
rect 19684 24614 19708 24616
rect 19764 24614 19788 24616
rect 19844 24614 19868 24616
rect 19628 24594 19924 24614
rect 19628 23338 19924 23358
rect 19684 23336 19708 23338
rect 19764 23336 19788 23338
rect 19844 23336 19868 23338
rect 19706 23284 19708 23336
rect 19770 23284 19782 23336
rect 19844 23284 19846 23336
rect 19684 23282 19708 23284
rect 19764 23282 19788 23284
rect 19844 23282 19868 23284
rect 19628 23262 19924 23282
rect 19628 22006 19924 22026
rect 19684 22004 19708 22006
rect 19764 22004 19788 22006
rect 19844 22004 19868 22006
rect 19706 21952 19708 22004
rect 19770 21952 19782 22004
rect 19844 21952 19846 22004
rect 19684 21950 19708 21952
rect 19764 21950 19788 21952
rect 19844 21950 19868 21952
rect 19628 21930 19924 21950
rect 19628 20674 19924 20694
rect 19684 20672 19708 20674
rect 19764 20672 19788 20674
rect 19844 20672 19868 20674
rect 19706 20620 19708 20672
rect 19770 20620 19782 20672
rect 19844 20620 19846 20672
rect 19684 20618 19708 20620
rect 19764 20618 19788 20620
rect 19844 20618 19868 20620
rect 19628 20598 19924 20618
rect 19628 19342 19924 19362
rect 19684 19340 19708 19342
rect 19764 19340 19788 19342
rect 19844 19340 19868 19342
rect 19706 19288 19708 19340
rect 19770 19288 19782 19340
rect 19844 19288 19846 19340
rect 19684 19286 19708 19288
rect 19764 19286 19788 19288
rect 19844 19286 19868 19288
rect 19628 19266 19924 19286
rect 19628 18010 19924 18030
rect 19684 18008 19708 18010
rect 19764 18008 19788 18010
rect 19844 18008 19868 18010
rect 19706 17956 19708 18008
rect 19770 17956 19782 18008
rect 19844 17956 19846 18008
rect 19684 17954 19708 17956
rect 19764 17954 19788 17956
rect 19844 17954 19868 17956
rect 19628 17934 19924 17954
rect 19628 16678 19924 16698
rect 19684 16676 19708 16678
rect 19764 16676 19788 16678
rect 19844 16676 19868 16678
rect 19706 16624 19708 16676
rect 19770 16624 19782 16676
rect 19844 16624 19846 16676
rect 19684 16622 19708 16624
rect 19764 16622 19788 16624
rect 19844 16622 19868 16624
rect 19628 16602 19924 16622
rect 19628 15346 19924 15366
rect 19684 15344 19708 15346
rect 19764 15344 19788 15346
rect 19844 15344 19868 15346
rect 19706 15292 19708 15344
rect 19770 15292 19782 15344
rect 19844 15292 19846 15344
rect 19684 15290 19708 15292
rect 19764 15290 19788 15292
rect 19844 15290 19868 15292
rect 19628 15270 19924 15290
rect 19628 14014 19924 14034
rect 19684 14012 19708 14014
rect 19764 14012 19788 14014
rect 19844 14012 19868 14014
rect 19706 13960 19708 14012
rect 19770 13960 19782 14012
rect 19844 13960 19846 14012
rect 19684 13958 19708 13960
rect 19764 13958 19788 13960
rect 19844 13958 19868 13960
rect 19628 13938 19924 13958
rect 19628 12682 19924 12702
rect 19684 12680 19708 12682
rect 19764 12680 19788 12682
rect 19844 12680 19868 12682
rect 19706 12628 19708 12680
rect 19770 12628 19782 12680
rect 19844 12628 19846 12680
rect 19684 12626 19708 12628
rect 19764 12626 19788 12628
rect 19844 12626 19868 12628
rect 19628 12606 19924 12626
rect 19628 11350 19924 11370
rect 19684 11348 19708 11350
rect 19764 11348 19788 11350
rect 19844 11348 19868 11350
rect 19706 11296 19708 11348
rect 19770 11296 19782 11348
rect 19844 11296 19846 11348
rect 19684 11294 19708 11296
rect 19764 11294 19788 11296
rect 19844 11294 19868 11296
rect 19628 11274 19924 11294
rect 19628 10018 19924 10038
rect 19684 10016 19708 10018
rect 19764 10016 19788 10018
rect 19844 10016 19868 10018
rect 19706 9964 19708 10016
rect 19770 9964 19782 10016
rect 19844 9964 19846 10016
rect 19684 9962 19708 9964
rect 19764 9962 19788 9964
rect 19844 9962 19868 9964
rect 19628 9942 19924 9962
rect 19318 9461 19370 9467
rect 19318 9403 19370 9409
rect 19628 8686 19924 8706
rect 19684 8684 19708 8686
rect 19764 8684 19788 8686
rect 19844 8684 19868 8686
rect 19706 8632 19708 8684
rect 19770 8632 19782 8684
rect 19844 8632 19846 8684
rect 19684 8630 19708 8632
rect 19764 8630 19788 8632
rect 19844 8630 19868 8632
rect 19628 8610 19924 8630
rect 19628 7354 19924 7374
rect 19684 7352 19708 7354
rect 19764 7352 19788 7354
rect 19844 7352 19868 7354
rect 19706 7300 19708 7352
rect 19770 7300 19782 7352
rect 19844 7300 19846 7352
rect 19684 7298 19708 7300
rect 19764 7298 19788 7300
rect 19844 7298 19868 7300
rect 19628 7278 19924 7298
rect 19222 6945 19274 6951
rect 19222 6887 19274 6893
rect 19030 6501 19082 6507
rect 19030 6443 19082 6449
rect 19604 6466 19660 6475
rect 20002 6433 20030 45145
rect 20386 15905 20414 55505
rect 20578 32555 20606 56171
rect 20566 32549 20618 32555
rect 20566 32491 20618 32497
rect 20470 28109 20522 28115
rect 20470 28051 20522 28057
rect 20374 15899 20426 15905
rect 20374 15841 20426 15847
rect 20482 7363 20510 28051
rect 20662 18341 20714 18347
rect 20662 18283 20714 18289
rect 20674 17294 20702 18283
rect 20578 17266 20702 17294
rect 20578 8431 20606 17266
rect 20866 9023 20894 56837
rect 21250 56531 21278 59200
rect 21730 56531 21758 59200
rect 22306 56975 22334 59200
rect 22294 56969 22346 56975
rect 22294 56911 22346 56917
rect 22294 56821 22346 56827
rect 22294 56763 22346 56769
rect 21238 56525 21290 56531
rect 21238 56467 21290 56473
rect 21718 56525 21770 56531
rect 21718 56467 21770 56473
rect 21046 56229 21098 56235
rect 21046 56171 21098 56177
rect 20950 9239 21002 9245
rect 20950 9181 21002 9187
rect 20854 9017 20906 9023
rect 20854 8959 20906 8965
rect 20566 8425 20618 8431
rect 20566 8367 20618 8373
rect 20962 7765 20990 9181
rect 20950 7759 21002 7765
rect 20950 7701 21002 7707
rect 21058 7691 21086 56171
rect 21334 44907 21386 44913
rect 21334 44849 21386 44855
rect 21046 7685 21098 7691
rect 21046 7627 21098 7633
rect 20758 7463 20810 7469
rect 20758 7405 20810 7411
rect 20468 7354 20524 7363
rect 20468 7289 20524 7298
rect 20470 7167 20522 7173
rect 20470 7109 20522 7115
rect 20182 7093 20234 7099
rect 20482 7044 20510 7109
rect 20234 7041 20510 7044
rect 20182 7035 20510 7041
rect 20194 7016 20510 7035
rect 20482 6951 20510 7016
rect 20086 6945 20138 6951
rect 20086 6887 20138 6893
rect 20278 6945 20330 6951
rect 20470 6945 20522 6951
rect 20330 6905 20414 6933
rect 20278 6887 20330 6893
rect 20098 6433 20126 6887
rect 19604 6401 19606 6410
rect 19658 6401 19660 6410
rect 19990 6427 20042 6433
rect 19606 6369 19658 6375
rect 19990 6369 20042 6375
rect 20086 6427 20138 6433
rect 20086 6369 20138 6375
rect 19318 6353 19370 6359
rect 19318 6295 19370 6301
rect 18742 5687 18794 5693
rect 18742 5629 18794 5635
rect 18754 800 18782 5629
rect 19030 5021 19082 5027
rect 19030 4963 19082 4969
rect 19126 5021 19178 5027
rect 19126 4963 19178 4969
rect 19042 3917 19070 4963
rect 19030 3911 19082 3917
rect 19030 3853 19082 3859
rect 18934 3837 18986 3843
rect 18934 3779 18986 3785
rect 18946 3251 18974 3779
rect 19030 3541 19082 3547
rect 19030 3483 19082 3489
rect 18934 3245 18986 3251
rect 18934 3187 18986 3193
rect 18850 3029 18974 3048
rect 18850 3023 18986 3029
rect 18850 3020 18934 3023
rect 18850 800 18878 3020
rect 18934 2965 18986 2971
rect 19042 2894 19070 3483
rect 18946 2866 19070 2894
rect 18946 800 18974 2866
rect 19138 1272 19166 4963
rect 19220 4246 19276 4255
rect 19220 4181 19276 4190
rect 19234 3917 19262 4181
rect 19222 3911 19274 3917
rect 19222 3853 19274 3859
rect 19222 3689 19274 3695
rect 19222 3631 19274 3637
rect 19042 1244 19166 1272
rect 19042 800 19070 1244
rect 19234 800 19262 3631
rect 19330 800 19358 6295
rect 19510 6131 19562 6137
rect 19510 6073 19562 6079
rect 19414 3911 19466 3917
rect 19414 3853 19466 3859
rect 19426 800 19454 3853
rect 19522 3547 19550 6073
rect 19628 6022 19924 6042
rect 19684 6020 19708 6022
rect 19764 6020 19788 6022
rect 19844 6020 19868 6022
rect 19706 5968 19708 6020
rect 19770 5968 19782 6020
rect 19844 5968 19846 6020
rect 19684 5966 19708 5968
rect 19764 5966 19788 5968
rect 19844 5966 19868 5968
rect 19628 5946 19924 5966
rect 20182 5687 20234 5693
rect 20182 5629 20234 5635
rect 19628 4690 19924 4710
rect 19684 4688 19708 4690
rect 19764 4688 19788 4690
rect 19844 4688 19868 4690
rect 19706 4636 19708 4688
rect 19770 4636 19782 4688
rect 19844 4636 19846 4688
rect 19684 4634 19708 4636
rect 19764 4634 19788 4636
rect 19844 4634 19868 4636
rect 19628 4614 19924 4634
rect 19990 3689 20042 3695
rect 19990 3631 20042 3637
rect 19510 3541 19562 3547
rect 19510 3483 19562 3489
rect 19628 3358 19924 3378
rect 19684 3356 19708 3358
rect 19764 3356 19788 3358
rect 19844 3356 19868 3358
rect 19706 3304 19708 3356
rect 19770 3304 19782 3356
rect 19844 3304 19846 3356
rect 19684 3302 19708 3304
rect 19764 3302 19788 3304
rect 19844 3302 19868 3304
rect 19628 3282 19924 3302
rect 19702 3245 19754 3251
rect 19702 3187 19754 3193
rect 19510 3097 19562 3103
rect 19510 3039 19562 3045
rect 19522 2807 19550 3039
rect 19606 2949 19658 2955
rect 19606 2891 19658 2897
rect 19510 2801 19562 2807
rect 19510 2743 19562 2749
rect 19618 800 19646 2891
rect 19714 800 19742 3187
rect 19798 3171 19850 3177
rect 19798 3113 19850 3119
rect 19810 800 19838 3113
rect 20002 1864 20030 3631
rect 20194 3177 20222 5629
rect 20278 4355 20330 4361
rect 20278 4297 20330 4303
rect 20182 3171 20234 3177
rect 20182 3113 20234 3119
rect 20086 2801 20138 2807
rect 20086 2743 20138 2749
rect 19906 1836 20030 1864
rect 19906 800 19934 1836
rect 20098 800 20126 2743
rect 20182 2579 20234 2585
rect 20182 2521 20234 2527
rect 20194 800 20222 2521
rect 20290 800 20318 4297
rect 20386 3251 20414 6905
rect 20470 6887 20522 6893
rect 20470 6279 20522 6285
rect 20470 6221 20522 6227
rect 20566 6279 20618 6285
rect 20566 6221 20618 6227
rect 20482 5545 20510 6221
rect 20578 5841 20606 6221
rect 20566 5835 20618 5841
rect 20566 5777 20618 5783
rect 20566 5687 20618 5693
rect 20566 5629 20618 5635
rect 20470 5539 20522 5545
rect 20470 5481 20522 5487
rect 20470 5021 20522 5027
rect 20470 4963 20522 4969
rect 20482 3917 20510 4963
rect 20470 3911 20522 3917
rect 20470 3853 20522 3859
rect 20470 3763 20522 3769
rect 20470 3705 20522 3711
rect 20374 3245 20426 3251
rect 20374 3187 20426 3193
rect 20482 800 20510 3705
rect 20578 800 20606 5629
rect 20662 3689 20714 3695
rect 20662 3631 20714 3637
rect 20674 800 20702 3631
rect 20770 800 20798 7405
rect 20854 6945 20906 6951
rect 20854 6887 20906 6893
rect 20866 3769 20894 6887
rect 21346 6031 21374 44849
rect 21910 38765 21962 38771
rect 21910 38707 21962 38713
rect 21922 7099 21950 38707
rect 22306 11095 22334 56763
rect 22786 56531 22814 59200
rect 22774 56525 22826 56531
rect 22774 56467 22826 56473
rect 22870 56229 22922 56235
rect 22870 56171 22922 56177
rect 22678 29219 22730 29225
rect 22678 29161 22730 29167
rect 22294 11089 22346 11095
rect 22294 11031 22346 11037
rect 22690 7099 22718 29161
rect 22882 21751 22910 56171
rect 23362 55717 23390 59200
rect 23842 56975 23870 59200
rect 23830 56969 23882 56975
rect 23830 56911 23882 56917
rect 24418 56531 24446 59200
rect 24406 56525 24458 56531
rect 24406 56467 24458 56473
rect 24310 56229 24362 56235
rect 24310 56171 24362 56177
rect 23350 55711 23402 55717
rect 23350 55653 23402 55659
rect 23446 55563 23498 55569
rect 23446 55505 23498 55511
rect 22870 21745 22922 21751
rect 22870 21687 22922 21693
rect 22966 18785 23018 18791
rect 22966 18727 23018 18733
rect 21910 7093 21962 7099
rect 21910 7035 21962 7041
rect 22678 7093 22730 7099
rect 22678 7035 22730 7041
rect 21826 6979 22046 7007
rect 21826 6951 21854 6979
rect 21814 6945 21866 6951
rect 21814 6887 21866 6893
rect 21910 6945 21962 6951
rect 21910 6887 21962 6893
rect 21430 6131 21482 6137
rect 21430 6073 21482 6079
rect 21526 6131 21578 6137
rect 21526 6073 21578 6079
rect 21332 6022 21388 6031
rect 21332 5957 21388 5966
rect 20950 5021 21002 5027
rect 20950 4963 21002 4969
rect 20854 3763 20906 3769
rect 20854 3705 20906 3711
rect 20852 3506 20908 3515
rect 20852 3441 20854 3450
rect 20906 3441 20908 3450
rect 20854 3409 20906 3415
rect 20962 3344 20990 4963
rect 21046 4355 21098 4361
rect 21046 4297 21098 4303
rect 20866 3316 20990 3344
rect 20866 2585 20894 3316
rect 20950 3245 21002 3251
rect 20950 3187 21002 3193
rect 20854 2579 20906 2585
rect 20854 2521 20906 2527
rect 20962 800 20990 3187
rect 21058 800 21086 4297
rect 21238 4281 21290 4287
rect 21238 4223 21290 4229
rect 21140 3210 21196 3219
rect 21140 3145 21142 3154
rect 21194 3145 21196 3154
rect 21142 3113 21194 3119
rect 21142 2949 21194 2955
rect 21140 2914 21142 2923
rect 21194 2914 21196 2923
rect 21140 2849 21196 2858
rect 21250 2752 21278 4223
rect 21334 3911 21386 3917
rect 21334 3853 21386 3859
rect 21154 2724 21278 2752
rect 21154 800 21182 2724
rect 21346 2604 21374 3853
rect 21442 3177 21470 6073
rect 21430 3171 21482 3177
rect 21430 3113 21482 3119
rect 21430 3023 21482 3029
rect 21430 2965 21482 2971
rect 21250 2576 21374 2604
rect 21250 800 21278 2576
rect 21442 800 21470 2965
rect 21538 800 21566 6073
rect 21718 5687 21770 5693
rect 21718 5629 21770 5635
rect 21622 5613 21674 5619
rect 21622 5555 21674 5561
rect 21634 800 21662 5555
rect 21730 3251 21758 5629
rect 21814 4355 21866 4361
rect 21814 4297 21866 4303
rect 21718 3245 21770 3251
rect 21718 3187 21770 3193
rect 21826 800 21854 4297
rect 21922 800 21950 6887
rect 22018 4287 22046 6979
rect 22678 6945 22730 6951
rect 22594 6905 22678 6933
rect 22102 5021 22154 5027
rect 22102 4963 22154 4969
rect 22006 4281 22058 4287
rect 22006 4223 22058 4229
rect 22114 3917 22142 4963
rect 22294 4207 22346 4213
rect 22294 4149 22346 4155
rect 22102 3911 22154 3917
rect 22102 3853 22154 3859
rect 22102 3689 22154 3695
rect 22102 3631 22154 3637
rect 22006 3245 22058 3251
rect 22006 3187 22058 3193
rect 22018 800 22046 3187
rect 22114 800 22142 3631
rect 22306 800 22334 4149
rect 22390 3097 22442 3103
rect 22390 3039 22442 3045
rect 22402 800 22430 3039
rect 22486 2949 22538 2955
rect 22486 2891 22538 2897
rect 22498 800 22526 2891
rect 22594 800 22622 6905
rect 22678 6887 22730 6893
rect 22870 6797 22922 6803
rect 22870 6739 22922 6745
rect 22676 6466 22732 6475
rect 22676 6401 22732 6410
rect 22690 5735 22718 6401
rect 22774 6279 22826 6285
rect 22774 6221 22826 6227
rect 22676 5726 22732 5735
rect 22676 5661 22732 5670
rect 22786 4287 22814 6221
rect 22882 5767 22910 6739
rect 22978 6285 23006 18727
rect 23458 9911 23486 55505
rect 23638 46757 23690 46763
rect 23638 46699 23690 46705
rect 23446 9905 23498 9911
rect 23446 9847 23498 9853
rect 23062 8795 23114 8801
rect 23062 8737 23114 8743
rect 23074 7173 23102 8737
rect 23156 7354 23212 7363
rect 23156 7289 23212 7298
rect 23170 7173 23198 7289
rect 23062 7167 23114 7173
rect 23062 7109 23114 7115
rect 23158 7167 23210 7173
rect 23158 7109 23210 7115
rect 23542 6945 23594 6951
rect 23542 6887 23594 6893
rect 23350 6797 23402 6803
rect 23350 6739 23402 6745
rect 22966 6279 23018 6285
rect 22966 6221 23018 6227
rect 22966 6131 23018 6137
rect 22966 6073 23018 6079
rect 22870 5761 22922 5767
rect 22870 5703 22922 5709
rect 22774 4281 22826 4287
rect 22774 4223 22826 4229
rect 22978 4213 23006 6073
rect 23062 5687 23114 5693
rect 23062 5629 23114 5635
rect 22966 4207 23018 4213
rect 22966 4149 23018 4155
rect 23074 3788 23102 5629
rect 23158 4947 23210 4953
rect 23158 4889 23210 4895
rect 22786 3760 23102 3788
rect 22786 800 22814 3760
rect 22870 3689 22922 3695
rect 22870 3631 22922 3637
rect 22882 800 22910 3631
rect 22966 3171 23018 3177
rect 22966 3113 23018 3119
rect 22978 800 23006 3113
rect 23170 800 23198 4889
rect 23254 4355 23306 4361
rect 23254 4297 23306 4303
rect 23266 800 23294 4297
rect 23362 800 23390 6739
rect 23554 5767 23582 6887
rect 23650 6623 23678 46699
rect 24022 34251 24074 34257
rect 24022 34193 24074 34199
rect 24034 7765 24062 34193
rect 24322 26857 24350 56171
rect 24898 55717 24926 59200
rect 25474 56975 25502 59200
rect 25462 56969 25514 56975
rect 25462 56911 25514 56917
rect 25174 56895 25226 56901
rect 25174 56837 25226 56843
rect 24886 55711 24938 55717
rect 24886 55653 24938 55659
rect 25078 55563 25130 55569
rect 25078 55505 25130 55511
rect 25090 27597 25118 55505
rect 25078 27591 25130 27597
rect 25078 27533 25130 27539
rect 24310 26851 24362 26857
rect 24310 26793 24362 26799
rect 24214 26259 24266 26265
rect 24214 26201 24266 26207
rect 24226 8135 24254 26201
rect 24502 16935 24554 16941
rect 24502 16877 24554 16883
rect 24406 11607 24458 11613
rect 24406 11549 24458 11555
rect 24418 8135 24446 11549
rect 24214 8129 24266 8135
rect 24214 8071 24266 8077
rect 24406 8129 24458 8135
rect 24406 8071 24458 8077
rect 24022 7759 24074 7765
rect 24022 7701 24074 7707
rect 23734 7463 23786 7469
rect 23734 7405 23786 7411
rect 24118 7463 24170 7469
rect 24118 7405 24170 7411
rect 23636 6614 23692 6623
rect 23636 6549 23692 6558
rect 23542 5761 23594 5767
rect 23542 5703 23594 5709
rect 23446 5687 23498 5693
rect 23446 5629 23498 5635
rect 23458 800 23486 5629
rect 23542 5021 23594 5027
rect 23542 4963 23594 4969
rect 23554 3103 23582 4963
rect 23638 3689 23690 3695
rect 23638 3631 23690 3637
rect 23542 3097 23594 3103
rect 23542 3039 23594 3045
rect 23650 800 23678 3631
rect 23746 800 23774 7405
rect 23828 7354 23884 7363
rect 23828 7289 23884 7298
rect 23842 6877 23870 7289
rect 23926 7093 23978 7099
rect 23926 7035 23978 7041
rect 23830 6871 23882 6877
rect 23830 6813 23882 6819
rect 23830 3911 23882 3917
rect 23830 3853 23882 3859
rect 23842 800 23870 3853
rect 23938 2807 23966 7035
rect 24022 6575 24074 6581
rect 24022 6517 24074 6523
rect 24034 6327 24062 6517
rect 24020 6318 24076 6327
rect 24020 6253 24076 6262
rect 24022 4355 24074 4361
rect 24022 4297 24074 4303
rect 24034 3251 24062 4297
rect 24022 3245 24074 3251
rect 24022 3187 24074 3193
rect 24022 3023 24074 3029
rect 24022 2965 24074 2971
rect 23926 2801 23978 2807
rect 23926 2743 23978 2749
rect 24034 800 24062 2965
rect 24130 800 24158 7405
rect 24514 6433 24542 16877
rect 24694 14789 24746 14795
rect 24694 14731 24746 14737
rect 24706 7765 24734 14731
rect 25186 11687 25214 56837
rect 25558 56821 25610 56827
rect 25558 56763 25610 56769
rect 25270 54749 25322 54755
rect 25270 54691 25322 54697
rect 25174 11681 25226 11687
rect 25174 11623 25226 11629
rect 24694 7759 24746 7765
rect 24694 7701 24746 7707
rect 25282 7691 25310 54691
rect 25366 40763 25418 40769
rect 25366 40705 25418 40711
rect 25270 7685 25322 7691
rect 25270 7627 25322 7633
rect 24790 7463 24842 7469
rect 24790 7405 24842 7411
rect 24598 6945 24650 6951
rect 24598 6887 24650 6893
rect 24502 6427 24554 6433
rect 24502 6369 24554 6375
rect 24406 6279 24458 6285
rect 24406 6221 24458 6227
rect 24310 6131 24362 6137
rect 24310 6073 24362 6079
rect 24214 4281 24266 4287
rect 24214 4223 24266 4229
rect 24226 800 24254 4223
rect 24322 3177 24350 6073
rect 24418 4435 24446 6221
rect 24610 5749 24638 6887
rect 24514 5721 24638 5749
rect 24406 4429 24458 4435
rect 24406 4371 24458 4377
rect 24406 3689 24458 3695
rect 24406 3631 24458 3637
rect 24310 3171 24362 3177
rect 24310 3113 24362 3119
rect 24418 1864 24446 3631
rect 24322 1836 24446 1864
rect 24322 800 24350 1836
rect 24514 800 24542 5721
rect 24598 5687 24650 5693
rect 24598 5629 24650 5635
rect 24610 800 24638 5629
rect 24694 3615 24746 3621
rect 24694 3557 24746 3563
rect 24706 800 24734 3557
rect 24802 800 24830 7405
rect 25378 7173 25406 40705
rect 25462 30403 25514 30409
rect 25462 30345 25514 30351
rect 25474 7765 25502 30345
rect 25570 14203 25598 56763
rect 25954 56531 25982 59200
rect 26530 56531 26558 59200
rect 27010 56975 27038 59200
rect 26998 56969 27050 56975
rect 26998 56911 27050 56917
rect 27586 56531 27614 59200
rect 28066 56531 28094 59200
rect 28642 56975 28670 59200
rect 29122 57049 29150 59200
rect 29110 57043 29162 57049
rect 29110 56985 29162 56991
rect 28630 56969 28682 56975
rect 28630 56911 28682 56917
rect 29698 56531 29726 59200
rect 30178 56957 30206 59200
rect 30262 56969 30314 56975
rect 30178 56929 30262 56957
rect 30262 56911 30314 56917
rect 30070 56895 30122 56901
rect 30070 56837 30122 56843
rect 25942 56525 25994 56531
rect 25942 56467 25994 56473
rect 26518 56525 26570 56531
rect 26518 56467 26570 56473
rect 27574 56525 27626 56531
rect 27574 56467 27626 56473
rect 28054 56525 28106 56531
rect 28054 56467 28106 56473
rect 29686 56525 29738 56531
rect 29686 56467 29738 56473
rect 26518 56229 26570 56235
rect 26518 56171 26570 56177
rect 27670 56229 27722 56235
rect 27670 56171 27722 56177
rect 28150 56229 28202 56235
rect 28150 56171 28202 56177
rect 29302 56229 29354 56235
rect 29302 56171 29354 56177
rect 26134 40911 26186 40917
rect 26134 40853 26186 40859
rect 26146 17294 26174 40853
rect 26422 27887 26474 27893
rect 26422 27829 26474 27835
rect 25954 17266 26174 17294
rect 25558 14197 25610 14203
rect 25558 14139 25610 14145
rect 25654 8203 25706 8209
rect 25654 8145 25706 8151
rect 25666 7839 25694 8145
rect 25954 7913 25982 17266
rect 25942 7907 25994 7913
rect 25942 7849 25994 7855
rect 25654 7833 25706 7839
rect 26230 7833 26282 7839
rect 25654 7775 25706 7781
rect 25858 7781 26230 7784
rect 25858 7775 26282 7781
rect 25462 7759 25514 7765
rect 25462 7701 25514 7707
rect 25858 7756 26270 7775
rect 25654 7685 25706 7691
rect 25858 7636 25886 7756
rect 25706 7633 25886 7636
rect 25654 7627 25886 7633
rect 25666 7608 25886 7627
rect 25942 7463 25994 7469
rect 25942 7405 25994 7411
rect 25174 7167 25226 7173
rect 25174 7109 25226 7115
rect 25366 7167 25418 7173
rect 25366 7109 25418 7115
rect 25654 7167 25706 7173
rect 25654 7109 25706 7115
rect 25186 6507 25214 7109
rect 25666 6951 25694 7109
rect 25654 6945 25706 6951
rect 25654 6887 25706 6893
rect 25174 6501 25226 6507
rect 25174 6443 25226 6449
rect 25654 6353 25706 6359
rect 25654 6295 25706 6301
rect 25078 5021 25130 5027
rect 25078 4963 25130 4969
rect 25090 3917 25118 4963
rect 25462 4355 25514 4361
rect 25462 4297 25514 4303
rect 25366 4207 25418 4213
rect 25366 4149 25418 4155
rect 25078 3911 25130 3917
rect 25078 3853 25130 3859
rect 25174 3763 25226 3769
rect 25174 3705 25226 3711
rect 24982 3245 25034 3251
rect 24982 3187 25034 3193
rect 24994 800 25022 3187
rect 25078 2949 25130 2955
rect 25078 2891 25130 2897
rect 25090 800 25118 2891
rect 25186 800 25214 3705
rect 25378 800 25406 4149
rect 25474 800 25502 4297
rect 25558 4133 25610 4139
rect 25558 4075 25610 4081
rect 25570 800 25598 4075
rect 25666 800 25694 6295
rect 25846 5021 25898 5027
rect 25846 4963 25898 4969
rect 25858 4287 25886 4963
rect 25846 4281 25898 4287
rect 25846 4223 25898 4229
rect 25954 4139 25982 7405
rect 26434 7099 26462 27829
rect 26530 10947 26558 56171
rect 27094 20117 27146 20123
rect 27094 20059 27146 20065
rect 27106 11687 27134 20059
rect 27190 19599 27242 19605
rect 27190 19541 27242 19547
rect 27094 11681 27146 11687
rect 27094 11623 27146 11629
rect 26518 10941 26570 10947
rect 26518 10883 26570 10889
rect 27094 7611 27146 7617
rect 27094 7553 27146 7559
rect 26710 7463 26762 7469
rect 26710 7405 26762 7411
rect 26422 7093 26474 7099
rect 26422 7035 26474 7041
rect 26326 6945 26378 6951
rect 26326 6887 26378 6893
rect 26230 5687 26282 5693
rect 26230 5629 26282 5635
rect 26038 5613 26090 5619
rect 26038 5555 26090 5561
rect 25942 4133 25994 4139
rect 25942 4075 25994 4081
rect 25942 3911 25994 3917
rect 25942 3853 25994 3859
rect 25846 3541 25898 3547
rect 25846 3483 25898 3489
rect 25858 800 25886 3483
rect 25954 800 25982 3853
rect 26050 800 26078 5555
rect 26134 4355 26186 4361
rect 26134 4297 26186 4303
rect 26146 800 26174 4297
rect 26242 4213 26270 5629
rect 26230 4207 26282 4213
rect 26230 4149 26282 4155
rect 26338 3769 26366 6887
rect 26614 5021 26666 5027
rect 26614 4963 26666 4969
rect 26518 4355 26570 4361
rect 26518 4297 26570 4303
rect 26422 4133 26474 4139
rect 26422 4075 26474 4081
rect 26326 3763 26378 3769
rect 26326 3705 26378 3711
rect 26326 3467 26378 3473
rect 26326 3409 26378 3415
rect 26338 800 26366 3409
rect 26434 800 26462 4075
rect 26530 800 26558 4297
rect 26626 3251 26654 4963
rect 26614 3245 26666 3251
rect 26614 3187 26666 3193
rect 26722 800 26750 7405
rect 26902 7093 26954 7099
rect 26902 7035 26954 7041
rect 26806 6353 26858 6359
rect 26806 6295 26858 6301
rect 26818 800 26846 6295
rect 26914 3917 26942 7035
rect 27106 7025 27134 7553
rect 27202 7099 27230 19541
rect 27682 15609 27710 56171
rect 27670 15603 27722 15609
rect 27670 15545 27722 15551
rect 28162 11095 28190 56171
rect 28246 55563 28298 55569
rect 28246 55505 28298 55511
rect 28258 55051 28286 55505
rect 29014 55415 29066 55421
rect 29014 55357 29066 55363
rect 28246 55045 28298 55051
rect 28246 54987 28298 54993
rect 28822 49865 28874 49871
rect 28822 49807 28874 49813
rect 28246 33659 28298 33665
rect 28246 33601 28298 33607
rect 28258 33147 28286 33601
rect 28342 33511 28394 33517
rect 28342 33453 28394 33459
rect 28246 33141 28298 33147
rect 28246 33083 28298 33089
rect 28354 27374 28382 33453
rect 28258 27346 28382 27374
rect 28150 11089 28202 11095
rect 28150 11031 28202 11037
rect 28052 7946 28108 7955
rect 28052 7881 28108 7890
rect 28066 7363 28094 7881
rect 28150 7463 28202 7469
rect 28150 7405 28202 7411
rect 27284 7354 27340 7363
rect 27284 7289 27340 7298
rect 28052 7354 28108 7363
rect 28052 7289 28108 7298
rect 27298 7173 27326 7289
rect 27286 7167 27338 7173
rect 27286 7109 27338 7115
rect 27190 7093 27242 7099
rect 27190 7035 27242 7041
rect 27094 7019 27146 7025
rect 27094 6961 27146 6967
rect 27958 6945 28010 6951
rect 27682 6905 27958 6933
rect 26998 6871 27050 6877
rect 26998 6813 27050 6819
rect 26902 3911 26954 3917
rect 26902 3853 26954 3859
rect 26902 3023 26954 3029
rect 26902 2965 26954 2971
rect 26914 800 26942 2965
rect 27010 800 27038 6813
rect 27682 6507 27710 6905
rect 27958 6887 28010 6893
rect 27958 6575 28010 6581
rect 27958 6517 28010 6523
rect 27670 6501 27722 6507
rect 27670 6443 27722 6449
rect 27574 6131 27626 6137
rect 27574 6073 27626 6079
rect 27382 5687 27434 5693
rect 27382 5629 27434 5635
rect 27394 4269 27422 5629
rect 27202 4241 27422 4269
rect 27202 800 27230 4241
rect 27478 3911 27530 3917
rect 27478 3853 27530 3859
rect 27382 3763 27434 3769
rect 27382 3705 27434 3711
rect 27286 3689 27338 3695
rect 27286 3631 27338 3637
rect 27298 800 27326 3631
rect 27394 800 27422 3705
rect 27490 800 27518 3853
rect 27586 3473 27614 6073
rect 27862 5687 27914 5693
rect 27862 5629 27914 5635
rect 27574 3467 27626 3473
rect 27574 3409 27626 3415
rect 27574 2949 27626 2955
rect 27574 2891 27626 2897
rect 27586 1568 27614 2891
rect 27766 2801 27818 2807
rect 27766 2743 27818 2749
rect 27586 1540 27710 1568
rect 27682 800 27710 1540
rect 27778 800 27806 2743
rect 27874 800 27902 5629
rect 27970 2807 27998 6517
rect 28054 5021 28106 5027
rect 28054 4963 28106 4969
rect 28066 4139 28094 4963
rect 28054 4133 28106 4139
rect 28054 4075 28106 4081
rect 28054 3541 28106 3547
rect 28054 3483 28106 3489
rect 27958 2801 28010 2807
rect 27958 2743 28010 2749
rect 28066 800 28094 3483
rect 28162 800 28190 7405
rect 28258 6433 28286 27346
rect 28630 26777 28682 26783
rect 28630 26719 28682 26725
rect 28342 20931 28394 20937
rect 28342 20873 28394 20879
rect 28354 17294 28382 20873
rect 28354 17266 28478 17294
rect 28450 6623 28478 17266
rect 28642 9615 28670 26719
rect 28726 22263 28778 22269
rect 28726 22205 28778 22211
rect 28630 9609 28682 9615
rect 28630 9551 28682 9557
rect 28534 7685 28586 7691
rect 28534 7627 28586 7633
rect 28546 7543 28574 7627
rect 28534 7537 28586 7543
rect 28534 7479 28586 7485
rect 28738 7099 28766 22205
rect 28726 7093 28778 7099
rect 28726 7035 28778 7041
rect 28630 6945 28682 6951
rect 28630 6887 28682 6893
rect 28534 6797 28586 6803
rect 28534 6739 28586 6745
rect 28436 6614 28492 6623
rect 28436 6549 28492 6558
rect 28246 6427 28298 6433
rect 28246 6369 28298 6375
rect 28438 6131 28490 6137
rect 28438 6073 28490 6079
rect 28342 4355 28394 4361
rect 28342 4297 28394 4303
rect 28246 4133 28298 4139
rect 28246 4075 28298 4081
rect 28258 800 28286 4075
rect 28354 800 28382 4297
rect 28450 3769 28478 6073
rect 28438 3763 28490 3769
rect 28438 3705 28490 3711
rect 28546 800 28574 6739
rect 28642 6581 28670 6887
rect 28834 6581 28862 49807
rect 29026 8801 29054 55357
rect 29110 40097 29162 40103
rect 29110 40039 29162 40045
rect 29014 8795 29066 8801
rect 29014 8737 29066 8743
rect 29122 7913 29150 40039
rect 29314 11835 29342 56171
rect 29974 30329 30026 30335
rect 29974 30271 30026 30277
rect 29302 11829 29354 11835
rect 29302 11771 29354 11777
rect 29782 10941 29834 10947
rect 29782 10883 29834 10889
rect 29206 8573 29258 8579
rect 29206 8515 29258 8521
rect 29218 7913 29246 8515
rect 29794 8209 29822 10883
rect 29782 8203 29834 8209
rect 29782 8145 29834 8151
rect 29986 8135 30014 30271
rect 30082 12871 30110 56837
rect 30658 56531 30686 59200
rect 31234 56531 31262 59200
rect 31714 56975 31742 59200
rect 31702 56969 31754 56975
rect 31702 56911 31754 56917
rect 32290 56531 32318 59200
rect 32662 56895 32714 56901
rect 32662 56837 32714 56843
rect 30646 56525 30698 56531
rect 30646 56467 30698 56473
rect 31222 56525 31274 56531
rect 31222 56467 31274 56473
rect 32278 56525 32330 56531
rect 32278 56467 32330 56473
rect 30262 56303 30314 56309
rect 30262 56245 30314 56251
rect 30274 51721 30302 56245
rect 30934 56229 30986 56235
rect 30934 56171 30986 56177
rect 32470 56229 32522 56235
rect 32470 56171 32522 56177
rect 30262 51715 30314 51721
rect 30262 51657 30314 51663
rect 30646 39505 30698 39511
rect 30646 39447 30698 39453
rect 30166 24113 30218 24119
rect 30166 24055 30218 24061
rect 30070 12865 30122 12871
rect 30070 12807 30122 12813
rect 29302 8129 29354 8135
rect 29302 8071 29354 8077
rect 29974 8129 30026 8135
rect 29974 8071 30026 8077
rect 29110 7907 29162 7913
rect 29110 7849 29162 7855
rect 29206 7907 29258 7913
rect 29206 7849 29258 7855
rect 29314 7839 29342 8071
rect 29302 7833 29354 7839
rect 29302 7775 29354 7781
rect 30178 7765 30206 24055
rect 30166 7759 30218 7765
rect 30166 7701 30218 7707
rect 29686 7611 29738 7617
rect 29686 7553 29738 7559
rect 29206 7463 29258 7469
rect 29206 7405 29258 7411
rect 29590 7463 29642 7469
rect 29590 7405 29642 7411
rect 28630 6575 28682 6581
rect 28630 6517 28682 6523
rect 28822 6575 28874 6581
rect 29110 6575 29162 6581
rect 28874 6535 29054 6563
rect 28822 6517 28874 6523
rect 29026 6433 29054 6535
rect 29110 6517 29162 6523
rect 29014 6427 29066 6433
rect 29014 6369 29066 6375
rect 28822 5687 28874 5693
rect 28822 5629 28874 5635
rect 28834 4269 28862 5629
rect 29122 5545 29150 6517
rect 29110 5539 29162 5545
rect 29110 5481 29162 5487
rect 28918 5021 28970 5027
rect 28918 4963 28970 4969
rect 29014 5021 29066 5027
rect 29014 4963 29066 4969
rect 28642 4241 28862 4269
rect 28642 800 28670 4241
rect 28930 3917 28958 4963
rect 29026 4139 29054 4963
rect 29110 4355 29162 4361
rect 29110 4297 29162 4303
rect 29014 4133 29066 4139
rect 29014 4075 29066 4081
rect 28918 3911 28970 3917
rect 28918 3853 28970 3859
rect 29014 3911 29066 3917
rect 29014 3853 29066 3859
rect 28726 3763 28778 3769
rect 28726 3705 28778 3711
rect 28738 800 28766 3705
rect 28918 3467 28970 3473
rect 28918 3409 28970 3415
rect 28930 800 28958 3409
rect 29026 800 29054 3853
rect 29122 800 29150 4297
rect 29218 800 29246 7405
rect 29302 7241 29354 7247
rect 29494 7241 29546 7247
rect 29354 7189 29494 7192
rect 29302 7183 29546 7189
rect 29314 7164 29534 7183
rect 29302 4133 29354 4139
rect 29302 4075 29354 4081
rect 29314 2604 29342 4075
rect 29494 3615 29546 3621
rect 29494 3557 29546 3563
rect 29314 2576 29438 2604
rect 29410 800 29438 2576
rect 29506 800 29534 3557
rect 29602 800 29630 7405
rect 29698 7025 29726 7553
rect 29782 7093 29834 7099
rect 29782 7035 29834 7041
rect 29878 7093 29930 7099
rect 29878 7035 29930 7041
rect 29686 7019 29738 7025
rect 29686 6961 29738 6967
rect 29794 6803 29822 7035
rect 29782 6797 29834 6803
rect 29782 6739 29834 6745
rect 29686 6353 29738 6359
rect 29686 6295 29738 6301
rect 29698 800 29726 6295
rect 29782 6131 29834 6137
rect 29782 6073 29834 6079
rect 29794 3473 29822 6073
rect 29890 5767 29918 7035
rect 29974 6945 30026 6951
rect 29974 6887 30026 6893
rect 29878 5761 29930 5767
rect 29878 5703 29930 5709
rect 29782 3467 29834 3473
rect 29782 3409 29834 3415
rect 29878 3023 29930 3029
rect 29878 2965 29930 2971
rect 29890 800 29918 2965
rect 29986 800 30014 6887
rect 30070 6871 30122 6877
rect 30070 6813 30122 6819
rect 30082 5735 30110 6813
rect 30658 6433 30686 39447
rect 30946 20493 30974 56171
rect 31318 52159 31370 52165
rect 31318 52101 31370 52107
rect 31030 35731 31082 35737
rect 31030 35673 31082 35679
rect 30934 20487 30986 20493
rect 30934 20429 30986 20435
rect 30836 8094 30892 8103
rect 30836 8029 30892 8038
rect 30850 7765 30878 8029
rect 30838 7759 30890 7765
rect 30838 7701 30890 7707
rect 30742 7167 30794 7173
rect 30742 7109 30794 7115
rect 30754 6433 30782 7109
rect 31042 7099 31070 35673
rect 31222 32105 31274 32111
rect 31222 32047 31274 32053
rect 31234 8579 31262 32047
rect 31222 8573 31274 8579
rect 31222 8515 31274 8521
rect 31126 7463 31178 7469
rect 31126 7405 31178 7411
rect 31030 7093 31082 7099
rect 31030 7035 31082 7041
rect 30646 6427 30698 6433
rect 30646 6369 30698 6375
rect 30742 6427 30794 6433
rect 30742 6369 30794 6375
rect 30646 6131 30698 6137
rect 30646 6073 30698 6079
rect 30068 5726 30124 5735
rect 30068 5661 30124 5670
rect 30262 5687 30314 5693
rect 30262 5629 30314 5635
rect 30274 2894 30302 5629
rect 30358 5021 30410 5027
rect 30358 4963 30410 4969
rect 30454 5021 30506 5027
rect 30454 4963 30506 4969
rect 30370 3917 30398 4963
rect 30466 4139 30494 4963
rect 30454 4133 30506 4139
rect 30454 4075 30506 4081
rect 30358 3911 30410 3917
rect 30358 3853 30410 3859
rect 30454 3689 30506 3695
rect 30082 2866 30302 2894
rect 30370 3649 30454 3677
rect 30082 800 30110 2866
rect 30370 1864 30398 3649
rect 30454 3631 30506 3637
rect 30454 3541 30506 3547
rect 30454 3483 30506 3489
rect 30274 1836 30398 1864
rect 30274 800 30302 1836
rect 30358 1765 30410 1771
rect 30358 1707 30410 1713
rect 30370 800 30398 1707
rect 30466 800 30494 3483
rect 30550 2949 30602 2955
rect 30550 2891 30602 2897
rect 30562 800 30590 2891
rect 30658 1771 30686 6073
rect 30838 5687 30890 5693
rect 30838 5629 30890 5635
rect 30742 3911 30794 3917
rect 30742 3853 30794 3859
rect 30646 1765 30698 1771
rect 30646 1707 30698 1713
rect 30754 800 30782 3853
rect 30850 800 30878 5629
rect 30934 4355 30986 4361
rect 30934 4297 30986 4303
rect 30946 800 30974 4297
rect 31138 2894 31166 7405
rect 31330 7173 31358 52101
rect 32086 48977 32138 48983
rect 32086 48919 32138 48925
rect 31702 10793 31754 10799
rect 31702 10735 31754 10741
rect 31318 7167 31370 7173
rect 31318 7109 31370 7115
rect 31510 7093 31562 7099
rect 31714 7081 31742 10735
rect 31562 7053 31742 7081
rect 31510 7035 31562 7041
rect 31990 6945 32042 6951
rect 31990 6887 32042 6893
rect 31222 6353 31274 6359
rect 31222 6295 31274 6301
rect 31042 2866 31166 2894
rect 31042 800 31070 2866
rect 31234 800 31262 6295
rect 31702 5687 31754 5693
rect 31702 5629 31754 5635
rect 31714 4528 31742 5629
rect 31894 5021 31946 5027
rect 31894 4963 31946 4969
rect 31618 4500 31742 4528
rect 31414 4207 31466 4213
rect 31414 4149 31466 4155
rect 31318 3689 31370 3695
rect 31318 3631 31370 3637
rect 31330 800 31358 3631
rect 31426 800 31454 4149
rect 31618 800 31646 4500
rect 31702 4355 31754 4361
rect 31702 4297 31754 4303
rect 31714 800 31742 4297
rect 31798 4133 31850 4139
rect 31798 4075 31850 4081
rect 31810 800 31838 4075
rect 31906 3547 31934 4963
rect 32002 3917 32030 6887
rect 32098 6433 32126 48919
rect 32482 39585 32510 56171
rect 32674 49057 32702 56837
rect 32770 56161 32798 59200
rect 33346 56975 33374 59200
rect 33334 56969 33386 56975
rect 33334 56911 33386 56917
rect 33826 56531 33854 59200
rect 34402 57614 34430 59200
rect 34402 57586 34622 57614
rect 34594 56531 34622 57586
rect 34882 56975 34910 59200
rect 34988 57304 35284 57324
rect 35044 57302 35068 57304
rect 35124 57302 35148 57304
rect 35204 57302 35228 57304
rect 35066 57250 35068 57302
rect 35130 57250 35142 57302
rect 35204 57250 35206 57302
rect 35044 57248 35068 57250
rect 35124 57248 35148 57250
rect 35204 57248 35228 57250
rect 34988 57228 35284 57248
rect 34870 56969 34922 56975
rect 34870 56911 34922 56917
rect 35458 56531 35486 59200
rect 35938 57614 35966 59200
rect 35938 57586 36254 57614
rect 36226 56531 36254 57586
rect 36514 56901 36542 59200
rect 36994 57614 37022 59200
rect 36994 57586 37118 57614
rect 36502 56895 36554 56901
rect 36502 56837 36554 56843
rect 36694 56747 36746 56753
rect 36694 56689 36746 56695
rect 33814 56525 33866 56531
rect 33814 56467 33866 56473
rect 34582 56525 34634 56531
rect 34582 56467 34634 56473
rect 35446 56525 35498 56531
rect 35446 56467 35498 56473
rect 36214 56525 36266 56531
rect 36214 56467 36266 56473
rect 33046 56229 33098 56235
rect 33046 56171 33098 56177
rect 34390 56229 34442 56235
rect 34390 56171 34442 56177
rect 36214 56229 36266 56235
rect 36214 56171 36266 56177
rect 36598 56229 36650 56235
rect 36598 56171 36650 56177
rect 32758 56155 32810 56161
rect 32758 56097 32810 56103
rect 32662 49051 32714 49057
rect 32662 48993 32714 48999
rect 32662 42539 32714 42545
rect 32662 42481 32714 42487
rect 32470 39579 32522 39585
rect 32470 39521 32522 39527
rect 32278 8943 32330 8949
rect 32278 8885 32330 8891
rect 32290 6581 32318 8885
rect 32674 7099 32702 42481
rect 32758 34769 32810 34775
rect 32758 34711 32810 34717
rect 32662 7093 32714 7099
rect 32662 7035 32714 7041
rect 32374 6945 32426 6951
rect 32374 6887 32426 6893
rect 32470 6945 32522 6951
rect 32470 6887 32522 6893
rect 32278 6575 32330 6581
rect 32278 6517 32330 6523
rect 32086 6427 32138 6433
rect 32086 6369 32138 6375
rect 32386 4213 32414 6887
rect 32374 4207 32426 4213
rect 32374 4149 32426 4155
rect 32482 4084 32510 6887
rect 32770 6327 32798 34711
rect 33058 13167 33086 56171
rect 33526 35583 33578 35589
rect 33526 35525 33578 35531
rect 33046 13161 33098 13167
rect 33046 13103 33098 13109
rect 32950 8129 33002 8135
rect 32950 8071 33002 8077
rect 33238 8129 33290 8135
rect 33238 8071 33290 8077
rect 32854 7167 32906 7173
rect 32854 7109 32906 7115
rect 32866 6623 32894 7109
rect 32852 6614 32908 6623
rect 32852 6549 32908 6558
rect 32756 6318 32812 6327
rect 32756 6253 32812 6262
rect 32962 5767 32990 8071
rect 33250 6803 33278 8071
rect 33238 6797 33290 6803
rect 33044 6762 33100 6771
rect 33238 6739 33290 6745
rect 33044 6697 33100 6706
rect 33058 6327 33086 6697
rect 33140 6614 33196 6623
rect 33538 6581 33566 35525
rect 34402 18495 34430 56171
rect 34988 55972 35284 55992
rect 35044 55970 35068 55972
rect 35124 55970 35148 55972
rect 35204 55970 35228 55972
rect 35066 55918 35068 55970
rect 35130 55918 35142 55970
rect 35204 55918 35206 55970
rect 35044 55916 35068 55918
rect 35124 55916 35148 55918
rect 35204 55916 35228 55918
rect 34988 55896 35284 55916
rect 35350 55119 35402 55125
rect 35350 55061 35402 55067
rect 34988 54640 35284 54660
rect 35044 54638 35068 54640
rect 35124 54638 35148 54640
rect 35204 54638 35228 54640
rect 35066 54586 35068 54638
rect 35130 54586 35142 54638
rect 35204 54586 35206 54638
rect 35044 54584 35068 54586
rect 35124 54584 35148 54586
rect 35204 54584 35228 54586
rect 34988 54564 35284 54584
rect 34988 53308 35284 53328
rect 35044 53306 35068 53308
rect 35124 53306 35148 53308
rect 35204 53306 35228 53308
rect 35066 53254 35068 53306
rect 35130 53254 35142 53306
rect 35204 53254 35206 53306
rect 35044 53252 35068 53254
rect 35124 53252 35148 53254
rect 35204 53252 35228 53254
rect 34988 53232 35284 53252
rect 34988 51976 35284 51996
rect 35044 51974 35068 51976
rect 35124 51974 35148 51976
rect 35204 51974 35228 51976
rect 35066 51922 35068 51974
rect 35130 51922 35142 51974
rect 35204 51922 35206 51974
rect 35044 51920 35068 51922
rect 35124 51920 35148 51922
rect 35204 51920 35228 51922
rect 34988 51900 35284 51920
rect 34988 50644 35284 50664
rect 35044 50642 35068 50644
rect 35124 50642 35148 50644
rect 35204 50642 35228 50644
rect 35066 50590 35068 50642
rect 35130 50590 35142 50642
rect 35204 50590 35206 50642
rect 35044 50588 35068 50590
rect 35124 50588 35148 50590
rect 35204 50588 35228 50590
rect 34988 50568 35284 50588
rect 34988 49312 35284 49332
rect 35044 49310 35068 49312
rect 35124 49310 35148 49312
rect 35204 49310 35228 49312
rect 35066 49258 35068 49310
rect 35130 49258 35142 49310
rect 35204 49258 35206 49310
rect 35044 49256 35068 49258
rect 35124 49256 35148 49258
rect 35204 49256 35228 49258
rect 34988 49236 35284 49256
rect 34988 47980 35284 48000
rect 35044 47978 35068 47980
rect 35124 47978 35148 47980
rect 35204 47978 35228 47980
rect 35066 47926 35068 47978
rect 35130 47926 35142 47978
rect 35204 47926 35206 47978
rect 35044 47924 35068 47926
rect 35124 47924 35148 47926
rect 35204 47924 35228 47926
rect 34988 47904 35284 47924
rect 34582 47571 34634 47577
rect 34582 47513 34634 47519
rect 34390 18489 34442 18495
rect 34390 18431 34442 18437
rect 34294 10867 34346 10873
rect 34294 10809 34346 10815
rect 33814 10571 33866 10577
rect 33814 10513 33866 10519
rect 33826 7617 33854 10513
rect 33814 7611 33866 7617
rect 33814 7553 33866 7559
rect 33622 7463 33674 7469
rect 33622 7405 33674 7411
rect 33140 6549 33196 6558
rect 33526 6575 33578 6581
rect 33044 6318 33100 6327
rect 33044 6253 33100 6262
rect 33154 6211 33182 6549
rect 33526 6517 33578 6523
rect 33250 6276 33470 6304
rect 33142 6205 33194 6211
rect 33142 6147 33194 6153
rect 33250 6008 33278 6276
rect 33334 6205 33386 6211
rect 33334 6147 33386 6153
rect 33058 5980 33278 6008
rect 32950 5761 33002 5767
rect 32950 5703 33002 5709
rect 32950 4503 33002 4509
rect 32950 4445 33002 4451
rect 32758 4355 32810 4361
rect 32758 4297 32810 4303
rect 32194 4056 32510 4084
rect 31990 3911 32042 3917
rect 31990 3853 32042 3859
rect 31894 3541 31946 3547
rect 31894 3483 31946 3489
rect 31894 3097 31946 3103
rect 31894 3039 31946 3045
rect 31906 800 31934 3039
rect 32086 3023 32138 3029
rect 32086 2965 32138 2971
rect 32098 800 32126 2965
rect 32194 800 32222 4056
rect 32470 3689 32522 3695
rect 32470 3631 32522 3637
rect 32278 2949 32330 2955
rect 32278 2891 32330 2897
rect 32290 800 32318 2891
rect 32482 800 32510 3631
rect 32566 3467 32618 3473
rect 32566 3409 32618 3415
rect 32578 800 32606 3409
rect 32662 3245 32714 3251
rect 32662 3187 32714 3193
rect 32674 800 32702 3187
rect 32770 800 32798 4297
rect 32962 800 32990 4445
rect 33058 4139 33086 5980
rect 33346 5860 33374 6147
rect 33442 6137 33470 6276
rect 33430 6131 33482 6137
rect 33430 6073 33482 6079
rect 33154 5841 33374 5860
rect 33142 5835 33374 5841
rect 33194 5832 33374 5835
rect 33142 5777 33194 5783
rect 33142 5687 33194 5693
rect 33142 5629 33194 5635
rect 33046 4133 33098 4139
rect 33046 4075 33098 4081
rect 33154 2955 33182 5629
rect 33238 5613 33290 5619
rect 33238 5555 33290 5561
rect 33142 2949 33194 2955
rect 33142 2891 33194 2897
rect 33250 2752 33278 5555
rect 33334 5021 33386 5027
rect 33334 4963 33386 4969
rect 33346 3103 33374 4963
rect 33430 3911 33482 3917
rect 33430 3853 33482 3859
rect 33334 3097 33386 3103
rect 33334 3039 33386 3045
rect 33334 2949 33386 2955
rect 33334 2891 33386 2897
rect 33058 2724 33278 2752
rect 33058 800 33086 2724
rect 33346 1420 33374 2891
rect 33154 1392 33374 1420
rect 33154 800 33182 1392
rect 33238 1321 33290 1327
rect 33238 1263 33290 1269
rect 33250 800 33278 1263
rect 33442 800 33470 3853
rect 33526 3689 33578 3695
rect 33526 3631 33578 3637
rect 33538 800 33566 3631
rect 33634 800 33662 7405
rect 33910 6945 33962 6951
rect 33910 6887 33962 6893
rect 34102 6945 34154 6951
rect 34102 6887 34154 6893
rect 34198 6945 34250 6951
rect 34198 6887 34250 6893
rect 33814 6871 33866 6877
rect 33814 6813 33866 6819
rect 33826 6771 33854 6813
rect 33812 6762 33868 6771
rect 33812 6697 33868 6706
rect 33718 6131 33770 6137
rect 33718 6073 33770 6079
rect 33730 3473 33758 6073
rect 33922 4509 33950 6887
rect 34114 6803 34142 6887
rect 34102 6797 34154 6803
rect 34102 6739 34154 6745
rect 34210 5120 34238 6887
rect 34306 6433 34334 10809
rect 34594 7765 34622 47513
rect 34988 46648 35284 46668
rect 35044 46646 35068 46648
rect 35124 46646 35148 46648
rect 35204 46646 35228 46648
rect 35066 46594 35068 46646
rect 35130 46594 35142 46646
rect 35204 46594 35206 46646
rect 35044 46592 35068 46594
rect 35124 46592 35148 46594
rect 35204 46592 35228 46594
rect 34988 46572 35284 46592
rect 35362 45727 35390 55061
rect 35350 45721 35402 45727
rect 35350 45663 35402 45669
rect 34988 45316 35284 45336
rect 35044 45314 35068 45316
rect 35124 45314 35148 45316
rect 35204 45314 35228 45316
rect 35066 45262 35068 45314
rect 35130 45262 35142 45314
rect 35204 45262 35206 45314
rect 35044 45260 35068 45262
rect 35124 45260 35148 45262
rect 35204 45260 35228 45262
rect 34988 45240 35284 45260
rect 34988 43984 35284 44004
rect 35044 43982 35068 43984
rect 35124 43982 35148 43984
rect 35204 43982 35228 43984
rect 35066 43930 35068 43982
rect 35130 43930 35142 43982
rect 35204 43930 35206 43982
rect 35044 43928 35068 43930
rect 35124 43928 35148 43930
rect 35204 43928 35228 43930
rect 34988 43908 35284 43928
rect 34988 42652 35284 42672
rect 35044 42650 35068 42652
rect 35124 42650 35148 42652
rect 35204 42650 35228 42652
rect 35066 42598 35068 42650
rect 35130 42598 35142 42650
rect 35204 42598 35206 42650
rect 35044 42596 35068 42598
rect 35124 42596 35148 42598
rect 35204 42596 35228 42598
rect 34988 42576 35284 42596
rect 34988 41320 35284 41340
rect 35044 41318 35068 41320
rect 35124 41318 35148 41320
rect 35204 41318 35228 41320
rect 35066 41266 35068 41318
rect 35130 41266 35142 41318
rect 35204 41266 35206 41318
rect 35044 41264 35068 41266
rect 35124 41264 35148 41266
rect 35204 41264 35228 41266
rect 34988 41244 35284 41264
rect 34988 39988 35284 40008
rect 35044 39986 35068 39988
rect 35124 39986 35148 39988
rect 35204 39986 35228 39988
rect 35066 39934 35068 39986
rect 35130 39934 35142 39986
rect 35204 39934 35206 39986
rect 35044 39932 35068 39934
rect 35124 39932 35148 39934
rect 35204 39932 35228 39934
rect 34988 39912 35284 39932
rect 34988 38656 35284 38676
rect 35044 38654 35068 38656
rect 35124 38654 35148 38656
rect 35204 38654 35228 38656
rect 35066 38602 35068 38654
rect 35130 38602 35142 38654
rect 35204 38602 35206 38654
rect 35044 38600 35068 38602
rect 35124 38600 35148 38602
rect 35204 38600 35228 38602
rect 34988 38580 35284 38600
rect 34988 37324 35284 37344
rect 35044 37322 35068 37324
rect 35124 37322 35148 37324
rect 35204 37322 35228 37324
rect 35066 37270 35068 37322
rect 35130 37270 35142 37322
rect 35204 37270 35206 37322
rect 35044 37268 35068 37270
rect 35124 37268 35148 37270
rect 35204 37268 35228 37270
rect 34988 37248 35284 37268
rect 34988 35992 35284 36012
rect 35044 35990 35068 35992
rect 35124 35990 35148 35992
rect 35204 35990 35228 35992
rect 35066 35938 35068 35990
rect 35130 35938 35142 35990
rect 35204 35938 35206 35990
rect 35044 35936 35068 35938
rect 35124 35936 35148 35938
rect 35204 35936 35228 35938
rect 34988 35916 35284 35936
rect 34988 34660 35284 34680
rect 35044 34658 35068 34660
rect 35124 34658 35148 34660
rect 35204 34658 35228 34660
rect 35066 34606 35068 34658
rect 35130 34606 35142 34658
rect 35204 34606 35206 34658
rect 35044 34604 35068 34606
rect 35124 34604 35148 34606
rect 35204 34604 35228 34606
rect 34988 34584 35284 34604
rect 34988 33328 35284 33348
rect 35044 33326 35068 33328
rect 35124 33326 35148 33328
rect 35204 33326 35228 33328
rect 35066 33274 35068 33326
rect 35130 33274 35142 33326
rect 35204 33274 35206 33326
rect 35044 33272 35068 33274
rect 35124 33272 35148 33274
rect 35204 33272 35228 33274
rect 34988 33252 35284 33272
rect 34774 32105 34826 32111
rect 34774 32047 34826 32053
rect 34582 7759 34634 7765
rect 34582 7701 34634 7707
rect 34390 7463 34442 7469
rect 34390 7405 34442 7411
rect 34294 6427 34346 6433
rect 34294 6369 34346 6375
rect 34294 6131 34346 6137
rect 34294 6073 34346 6079
rect 34018 5092 34238 5120
rect 33910 4503 33962 4509
rect 33910 4445 33962 4451
rect 33910 4355 33962 4361
rect 33910 4297 33962 4303
rect 33814 4133 33866 4139
rect 33814 4075 33866 4081
rect 33718 3467 33770 3473
rect 33718 3409 33770 3415
rect 33716 3358 33772 3367
rect 33716 3293 33772 3302
rect 33730 1327 33758 3293
rect 33718 1321 33770 1327
rect 33718 1263 33770 1269
rect 33826 800 33854 4075
rect 33922 800 33950 4297
rect 34018 800 34046 5092
rect 34102 5021 34154 5027
rect 34102 4963 34154 4969
rect 34114 3251 34142 4963
rect 34198 4281 34250 4287
rect 34198 4223 34250 4229
rect 34102 3245 34154 3251
rect 34102 3187 34154 3193
rect 34210 2894 34238 4223
rect 34306 3811 34334 6073
rect 34292 3802 34348 3811
rect 34292 3737 34348 3746
rect 34294 3689 34346 3695
rect 34294 3631 34346 3637
rect 34114 2866 34238 2894
rect 34114 800 34142 2866
rect 34306 800 34334 3631
rect 34402 800 34430 7405
rect 34786 7099 34814 32047
rect 34988 31996 35284 32016
rect 35044 31994 35068 31996
rect 35124 31994 35148 31996
rect 35204 31994 35228 31996
rect 35066 31942 35068 31994
rect 35130 31942 35142 31994
rect 35204 31942 35206 31994
rect 35044 31940 35068 31942
rect 35124 31940 35148 31942
rect 35204 31940 35228 31942
rect 34988 31920 35284 31940
rect 34988 30664 35284 30684
rect 35044 30662 35068 30664
rect 35124 30662 35148 30664
rect 35204 30662 35228 30664
rect 35066 30610 35068 30662
rect 35130 30610 35142 30662
rect 35204 30610 35206 30662
rect 35044 30608 35068 30610
rect 35124 30608 35148 30610
rect 35204 30608 35228 30610
rect 34988 30588 35284 30608
rect 34988 29332 35284 29352
rect 35044 29330 35068 29332
rect 35124 29330 35148 29332
rect 35204 29330 35228 29332
rect 35066 29278 35068 29330
rect 35130 29278 35142 29330
rect 35204 29278 35206 29330
rect 35044 29276 35068 29278
rect 35124 29276 35148 29278
rect 35204 29276 35228 29278
rect 34988 29256 35284 29276
rect 34988 28000 35284 28020
rect 35044 27998 35068 28000
rect 35124 27998 35148 28000
rect 35204 27998 35228 28000
rect 35066 27946 35068 27998
rect 35130 27946 35142 27998
rect 35204 27946 35206 27998
rect 35044 27944 35068 27946
rect 35124 27944 35148 27946
rect 35204 27944 35228 27946
rect 34988 27924 35284 27944
rect 34988 26668 35284 26688
rect 35044 26666 35068 26668
rect 35124 26666 35148 26668
rect 35204 26666 35228 26668
rect 35066 26614 35068 26666
rect 35130 26614 35142 26666
rect 35204 26614 35206 26666
rect 35044 26612 35068 26614
rect 35124 26612 35148 26614
rect 35204 26612 35228 26614
rect 34988 26592 35284 26612
rect 36118 26259 36170 26265
rect 36118 26201 36170 26207
rect 34988 25336 35284 25356
rect 35044 25334 35068 25336
rect 35124 25334 35148 25336
rect 35204 25334 35228 25336
rect 35066 25282 35068 25334
rect 35130 25282 35142 25334
rect 35204 25282 35206 25334
rect 35044 25280 35068 25282
rect 35124 25280 35148 25282
rect 35204 25280 35228 25282
rect 34988 25260 35284 25280
rect 34870 24187 34922 24193
rect 34870 24129 34922 24135
rect 34882 23897 34910 24129
rect 34988 24004 35284 24024
rect 35044 24002 35068 24004
rect 35124 24002 35148 24004
rect 35204 24002 35228 24004
rect 35066 23950 35068 24002
rect 35130 23950 35142 24002
rect 35204 23950 35206 24002
rect 35044 23948 35068 23950
rect 35124 23948 35148 23950
rect 35204 23948 35228 23950
rect 34988 23928 35284 23948
rect 34870 23891 34922 23897
rect 34870 23833 34922 23839
rect 34988 22672 35284 22692
rect 35044 22670 35068 22672
rect 35124 22670 35148 22672
rect 35204 22670 35228 22672
rect 35066 22618 35068 22670
rect 35130 22618 35142 22670
rect 35204 22618 35206 22670
rect 35044 22616 35068 22618
rect 35124 22616 35148 22618
rect 35204 22616 35228 22618
rect 34988 22596 35284 22616
rect 34870 22263 34922 22269
rect 34870 22205 34922 22211
rect 34882 7913 34910 22205
rect 34988 21340 35284 21360
rect 35044 21338 35068 21340
rect 35124 21338 35148 21340
rect 35204 21338 35228 21340
rect 35066 21286 35068 21338
rect 35130 21286 35142 21338
rect 35204 21286 35206 21338
rect 35044 21284 35068 21286
rect 35124 21284 35148 21286
rect 35204 21284 35228 21286
rect 34988 21264 35284 21284
rect 34988 20008 35284 20028
rect 35044 20006 35068 20008
rect 35124 20006 35148 20008
rect 35204 20006 35228 20008
rect 35066 19954 35068 20006
rect 35130 19954 35142 20006
rect 35204 19954 35206 20006
rect 35044 19952 35068 19954
rect 35124 19952 35148 19954
rect 35204 19952 35228 19954
rect 34988 19932 35284 19952
rect 34988 18676 35284 18696
rect 35044 18674 35068 18676
rect 35124 18674 35148 18676
rect 35204 18674 35228 18676
rect 35066 18622 35068 18674
rect 35130 18622 35142 18674
rect 35204 18622 35206 18674
rect 35044 18620 35068 18622
rect 35124 18620 35148 18622
rect 35204 18620 35228 18622
rect 34988 18600 35284 18620
rect 34988 17344 35284 17364
rect 35044 17342 35068 17344
rect 35124 17342 35148 17344
rect 35204 17342 35228 17344
rect 35066 17290 35068 17342
rect 35130 17290 35142 17342
rect 35204 17290 35206 17342
rect 35044 17288 35068 17290
rect 35124 17288 35148 17290
rect 35204 17288 35228 17290
rect 34988 17268 35284 17288
rect 34988 16012 35284 16032
rect 35044 16010 35068 16012
rect 35124 16010 35148 16012
rect 35204 16010 35228 16012
rect 35066 15958 35068 16010
rect 35130 15958 35142 16010
rect 35204 15958 35206 16010
rect 35044 15956 35068 15958
rect 35124 15956 35148 15958
rect 35204 15956 35228 15958
rect 34988 15936 35284 15956
rect 34988 14680 35284 14700
rect 35044 14678 35068 14680
rect 35124 14678 35148 14680
rect 35204 14678 35228 14680
rect 35066 14626 35068 14678
rect 35130 14626 35142 14678
rect 35204 14626 35206 14678
rect 35044 14624 35068 14626
rect 35124 14624 35148 14626
rect 35204 14624 35228 14626
rect 34988 14604 35284 14624
rect 34988 13348 35284 13368
rect 35044 13346 35068 13348
rect 35124 13346 35148 13348
rect 35204 13346 35228 13348
rect 35066 13294 35068 13346
rect 35130 13294 35142 13346
rect 35204 13294 35206 13346
rect 35044 13292 35068 13294
rect 35124 13292 35148 13294
rect 35204 13292 35228 13294
rect 34988 13272 35284 13292
rect 34988 12016 35284 12036
rect 35044 12014 35068 12016
rect 35124 12014 35148 12016
rect 35204 12014 35228 12016
rect 35066 11962 35068 12014
rect 35130 11962 35142 12014
rect 35204 11962 35206 12014
rect 35044 11960 35068 11962
rect 35124 11960 35148 11962
rect 35204 11960 35228 11962
rect 34988 11940 35284 11960
rect 34988 10684 35284 10704
rect 35044 10682 35068 10684
rect 35124 10682 35148 10684
rect 35204 10682 35228 10684
rect 35066 10630 35068 10682
rect 35130 10630 35142 10682
rect 35204 10630 35206 10682
rect 35044 10628 35068 10630
rect 35124 10628 35148 10630
rect 35204 10628 35228 10630
rect 34988 10608 35284 10628
rect 34988 9352 35284 9372
rect 35044 9350 35068 9352
rect 35124 9350 35148 9352
rect 35204 9350 35228 9352
rect 35066 9298 35068 9350
rect 35130 9298 35142 9350
rect 35204 9298 35206 9350
rect 35044 9296 35068 9298
rect 35124 9296 35148 9298
rect 35204 9296 35228 9298
rect 34988 9276 35284 9296
rect 34988 8020 35284 8040
rect 35044 8018 35068 8020
rect 35124 8018 35148 8020
rect 35204 8018 35228 8020
rect 35066 7966 35068 8018
rect 35130 7966 35142 8018
rect 35204 7966 35206 8018
rect 35044 7964 35068 7966
rect 35124 7964 35148 7966
rect 35204 7964 35228 7966
rect 34988 7944 35284 7964
rect 34870 7907 34922 7913
rect 34870 7849 34922 7855
rect 36130 7765 36158 26201
rect 36226 8801 36254 56171
rect 36610 14129 36638 56171
rect 36706 15239 36734 56689
rect 37090 56161 37118 57586
rect 37570 56531 37598 59200
rect 38050 56975 38078 59200
rect 38038 56969 38090 56975
rect 38038 56911 38090 56917
rect 38134 56969 38186 56975
rect 38134 56911 38186 56917
rect 37558 56525 37610 56531
rect 37558 56467 37610 56473
rect 37654 56229 37706 56235
rect 37654 56171 37706 56177
rect 37078 56155 37130 56161
rect 37078 56097 37130 56103
rect 37666 25451 37694 56171
rect 38146 52387 38174 56911
rect 38626 56531 38654 59200
rect 38614 56525 38666 56531
rect 38614 56467 38666 56473
rect 38614 56229 38666 56235
rect 38614 56171 38666 56177
rect 38134 52381 38186 52387
rect 38134 52323 38186 52329
rect 38626 38327 38654 56171
rect 39106 55717 39134 59200
rect 39478 57043 39530 57049
rect 39478 56985 39530 56991
rect 39490 56383 39518 56985
rect 39682 56901 39710 59200
rect 39670 56895 39722 56901
rect 39670 56837 39722 56843
rect 39766 56747 39818 56753
rect 39766 56689 39818 56695
rect 39478 56377 39530 56383
rect 39478 56319 39530 56325
rect 39574 56377 39626 56383
rect 39574 56319 39626 56325
rect 39094 55711 39146 55717
rect 39094 55653 39146 55659
rect 38806 55637 38858 55643
rect 38806 55579 38858 55585
rect 38818 45209 38846 55579
rect 38902 55415 38954 55421
rect 38902 55357 38954 55363
rect 38806 45203 38858 45209
rect 38806 45145 38858 45151
rect 38614 38321 38666 38327
rect 38614 38263 38666 38269
rect 38326 38099 38378 38105
rect 38326 38041 38378 38047
rect 37654 25445 37706 25451
rect 37654 25387 37706 25393
rect 36886 23595 36938 23601
rect 36886 23537 36938 23543
rect 36694 15233 36746 15239
rect 36694 15175 36746 15181
rect 36598 14123 36650 14129
rect 36598 14065 36650 14071
rect 36214 8795 36266 8801
rect 36214 8737 36266 8743
rect 36898 7765 36926 23537
rect 36982 22263 37034 22269
rect 36982 22205 37034 22211
rect 36118 7759 36170 7765
rect 36118 7701 36170 7707
rect 36886 7759 36938 7765
rect 36886 7701 36938 7707
rect 35254 7685 35306 7691
rect 35446 7685 35498 7691
rect 35306 7633 35446 7636
rect 35254 7627 35498 7633
rect 35158 7611 35210 7617
rect 35266 7608 35486 7627
rect 35542 7611 35594 7617
rect 35158 7553 35210 7559
rect 35542 7553 35594 7559
rect 35170 7525 35198 7553
rect 35554 7525 35582 7553
rect 35170 7497 35582 7525
rect 34870 7463 34922 7469
rect 34870 7405 34922 7411
rect 35830 7463 35882 7469
rect 35830 7405 35882 7411
rect 36598 7463 36650 7469
rect 36598 7405 36650 7411
rect 34774 7093 34826 7099
rect 34774 7035 34826 7041
rect 34486 7019 34538 7025
rect 34486 6961 34538 6967
rect 34498 6211 34526 6961
rect 34582 6871 34634 6877
rect 34582 6813 34634 6819
rect 34594 6771 34622 6813
rect 34580 6762 34636 6771
rect 34580 6697 34636 6706
rect 34676 6466 34732 6475
rect 34676 6401 34678 6410
rect 34730 6401 34732 6410
rect 34678 6369 34730 6375
rect 34486 6205 34538 6211
rect 34486 6147 34538 6153
rect 34678 5687 34730 5693
rect 34678 5629 34730 5635
rect 34582 4947 34634 4953
rect 34582 4889 34634 4895
rect 34594 4528 34622 4889
rect 34498 4500 34622 4528
rect 34498 800 34526 4500
rect 34582 4355 34634 4361
rect 34582 4297 34634 4303
rect 34594 800 34622 4297
rect 34690 4139 34718 5629
rect 34774 5021 34826 5027
rect 34774 4963 34826 4969
rect 34678 4133 34730 4139
rect 34678 4075 34730 4081
rect 34786 3917 34814 4963
rect 34774 3911 34826 3917
rect 34774 3853 34826 3859
rect 34678 3837 34730 3843
rect 34678 3779 34730 3785
rect 34690 1179 34718 3779
rect 34882 1420 34910 7405
rect 35542 6945 35594 6951
rect 35542 6887 35594 6893
rect 35446 6797 35498 6803
rect 35444 6762 35446 6771
rect 35498 6762 35500 6771
rect 34988 6688 35284 6708
rect 35444 6697 35500 6706
rect 35044 6686 35068 6688
rect 35124 6686 35148 6688
rect 35204 6686 35228 6688
rect 35066 6634 35068 6686
rect 35130 6634 35142 6686
rect 35204 6634 35206 6686
rect 35044 6632 35068 6634
rect 35124 6632 35148 6634
rect 35204 6632 35228 6634
rect 34988 6612 35284 6632
rect 35446 6131 35498 6137
rect 35446 6073 35498 6079
rect 34988 5356 35284 5376
rect 35044 5354 35068 5356
rect 35124 5354 35148 5356
rect 35204 5354 35228 5356
rect 35066 5302 35068 5354
rect 35130 5302 35142 5354
rect 35204 5302 35206 5354
rect 35044 5300 35068 5302
rect 35124 5300 35148 5302
rect 35204 5300 35228 5302
rect 34988 5280 35284 5300
rect 34988 4024 35284 4044
rect 35044 4022 35068 4024
rect 35124 4022 35148 4024
rect 35204 4022 35228 4024
rect 35066 3970 35068 4022
rect 35130 3970 35142 4022
rect 35204 3970 35206 4022
rect 35044 3968 35068 3970
rect 35124 3968 35148 3970
rect 35204 3968 35228 3970
rect 34988 3948 35284 3968
rect 35458 3843 35486 6073
rect 35446 3837 35498 3843
rect 35446 3779 35498 3785
rect 35350 3689 35402 3695
rect 35350 3631 35402 3637
rect 34988 2692 35284 2712
rect 35044 2690 35068 2692
rect 35124 2690 35148 2692
rect 35204 2690 35228 2692
rect 35066 2638 35068 2690
rect 35130 2638 35142 2690
rect 35204 2638 35206 2690
rect 35044 2636 35068 2638
rect 35124 2636 35148 2638
rect 35204 2636 35228 2638
rect 34988 2616 35284 2636
rect 35362 1568 35390 3631
rect 35446 3023 35498 3029
rect 35446 2965 35498 2971
rect 34786 1392 34910 1420
rect 35074 1540 35390 1568
rect 34678 1173 34730 1179
rect 34678 1115 34730 1121
rect 34786 800 34814 1392
rect 35074 1124 35102 1540
rect 35158 1469 35210 1475
rect 35458 1420 35486 2965
rect 35554 1475 35582 6887
rect 35638 3837 35690 3843
rect 35638 3779 35690 3785
rect 35158 1411 35210 1417
rect 34870 1099 34922 1105
rect 34870 1041 34922 1047
rect 34978 1096 35102 1124
rect 34882 800 34910 1041
rect 34978 800 35006 1096
rect 35170 800 35198 1411
rect 35266 1392 35486 1420
rect 35542 1469 35594 1475
rect 35542 1411 35594 1417
rect 35266 1124 35294 1392
rect 35446 1173 35498 1179
rect 35266 1096 35390 1124
rect 35446 1115 35498 1121
rect 35254 1025 35306 1031
rect 35254 967 35306 973
rect 35266 800 35294 967
rect 35362 800 35390 1096
rect 35458 800 35486 1115
rect 35650 800 35678 3779
rect 35734 3689 35786 3695
rect 35734 3631 35786 3637
rect 35746 800 35774 3631
rect 35842 800 35870 7405
rect 36406 6945 36458 6951
rect 36406 6887 36458 6893
rect 36310 6353 36362 6359
rect 36310 6295 36362 6301
rect 35926 6205 35978 6211
rect 35926 6147 35978 6153
rect 35938 5767 35966 6147
rect 35926 5761 35978 5767
rect 35926 5703 35978 5709
rect 36022 5687 36074 5693
rect 36022 5629 36074 5635
rect 36214 5687 36266 5693
rect 36214 5629 36266 5635
rect 36034 2894 36062 5629
rect 35938 2866 36062 2894
rect 36118 2949 36170 2955
rect 36118 2891 36170 2897
rect 35938 1031 35966 2866
rect 36130 1697 36158 2891
rect 36118 1691 36170 1697
rect 36118 1633 36170 1639
rect 36226 1420 36254 5629
rect 36322 1549 36350 6295
rect 36310 1543 36362 1549
rect 36310 1485 36362 1491
rect 36034 1392 36254 1420
rect 35926 1025 35978 1031
rect 35926 967 35978 973
rect 36034 800 36062 1392
rect 36118 1321 36170 1327
rect 36418 1272 36446 6887
rect 36502 5021 36554 5027
rect 36502 4963 36554 4969
rect 36514 3843 36542 4963
rect 36502 3837 36554 3843
rect 36502 3779 36554 3785
rect 36502 3689 36554 3695
rect 36502 3631 36554 3637
rect 36118 1263 36170 1269
rect 36130 800 36158 1263
rect 36226 1244 36446 1272
rect 36226 800 36254 1244
rect 36310 1173 36362 1179
rect 36310 1115 36362 1121
rect 36322 800 36350 1115
rect 36514 800 36542 3631
rect 36610 800 36638 7405
rect 36994 7099 37022 22205
rect 38050 8357 38270 8376
rect 38038 8351 38282 8357
rect 38090 8348 38230 8351
rect 38038 8293 38090 8299
rect 38230 8293 38282 8299
rect 38132 7946 38188 7955
rect 38132 7881 38188 7890
rect 38146 7659 38174 7881
rect 38132 7650 38188 7659
rect 38132 7585 38188 7594
rect 38038 7463 38090 7469
rect 38038 7405 38090 7411
rect 36982 7093 37034 7099
rect 36982 7035 37034 7041
rect 36694 7019 36746 7025
rect 36694 6961 36746 6967
rect 36706 3769 36734 6961
rect 36982 6945 37034 6951
rect 36982 6887 37034 6893
rect 37750 6945 37802 6951
rect 37750 6887 37802 6893
rect 36886 4947 36938 4953
rect 36886 4889 36938 4895
rect 36790 4355 36842 4361
rect 36790 4297 36842 4303
rect 36694 3763 36746 3769
rect 36694 3705 36746 3711
rect 36694 3615 36746 3621
rect 36694 3557 36746 3563
rect 36706 800 36734 3557
rect 36802 800 36830 4297
rect 36898 1105 36926 4889
rect 36886 1099 36938 1105
rect 36886 1041 36938 1047
rect 36994 800 37022 6887
rect 37270 6871 37322 6877
rect 37270 6813 37322 6819
rect 37366 6871 37418 6877
rect 37366 6813 37418 6819
rect 37282 6507 37310 6813
rect 37270 6501 37322 6507
rect 37270 6443 37322 6449
rect 37174 4281 37226 4287
rect 37174 4223 37226 4229
rect 37078 3911 37130 3917
rect 37078 3853 37130 3859
rect 37090 800 37118 3853
rect 37186 800 37214 4223
rect 37378 800 37406 6813
rect 37654 6797 37706 6803
rect 37654 6739 37706 6745
rect 37558 5687 37610 5693
rect 37558 5629 37610 5635
rect 37462 5613 37514 5619
rect 37462 5555 37514 5561
rect 37474 800 37502 5555
rect 37570 3621 37598 5629
rect 37558 3615 37610 3621
rect 37558 3557 37610 3563
rect 37558 3023 37610 3029
rect 37558 2965 37610 2971
rect 37570 800 37598 2965
rect 37666 800 37694 6739
rect 37762 5841 37790 6887
rect 37750 5835 37802 5841
rect 37750 5777 37802 5783
rect 37846 3837 37898 3843
rect 37846 3779 37898 3785
rect 37858 800 37886 3779
rect 37942 3689 37994 3695
rect 37942 3631 37994 3637
rect 37954 800 37982 3631
rect 38050 800 38078 7405
rect 38338 7025 38366 38041
rect 38914 15831 38942 55357
rect 39382 53417 39434 53423
rect 39382 53359 39434 53365
rect 38902 15825 38954 15831
rect 38902 15767 38954 15773
rect 38806 8277 38858 8283
rect 38806 8219 38858 8225
rect 38818 7765 38846 8219
rect 38806 7759 38858 7765
rect 38806 7701 38858 7707
rect 38806 7463 38858 7469
rect 38806 7405 38858 7411
rect 38326 7019 38378 7025
rect 38326 6961 38378 6967
rect 38614 7019 38666 7025
rect 38614 6961 38666 6967
rect 38518 6945 38570 6951
rect 38518 6887 38570 6893
rect 38530 6581 38558 6887
rect 38518 6575 38570 6581
rect 38518 6517 38570 6523
rect 38626 5120 38654 6961
rect 38434 5092 38654 5120
rect 38134 4281 38186 4287
rect 38134 4223 38186 4229
rect 38146 800 38174 4223
rect 38326 2949 38378 2955
rect 38326 2891 38378 2897
rect 38338 800 38366 2891
rect 38434 800 38462 5092
rect 38614 5021 38666 5027
rect 38614 4963 38666 4969
rect 38518 4133 38570 4139
rect 38518 4075 38570 4081
rect 38530 800 38558 4075
rect 38626 3917 38654 4963
rect 38614 3911 38666 3917
rect 38614 3853 38666 3859
rect 38710 3689 38762 3695
rect 38710 3631 38762 3637
rect 38722 800 38750 3631
rect 38818 800 38846 7405
rect 39394 7363 39422 53359
rect 39478 50235 39530 50241
rect 39478 50177 39530 50183
rect 39490 50093 39518 50177
rect 39478 50087 39530 50093
rect 39478 50029 39530 50035
rect 39380 7354 39436 7363
rect 39380 7289 39436 7298
rect 39382 7167 39434 7173
rect 39382 7109 39434 7115
rect 39286 6871 39338 6877
rect 39286 6813 39338 6819
rect 39298 6771 39326 6813
rect 39394 6803 39422 7109
rect 39382 6797 39434 6803
rect 39284 6762 39340 6771
rect 39382 6739 39434 6745
rect 39284 6697 39340 6706
rect 39490 6433 39518 50029
rect 39586 38549 39614 56319
rect 39574 38543 39626 38549
rect 39574 38485 39626 38491
rect 39778 17089 39806 56689
rect 40162 56531 40190 59200
rect 40150 56525 40202 56531
rect 40150 56467 40202 56473
rect 39862 56229 39914 56235
rect 39862 56171 39914 56177
rect 39874 17294 39902 56171
rect 40738 55717 40766 59200
rect 41218 56975 41246 59200
rect 41206 56969 41258 56975
rect 41206 56911 41258 56917
rect 41206 56821 41258 56827
rect 41206 56763 41258 56769
rect 40822 56747 40874 56753
rect 40822 56689 40874 56695
rect 40834 56161 40862 56689
rect 41110 56229 41162 56235
rect 41110 56171 41162 56177
rect 40822 56155 40874 56161
rect 40822 56097 40874 56103
rect 40726 55711 40778 55717
rect 40726 55653 40778 55659
rect 40822 55563 40874 55569
rect 40822 55505 40874 55511
rect 40054 52085 40106 52091
rect 40054 52027 40106 52033
rect 39874 17266 39998 17294
rect 39766 17083 39818 17089
rect 39766 17025 39818 17031
rect 39574 9683 39626 9689
rect 39574 9625 39626 9631
rect 39586 9171 39614 9625
rect 39574 9165 39626 9171
rect 39574 9107 39626 9113
rect 39574 8129 39626 8135
rect 39574 8071 39626 8077
rect 39586 7765 39614 8071
rect 39574 7759 39626 7765
rect 39574 7701 39626 7707
rect 39574 7463 39626 7469
rect 39574 7405 39626 7411
rect 39478 6427 39530 6433
rect 39478 6369 39530 6375
rect 38902 6353 38954 6359
rect 38902 6295 38954 6301
rect 38914 800 38942 6295
rect 39190 6131 39242 6137
rect 39190 6073 39242 6079
rect 39094 5687 39146 5693
rect 39094 5629 39146 5635
rect 38998 4355 39050 4361
rect 38998 4297 39050 4303
rect 39010 800 39038 4297
rect 39106 4287 39134 5629
rect 39094 4281 39146 4287
rect 39094 4223 39146 4229
rect 39202 800 39230 6073
rect 39286 5687 39338 5693
rect 39286 5629 39338 5635
rect 39298 800 39326 5629
rect 39382 5021 39434 5027
rect 39382 4963 39434 4969
rect 39394 3843 39422 4963
rect 39382 3837 39434 3843
rect 39382 3779 39434 3785
rect 39478 3689 39530 3695
rect 39478 3631 39530 3637
rect 39490 3344 39518 3631
rect 39394 3316 39518 3344
rect 39394 800 39422 3316
rect 39586 2894 39614 7405
rect 39862 7167 39914 7173
rect 39862 7109 39914 7115
rect 39766 4355 39818 4361
rect 39766 4297 39818 4303
rect 39670 3911 39722 3917
rect 39670 3853 39722 3859
rect 39490 2866 39614 2894
rect 39490 800 39518 2866
rect 39682 800 39710 3853
rect 39778 800 39806 4297
rect 39874 800 39902 7109
rect 39970 4805 39998 17266
rect 40066 9023 40094 52027
rect 40834 42767 40862 55505
rect 41014 44759 41066 44765
rect 41014 44701 41066 44707
rect 40822 42761 40874 42767
rect 40822 42703 40874 42709
rect 40342 29441 40394 29447
rect 40342 29383 40394 29389
rect 40054 9017 40106 9023
rect 40054 8959 40106 8965
rect 40354 8251 40382 29383
rect 41026 12974 41054 44701
rect 41122 31889 41150 56171
rect 41110 31883 41162 31889
rect 41110 31825 41162 31831
rect 40738 12946 41054 12974
rect 40630 9165 40682 9171
rect 40630 9107 40682 9113
rect 40340 8242 40396 8251
rect 40340 8177 40396 8186
rect 40054 7537 40106 7543
rect 40054 7479 40106 7485
rect 39958 4799 40010 4805
rect 39958 4741 40010 4747
rect 39958 3837 40010 3843
rect 39958 3779 40010 3785
rect 39970 2894 39998 3779
rect 40066 3251 40094 7479
rect 40642 6951 40670 9107
rect 40630 6945 40682 6951
rect 40630 6887 40682 6893
rect 40342 6353 40394 6359
rect 40342 6295 40394 6301
rect 40150 5021 40202 5027
rect 40150 4963 40202 4969
rect 40162 4139 40190 4963
rect 40150 4133 40202 4139
rect 40150 4075 40202 4081
rect 40246 3689 40298 3695
rect 40246 3631 40298 3637
rect 40258 3344 40286 3631
rect 40162 3316 40286 3344
rect 40054 3245 40106 3251
rect 40054 3187 40106 3193
rect 39970 2866 40094 2894
rect 40066 800 40094 2866
rect 40162 800 40190 3316
rect 40246 3245 40298 3251
rect 40246 3187 40298 3193
rect 40258 800 40286 3187
rect 40354 800 40382 6295
rect 40630 6279 40682 6285
rect 40630 6221 40682 6227
rect 40534 3023 40586 3029
rect 40534 2965 40586 2971
rect 40546 800 40574 2965
rect 40642 800 40670 6221
rect 40738 5883 40766 12946
rect 41110 8129 41162 8135
rect 41110 8071 41162 8077
rect 41122 7765 41150 8071
rect 41110 7759 41162 7765
rect 41110 7701 41162 7707
rect 41218 7044 41246 56763
rect 41794 56531 41822 59200
rect 42274 56531 42302 59200
rect 42850 56901 42878 59200
rect 42838 56895 42890 56901
rect 42838 56837 42890 56843
rect 42934 56747 42986 56753
rect 42934 56689 42986 56695
rect 41782 56525 41834 56531
rect 41782 56467 41834 56473
rect 42262 56525 42314 56531
rect 42262 56467 42314 56473
rect 42454 56377 42506 56383
rect 42454 56319 42506 56325
rect 41302 56303 41354 56309
rect 41302 56245 41354 56251
rect 41314 48539 41342 56245
rect 41302 48533 41354 48539
rect 41302 48475 41354 48481
rect 42466 45061 42494 56319
rect 42646 56229 42698 56235
rect 42646 56171 42698 56177
rect 42454 45055 42506 45061
rect 42454 44997 42506 45003
rect 42358 32919 42410 32925
rect 42358 32861 42410 32867
rect 41302 28997 41354 29003
rect 41302 28939 41354 28945
rect 40834 7016 41246 7044
rect 40724 5874 40780 5883
rect 40724 5809 40780 5818
rect 40726 5687 40778 5693
rect 40726 5629 40778 5635
rect 40738 800 40766 5629
rect 40834 3177 40862 7016
rect 41206 6575 41258 6581
rect 41206 6517 41258 6523
rect 40918 5021 40970 5027
rect 40918 4963 40970 4969
rect 41014 5021 41066 5027
rect 41014 4963 41066 4969
rect 40930 3917 40958 4963
rect 40918 3911 40970 3917
rect 40918 3853 40970 3859
rect 41026 3843 41054 4963
rect 41110 3911 41162 3917
rect 41110 3853 41162 3859
rect 41014 3837 41066 3843
rect 41014 3779 41066 3785
rect 41014 3689 41066 3695
rect 41014 3631 41066 3637
rect 40822 3171 40874 3177
rect 40822 3113 40874 3119
rect 41026 1420 41054 3631
rect 40930 1392 41054 1420
rect 40930 800 40958 1392
rect 41014 1321 41066 1327
rect 41014 1263 41066 1269
rect 41026 800 41054 1263
rect 41122 800 41150 3853
rect 41218 3251 41246 6517
rect 41314 6433 41342 28939
rect 41782 28109 41834 28115
rect 41782 28051 41834 28057
rect 41794 27893 41822 28051
rect 41782 27887 41834 27893
rect 41782 27829 41834 27835
rect 42370 17294 42398 32861
rect 42178 17266 42398 17294
rect 42178 12974 42206 17266
rect 42658 17237 42686 56171
rect 42742 23595 42794 23601
rect 42742 23537 42794 23543
rect 42646 17231 42698 17237
rect 42646 17173 42698 17179
rect 42754 12974 42782 23537
rect 42838 22781 42890 22787
rect 42838 22723 42890 22729
rect 42850 17294 42878 22723
rect 42946 17829 42974 56689
rect 43330 56531 43358 59200
rect 43798 57043 43850 57049
rect 43798 56985 43850 56991
rect 43318 56525 43370 56531
rect 43318 56467 43370 56473
rect 43126 53417 43178 53423
rect 43126 53359 43178 53365
rect 42934 17823 42986 17829
rect 42934 17765 42986 17771
rect 42850 17266 42974 17294
rect 41890 12946 42206 12974
rect 42274 12946 42782 12974
rect 41494 10275 41546 10281
rect 41494 10217 41546 10223
rect 41398 7463 41450 7469
rect 41398 7405 41450 7411
rect 41302 6427 41354 6433
rect 41302 6369 41354 6375
rect 41302 6279 41354 6285
rect 41302 6221 41354 6227
rect 41314 6137 41342 6221
rect 41302 6131 41354 6137
rect 41302 6073 41354 6079
rect 41302 3763 41354 3769
rect 41302 3705 41354 3711
rect 41206 3245 41258 3251
rect 41206 3187 41258 3193
rect 41206 2949 41258 2955
rect 41206 2891 41258 2897
rect 41218 800 41246 2891
rect 41314 1327 41342 3705
rect 41302 1321 41354 1327
rect 41302 1263 41354 1269
rect 41410 800 41438 7405
rect 41506 6285 41534 10217
rect 41590 9831 41642 9837
rect 41590 9773 41642 9779
rect 41602 7025 41630 9773
rect 41782 9757 41834 9763
rect 41782 9699 41834 9705
rect 41686 7167 41738 7173
rect 41686 7109 41738 7115
rect 41590 7019 41642 7025
rect 41590 6961 41642 6967
rect 41590 6871 41642 6877
rect 41590 6813 41642 6819
rect 41494 6279 41546 6285
rect 41494 6221 41546 6227
rect 41494 4281 41546 4287
rect 41494 4223 41546 4229
rect 41506 800 41534 4223
rect 41602 3769 41630 6813
rect 41590 3763 41642 3769
rect 41590 3705 41642 3711
rect 41590 3615 41642 3621
rect 41590 3557 41642 3563
rect 41602 800 41630 3557
rect 41698 800 41726 7109
rect 41794 7099 41822 9699
rect 41782 7093 41834 7099
rect 41782 7035 41834 7041
rect 41890 6475 41918 12946
rect 42274 7784 42302 12946
rect 42946 8949 42974 17266
rect 43138 12974 43166 53359
rect 43042 12946 43166 12974
rect 42934 8943 42986 8949
rect 42934 8885 42986 8891
rect 42646 8573 42698 8579
rect 42646 8515 42698 8521
rect 41986 7756 42302 7784
rect 42658 7765 42686 8515
rect 42646 7759 42698 7765
rect 41876 6466 41932 6475
rect 41876 6401 41932 6410
rect 41878 6353 41930 6359
rect 41878 6295 41930 6301
rect 41782 5687 41834 5693
rect 41782 5629 41834 5635
rect 41794 4287 41822 5629
rect 41782 4281 41834 4287
rect 41782 4223 41834 4229
rect 41890 800 41918 6295
rect 41986 5767 42014 7756
rect 42646 7701 42698 7707
rect 43042 7636 43070 12946
rect 42082 7608 43070 7636
rect 42082 6951 42110 7608
rect 42454 7463 42506 7469
rect 42454 7405 42506 7411
rect 42262 7093 42314 7099
rect 42262 7035 42314 7041
rect 42070 6945 42122 6951
rect 42070 6887 42122 6893
rect 42274 6507 42302 7035
rect 42358 6797 42410 6803
rect 42356 6762 42358 6771
rect 42410 6762 42412 6771
rect 42356 6697 42412 6706
rect 42262 6501 42314 6507
rect 42262 6443 42314 6449
rect 42358 6279 42410 6285
rect 42358 6221 42410 6227
rect 42370 6179 42398 6221
rect 42356 6170 42412 6179
rect 42356 6105 42412 6114
rect 41974 5761 42026 5767
rect 41974 5703 42026 5709
rect 42262 5687 42314 5693
rect 42262 5629 42314 5635
rect 42070 5021 42122 5027
rect 42070 4963 42122 4969
rect 41974 4355 42026 4361
rect 41974 4297 42026 4303
rect 41986 800 42014 4297
rect 42082 3917 42110 4963
rect 42070 3911 42122 3917
rect 42070 3853 42122 3859
rect 42070 3171 42122 3177
rect 42070 3113 42122 3119
rect 42082 800 42110 3113
rect 42274 800 42302 5629
rect 42358 4355 42410 4361
rect 42358 4297 42410 4303
rect 42370 800 42398 4297
rect 42466 800 42494 7405
rect 43222 7019 43274 7025
rect 43222 6961 43274 6967
rect 43126 6871 43178 6877
rect 43126 6813 43178 6819
rect 42646 6797 42698 6803
rect 42646 6739 42698 6745
rect 42658 6433 42686 6739
rect 42646 6427 42698 6433
rect 42646 6369 42698 6375
rect 42742 5909 42794 5915
rect 42742 5851 42794 5857
rect 42754 5619 42782 5851
rect 42742 5613 42794 5619
rect 42742 5555 42794 5561
rect 42742 3689 42794 3695
rect 42742 3631 42794 3637
rect 42550 3097 42602 3103
rect 42550 3039 42602 3045
rect 42562 800 42590 3039
rect 42754 800 42782 3631
rect 43138 3492 43166 6813
rect 43234 6581 43262 6961
rect 43222 6575 43274 6581
rect 43222 6517 43274 6523
rect 43700 6318 43756 6327
rect 43700 6253 43702 6262
rect 43754 6253 43756 6262
rect 43702 6221 43754 6227
rect 43318 5909 43370 5915
rect 43318 5851 43370 5857
rect 43222 5687 43274 5693
rect 43222 5629 43274 5635
rect 42850 3464 43166 3492
rect 42850 800 42878 3464
rect 43234 3196 43262 5629
rect 43330 5619 43358 5851
rect 43702 5687 43754 5693
rect 43702 5629 43754 5635
rect 43318 5613 43370 5619
rect 43318 5555 43370 5561
rect 43510 5021 43562 5027
rect 43510 4963 43562 4969
rect 43414 4355 43466 4361
rect 43414 4297 43466 4303
rect 43318 3911 43370 3917
rect 43318 3853 43370 3859
rect 42946 3168 43262 3196
rect 42946 800 42974 3168
rect 43030 3023 43082 3029
rect 43030 2965 43082 2971
rect 43042 800 43070 2965
rect 43222 2579 43274 2585
rect 43222 2521 43274 2527
rect 43234 800 43262 2521
rect 43330 800 43358 3853
rect 43426 800 43454 4297
rect 43522 3103 43550 4963
rect 43606 4281 43658 4287
rect 43606 4223 43658 4229
rect 43510 3097 43562 3103
rect 43510 3039 43562 3045
rect 43618 800 43646 4223
rect 43714 800 43742 5629
rect 43810 4583 43838 56985
rect 43906 56531 43934 59200
rect 43990 57413 44042 57419
rect 43990 57355 44042 57361
rect 43894 56525 43946 56531
rect 43894 56467 43946 56473
rect 43894 56377 43946 56383
rect 43894 56319 43946 56325
rect 43906 21603 43934 56319
rect 44002 41805 44030 57355
rect 44086 57043 44138 57049
rect 44086 56985 44138 56991
rect 44098 51499 44126 56985
rect 44386 56901 44414 59200
rect 44374 56895 44426 56901
rect 44374 56837 44426 56843
rect 44758 56747 44810 56753
rect 44758 56689 44810 56695
rect 44374 56229 44426 56235
rect 44374 56171 44426 56177
rect 44086 51493 44138 51499
rect 44086 51435 44138 51441
rect 44386 48761 44414 56171
rect 44470 53491 44522 53497
rect 44470 53433 44522 53439
rect 44374 48755 44426 48761
rect 44374 48697 44426 48703
rect 44374 44093 44426 44099
rect 44374 44035 44426 44041
rect 43990 41799 44042 41805
rect 43990 41741 44042 41747
rect 44086 39579 44138 39585
rect 44086 39521 44138 39527
rect 44098 39215 44126 39521
rect 44086 39209 44138 39215
rect 44086 39151 44138 39157
rect 43894 21597 43946 21603
rect 43894 21539 43946 21545
rect 44180 8094 44236 8103
rect 44180 8029 44236 8038
rect 44194 7839 44222 8029
rect 44386 7913 44414 44035
rect 44374 7907 44426 7913
rect 44374 7849 44426 7855
rect 44182 7833 44234 7839
rect 44182 7775 44234 7781
rect 43894 7463 43946 7469
rect 43894 7405 43946 7411
rect 43798 4577 43850 4583
rect 43798 4519 43850 4525
rect 43798 3615 43850 3621
rect 43798 3557 43850 3563
rect 43810 800 43838 3557
rect 43906 800 43934 7405
rect 44482 7099 44510 53433
rect 44566 40985 44618 40991
rect 44566 40927 44618 40933
rect 44470 7093 44522 7099
rect 44470 7035 44522 7041
rect 44278 6945 44330 6951
rect 44278 6887 44330 6893
rect 44374 6945 44426 6951
rect 44374 6887 44426 6893
rect 44182 6427 44234 6433
rect 44182 6369 44234 6375
rect 43990 6131 44042 6137
rect 43990 6073 44042 6079
rect 44002 2585 44030 6073
rect 44086 3837 44138 3843
rect 44086 3779 44138 3785
rect 43990 2579 44042 2585
rect 43990 2521 44042 2527
rect 44098 800 44126 3779
rect 44194 3177 44222 6369
rect 44182 3171 44234 3177
rect 44182 3113 44234 3119
rect 44182 2949 44234 2955
rect 44182 2891 44234 2897
rect 44194 800 44222 2891
rect 44290 800 44318 6887
rect 44386 4287 44414 6887
rect 44578 6581 44606 40927
rect 44770 18199 44798 56689
rect 44962 56531 44990 59200
rect 44950 56525 45002 56531
rect 44950 56467 45002 56473
rect 45442 55717 45470 59200
rect 45922 56901 45950 59200
rect 45910 56895 45962 56901
rect 45910 56837 45962 56843
rect 46102 56747 46154 56753
rect 46102 56689 46154 56695
rect 45430 55711 45482 55717
rect 45430 55653 45482 55659
rect 45142 55415 45194 55421
rect 45142 55357 45194 55363
rect 45154 30853 45182 55357
rect 45238 50753 45290 50759
rect 45238 50695 45290 50701
rect 45142 30847 45194 30853
rect 45142 30789 45194 30795
rect 44854 28923 44906 28929
rect 44854 28865 44906 28871
rect 44758 18193 44810 18199
rect 44758 18135 44810 18141
rect 44866 17294 44894 28865
rect 44866 17266 44990 17294
rect 44662 8943 44714 8949
rect 44662 8885 44714 8891
rect 44674 7839 44702 8885
rect 44662 7833 44714 7839
rect 44662 7775 44714 7781
rect 44662 7463 44714 7469
rect 44662 7405 44714 7411
rect 44566 6575 44618 6581
rect 44566 6517 44618 6523
rect 44578 6433 44606 6517
rect 44566 6427 44618 6433
rect 44566 6369 44618 6375
rect 44374 4281 44426 4287
rect 44374 4223 44426 4229
rect 44470 4281 44522 4287
rect 44470 4223 44522 4229
rect 44482 800 44510 4223
rect 44566 3541 44618 3547
rect 44566 3483 44618 3489
rect 44578 800 44606 3483
rect 44674 800 44702 7405
rect 44962 6507 44990 17266
rect 45142 13457 45194 13463
rect 45142 13399 45194 13405
rect 45154 13241 45182 13399
rect 45142 13235 45194 13241
rect 45142 13177 45194 13183
rect 45250 7913 45278 50695
rect 46114 18273 46142 56689
rect 46498 56531 46526 59200
rect 46486 56525 46538 56531
rect 46486 56467 46538 56473
rect 46870 56229 46922 56235
rect 46870 56171 46922 56177
rect 46390 42761 46442 42767
rect 46390 42703 46442 42709
rect 46198 36101 46250 36107
rect 46198 36043 46250 36049
rect 46294 36101 46346 36107
rect 46294 36043 46346 36049
rect 46102 18267 46154 18273
rect 46102 18209 46154 18215
rect 46102 8425 46154 8431
rect 46102 8367 46154 8373
rect 46114 8251 46142 8367
rect 46100 8242 46156 8251
rect 46100 8177 46156 8186
rect 46006 8129 46058 8135
rect 46006 8071 46058 8077
rect 45238 7907 45290 7913
rect 45238 7849 45290 7855
rect 46018 7839 46046 8071
rect 46006 7833 46058 7839
rect 46006 7775 46058 7781
rect 46006 7611 46058 7617
rect 46006 7553 46058 7559
rect 46018 7488 46046 7553
rect 46210 7488 46238 36043
rect 45046 7463 45098 7469
rect 45046 7405 45098 7411
rect 45814 7463 45866 7469
rect 46018 7460 46238 7488
rect 45814 7405 45866 7411
rect 44950 6501 45002 6507
rect 44950 6443 45002 6449
rect 44758 5021 44810 5027
rect 44758 4963 44810 4969
rect 44770 3917 44798 4963
rect 44950 4355 45002 4361
rect 44950 4297 45002 4303
rect 44758 3911 44810 3917
rect 44758 3853 44810 3859
rect 44854 3911 44906 3917
rect 44854 3853 44906 3859
rect 44866 2604 44894 3853
rect 44770 2576 44894 2604
rect 44770 800 44798 2576
rect 44962 800 44990 4297
rect 45058 800 45086 7405
rect 45334 6945 45386 6951
rect 45334 6887 45386 6893
rect 45142 5687 45194 5693
rect 45142 5629 45194 5635
rect 45154 4287 45182 5629
rect 45142 4281 45194 4287
rect 45142 4223 45194 4229
rect 45238 3763 45290 3769
rect 45238 3705 45290 3711
rect 45142 2579 45194 2585
rect 45142 2521 45194 2527
rect 45154 800 45182 2521
rect 45250 800 45278 3705
rect 45346 2807 45374 6887
rect 45622 6871 45674 6877
rect 45622 6813 45674 6819
rect 45526 6353 45578 6359
rect 45526 6295 45578 6301
rect 45430 5021 45482 5027
rect 45430 4963 45482 4969
rect 45442 3843 45470 4963
rect 45430 3837 45482 3843
rect 45430 3779 45482 3785
rect 45430 3467 45482 3473
rect 45430 3409 45482 3415
rect 45334 2801 45386 2807
rect 45334 2743 45386 2749
rect 45442 800 45470 3409
rect 45538 800 45566 6295
rect 45634 3473 45662 6813
rect 45718 3541 45770 3547
rect 45718 3483 45770 3489
rect 45622 3467 45674 3473
rect 45622 3409 45674 3415
rect 45622 3023 45674 3029
rect 45622 2965 45674 2971
rect 45634 800 45662 2965
rect 45730 2585 45758 3483
rect 45718 2579 45770 2585
rect 45718 2521 45770 2527
rect 45826 800 45854 7405
rect 46306 7067 46334 36043
rect 46402 12974 46430 42703
rect 46882 39881 46910 56171
rect 46978 55717 47006 59200
rect 47554 56975 47582 59200
rect 47542 56969 47594 56975
rect 47542 56911 47594 56917
rect 48034 56531 48062 59200
rect 48022 56525 48074 56531
rect 48022 56467 48074 56473
rect 48610 56161 48638 59200
rect 49090 56901 49118 59200
rect 49078 56895 49130 56901
rect 49078 56837 49130 56843
rect 48694 56747 48746 56753
rect 48694 56689 48746 56695
rect 48706 56457 48734 56689
rect 49666 56531 49694 59200
rect 50146 56531 50174 59200
rect 50722 56901 50750 59200
rect 51202 57614 51230 59200
rect 51202 57586 51326 57614
rect 50710 56895 50762 56901
rect 50710 56837 50762 56843
rect 50806 56747 50858 56753
rect 50806 56689 50858 56695
rect 50348 56638 50644 56658
rect 50404 56636 50428 56638
rect 50484 56636 50508 56638
rect 50564 56636 50588 56638
rect 50426 56584 50428 56636
rect 50490 56584 50502 56636
rect 50564 56584 50566 56636
rect 50404 56582 50428 56584
rect 50484 56582 50508 56584
rect 50564 56582 50588 56584
rect 50348 56562 50644 56582
rect 49654 56525 49706 56531
rect 49654 56467 49706 56473
rect 50134 56525 50186 56531
rect 50134 56467 50186 56473
rect 48694 56451 48746 56457
rect 48694 56393 48746 56399
rect 48886 56229 48938 56235
rect 48886 56171 48938 56177
rect 48598 56155 48650 56161
rect 48598 56097 48650 56103
rect 46966 55711 47018 55717
rect 46966 55653 47018 55659
rect 47158 55563 47210 55569
rect 47158 55505 47210 55511
rect 47170 55125 47198 55505
rect 47158 55119 47210 55125
rect 47158 55061 47210 55067
rect 46870 39875 46922 39881
rect 46870 39817 46922 39823
rect 47734 33437 47786 33443
rect 47734 33379 47786 33385
rect 47746 33221 47774 33379
rect 47734 33215 47786 33221
rect 47734 33157 47786 33163
rect 48310 31735 48362 31741
rect 48310 31677 48362 31683
rect 46402 12946 46526 12974
rect 46390 8795 46442 8801
rect 46390 8737 46442 8743
rect 46402 8357 46430 8737
rect 46498 8579 46526 12946
rect 48214 10793 48266 10799
rect 48214 10735 48266 10741
rect 48226 10577 48254 10735
rect 48214 10571 48266 10577
rect 48214 10513 48266 10519
rect 47542 9461 47594 9467
rect 47542 9403 47594 9409
rect 46486 8573 46538 8579
rect 46486 8515 46538 8521
rect 46390 8351 46442 8357
rect 46390 8293 46442 8299
rect 47554 8283 47582 9403
rect 47926 8573 47978 8579
rect 47926 8515 47978 8521
rect 47542 8277 47594 8283
rect 46484 8242 46540 8251
rect 47542 8219 47594 8225
rect 46484 8177 46540 8186
rect 46498 7839 46526 8177
rect 47938 8103 47966 8515
rect 48022 8277 48074 8283
rect 48022 8219 48074 8225
rect 47924 8094 47980 8103
rect 47924 8029 47980 8038
rect 46486 7833 46538 7839
rect 46486 7775 46538 7781
rect 47254 7759 47306 7765
rect 47254 7701 47306 7707
rect 46486 7463 46538 7469
rect 46486 7405 46538 7411
rect 46292 7058 46348 7067
rect 46292 6993 46348 7002
rect 46390 6945 46442 6951
rect 46390 6887 46442 6893
rect 46402 6803 46430 6887
rect 46390 6797 46442 6803
rect 46390 6739 46442 6745
rect 46402 6031 46430 6739
rect 46388 6022 46444 6031
rect 46388 5957 46444 5966
rect 46102 5687 46154 5693
rect 46102 5629 46154 5635
rect 46114 4232 46142 5629
rect 46198 5021 46250 5027
rect 46198 4963 46250 4969
rect 46390 5021 46442 5027
rect 46390 4963 46442 4969
rect 45922 4204 46142 4232
rect 45922 800 45950 4204
rect 46210 3917 46238 4963
rect 46198 3911 46250 3917
rect 46198 3853 46250 3859
rect 46294 3911 46346 3917
rect 46294 3853 46346 3859
rect 46006 3615 46058 3621
rect 46006 3557 46058 3563
rect 46018 800 46046 3557
rect 46102 2801 46154 2807
rect 46102 2743 46154 2749
rect 46114 800 46142 2743
rect 46306 800 46334 3853
rect 46402 3547 46430 4963
rect 46390 3541 46442 3547
rect 46390 3483 46442 3489
rect 46390 3097 46442 3103
rect 46390 3039 46442 3045
rect 46402 800 46430 3039
rect 46498 800 46526 7405
rect 46870 7019 46922 7025
rect 46870 6961 46922 6967
rect 46582 6575 46634 6581
rect 46582 6517 46634 6523
rect 46594 6211 46622 6517
rect 46582 6205 46634 6211
rect 46582 6147 46634 6153
rect 46678 5687 46730 5693
rect 46678 5629 46730 5635
rect 46690 2894 46718 5629
rect 46774 4355 46826 4361
rect 46774 4297 46826 4303
rect 46594 2866 46718 2894
rect 46594 800 46622 2866
rect 46786 800 46814 4297
rect 46882 800 46910 6961
rect 47158 6945 47210 6951
rect 47158 6887 47210 6893
rect 47062 6871 47114 6877
rect 47062 6813 47114 6819
rect 46966 6353 47018 6359
rect 46966 6295 47018 6301
rect 46978 800 47006 6295
rect 47074 2807 47102 6813
rect 47170 6803 47198 6887
rect 47158 6797 47210 6803
rect 47158 6739 47210 6745
rect 47170 5915 47198 6739
rect 47158 5909 47210 5915
rect 47158 5851 47210 5857
rect 47158 3689 47210 3695
rect 47158 3631 47210 3637
rect 47062 2801 47114 2807
rect 47062 2743 47114 2749
rect 47170 800 47198 3631
rect 47266 800 47294 7701
rect 47638 7611 47690 7617
rect 47638 7553 47690 7559
rect 47650 7469 47678 7553
rect 47638 7463 47690 7469
rect 47638 7405 47690 7411
rect 47542 5687 47594 5693
rect 47542 5629 47594 5635
rect 47554 4380 47582 5629
rect 47650 5471 47678 7405
rect 47734 6353 47786 6359
rect 47734 6295 47786 6301
rect 47638 5465 47690 5471
rect 47638 5407 47690 5413
rect 47638 5021 47690 5027
rect 47638 4963 47690 4969
rect 47362 4352 47582 4380
rect 47362 800 47390 4352
rect 47446 4281 47498 4287
rect 47446 4223 47498 4229
rect 47458 800 47486 4223
rect 47650 3917 47678 4963
rect 47638 3911 47690 3917
rect 47638 3853 47690 3859
rect 47542 3763 47594 3769
rect 47542 3705 47594 3711
rect 47554 2752 47582 3705
rect 47554 2724 47678 2752
rect 47650 800 47678 2724
rect 47746 800 47774 6295
rect 47830 4355 47882 4361
rect 47830 4297 47882 4303
rect 47842 800 47870 4297
rect 48034 800 48062 8219
rect 48322 7099 48350 31677
rect 48898 18347 48926 56171
rect 49174 55415 49226 55421
rect 49174 55357 49226 55363
rect 48886 18341 48938 18347
rect 48886 18283 48938 18289
rect 48886 17453 48938 17459
rect 48886 17395 48938 17401
rect 48898 8431 48926 17395
rect 49186 12974 49214 55357
rect 50348 55306 50644 55326
rect 50404 55304 50428 55306
rect 50484 55304 50508 55306
rect 50564 55304 50588 55306
rect 50426 55252 50428 55304
rect 50490 55252 50502 55304
rect 50564 55252 50566 55304
rect 50404 55250 50428 55252
rect 50484 55250 50508 55252
rect 50564 55250 50588 55252
rect 50348 55230 50644 55250
rect 50230 54823 50282 54829
rect 50230 54765 50282 54771
rect 50038 43427 50090 43433
rect 50038 43369 50090 43375
rect 49942 29441 49994 29447
rect 49942 29383 49994 29389
rect 49846 24927 49898 24933
rect 49846 24869 49898 24875
rect 49090 12946 49214 12974
rect 49090 9837 49118 12946
rect 49078 9831 49130 9837
rect 49078 9773 49130 9779
rect 49858 9171 49886 24869
rect 49954 9763 49982 29383
rect 49942 9757 49994 9763
rect 49942 9699 49994 9705
rect 49846 9165 49898 9171
rect 49846 9107 49898 9113
rect 48886 8425 48938 8431
rect 48886 8367 48938 8373
rect 48694 8277 48746 8283
rect 48694 8219 48746 8225
rect 49462 8277 49514 8283
rect 49462 8219 49514 8225
rect 48406 7759 48458 7765
rect 48406 7701 48458 7707
rect 48310 7093 48362 7099
rect 48310 7035 48362 7041
rect 48310 6945 48362 6951
rect 48310 6887 48362 6893
rect 48118 4133 48170 4139
rect 48118 4075 48170 4081
rect 48130 800 48158 4075
rect 48322 3769 48350 6887
rect 48310 3763 48362 3769
rect 48310 3705 48362 3711
rect 48214 3689 48266 3695
rect 48214 3631 48266 3637
rect 48226 800 48254 3631
rect 48418 2894 48446 7701
rect 48502 7019 48554 7025
rect 48502 6961 48554 6967
rect 48514 6771 48542 6961
rect 48500 6762 48556 6771
rect 48500 6697 48556 6706
rect 48598 4281 48650 4287
rect 48598 4223 48650 4229
rect 48502 3911 48554 3917
rect 48502 3853 48554 3859
rect 48322 2866 48446 2894
rect 48322 800 48350 2866
rect 48514 800 48542 3853
rect 48610 800 48638 4223
rect 48706 800 48734 8219
rect 48790 6353 48842 6359
rect 48790 6295 48842 6301
rect 48802 800 48830 6295
rect 48982 5687 49034 5693
rect 48982 5629 49034 5635
rect 48994 4139 49022 5629
rect 49366 5021 49418 5027
rect 49366 4963 49418 4969
rect 49174 4355 49226 4361
rect 49174 4297 49226 4303
rect 48982 4133 49034 4139
rect 48982 4075 49034 4081
rect 49186 3640 49214 4297
rect 49270 4133 49322 4139
rect 49270 4075 49322 4081
rect 48994 3612 49214 3640
rect 48994 800 49022 3612
rect 49078 3541 49130 3547
rect 49078 3483 49130 3489
rect 49090 800 49118 3483
rect 49282 2894 49310 4075
rect 49186 2866 49310 2894
rect 49186 800 49214 2866
rect 49378 800 49406 4963
rect 49474 800 49502 8219
rect 50050 7955 50078 43369
rect 50134 18267 50186 18273
rect 50134 18209 50186 18215
rect 50036 7946 50092 7955
rect 50036 7881 50092 7890
rect 50146 7765 50174 18209
rect 50134 7759 50186 7765
rect 50134 7701 50186 7707
rect 50038 7463 50090 7469
rect 50038 7405 50090 7411
rect 49558 6353 49610 6359
rect 49558 6295 49610 6301
rect 49570 800 49598 6295
rect 49846 6131 49898 6137
rect 49846 6073 49898 6079
rect 49654 5687 49706 5693
rect 49654 5629 49706 5635
rect 49666 3917 49694 5629
rect 49654 3911 49706 3917
rect 49654 3853 49706 3859
rect 49654 3023 49706 3029
rect 49654 2965 49706 2971
rect 49666 800 49694 2965
rect 49858 800 49886 6073
rect 49942 4281 49994 4287
rect 49942 4223 49994 4229
rect 49954 800 49982 4223
rect 50050 3547 50078 7405
rect 50242 7099 50270 54765
rect 50348 53974 50644 53994
rect 50404 53972 50428 53974
rect 50484 53972 50508 53974
rect 50564 53972 50588 53974
rect 50426 53920 50428 53972
rect 50490 53920 50502 53972
rect 50564 53920 50566 53972
rect 50404 53918 50428 53920
rect 50484 53918 50508 53920
rect 50564 53918 50588 53920
rect 50348 53898 50644 53918
rect 50348 52642 50644 52662
rect 50404 52640 50428 52642
rect 50484 52640 50508 52642
rect 50564 52640 50588 52642
rect 50426 52588 50428 52640
rect 50490 52588 50502 52640
rect 50564 52588 50566 52640
rect 50404 52586 50428 52588
rect 50484 52586 50508 52588
rect 50564 52586 50588 52588
rect 50348 52566 50644 52586
rect 50348 51310 50644 51330
rect 50404 51308 50428 51310
rect 50484 51308 50508 51310
rect 50564 51308 50588 51310
rect 50426 51256 50428 51308
rect 50490 51256 50502 51308
rect 50564 51256 50566 51308
rect 50404 51254 50428 51256
rect 50484 51254 50508 51256
rect 50564 51254 50588 51256
rect 50348 51234 50644 51254
rect 50348 49978 50644 49998
rect 50404 49976 50428 49978
rect 50484 49976 50508 49978
rect 50564 49976 50588 49978
rect 50426 49924 50428 49976
rect 50490 49924 50502 49976
rect 50564 49924 50566 49976
rect 50404 49922 50428 49924
rect 50484 49922 50508 49924
rect 50564 49922 50588 49924
rect 50348 49902 50644 49922
rect 50348 48646 50644 48666
rect 50404 48644 50428 48646
rect 50484 48644 50508 48646
rect 50564 48644 50588 48646
rect 50426 48592 50428 48644
rect 50490 48592 50502 48644
rect 50564 48592 50566 48644
rect 50404 48590 50428 48592
rect 50484 48590 50508 48592
rect 50564 48590 50588 48592
rect 50348 48570 50644 48590
rect 50348 47314 50644 47334
rect 50404 47312 50428 47314
rect 50484 47312 50508 47314
rect 50564 47312 50588 47314
rect 50426 47260 50428 47312
rect 50490 47260 50502 47312
rect 50564 47260 50566 47312
rect 50404 47258 50428 47260
rect 50484 47258 50508 47260
rect 50564 47258 50588 47260
rect 50348 47238 50644 47258
rect 50348 45982 50644 46002
rect 50404 45980 50428 45982
rect 50484 45980 50508 45982
rect 50564 45980 50588 45982
rect 50426 45928 50428 45980
rect 50490 45928 50502 45980
rect 50564 45928 50566 45980
rect 50404 45926 50428 45928
rect 50484 45926 50508 45928
rect 50564 45926 50588 45928
rect 50348 45906 50644 45926
rect 50348 44650 50644 44670
rect 50404 44648 50428 44650
rect 50484 44648 50508 44650
rect 50564 44648 50588 44650
rect 50426 44596 50428 44648
rect 50490 44596 50502 44648
rect 50564 44596 50566 44648
rect 50404 44594 50428 44596
rect 50484 44594 50508 44596
rect 50564 44594 50588 44596
rect 50348 44574 50644 44594
rect 50348 43318 50644 43338
rect 50404 43316 50428 43318
rect 50484 43316 50508 43318
rect 50564 43316 50588 43318
rect 50426 43264 50428 43316
rect 50490 43264 50502 43316
rect 50564 43264 50566 43316
rect 50404 43262 50428 43264
rect 50484 43262 50508 43264
rect 50564 43262 50588 43264
rect 50348 43242 50644 43262
rect 50348 41986 50644 42006
rect 50404 41984 50428 41986
rect 50484 41984 50508 41986
rect 50564 41984 50588 41986
rect 50426 41932 50428 41984
rect 50490 41932 50502 41984
rect 50564 41932 50566 41984
rect 50404 41930 50428 41932
rect 50484 41930 50508 41932
rect 50564 41930 50588 41932
rect 50348 41910 50644 41930
rect 50348 40654 50644 40674
rect 50404 40652 50428 40654
rect 50484 40652 50508 40654
rect 50564 40652 50588 40654
rect 50426 40600 50428 40652
rect 50490 40600 50502 40652
rect 50564 40600 50566 40652
rect 50404 40598 50428 40600
rect 50484 40598 50508 40600
rect 50564 40598 50588 40600
rect 50348 40578 50644 40598
rect 50348 39322 50644 39342
rect 50404 39320 50428 39322
rect 50484 39320 50508 39322
rect 50564 39320 50588 39322
rect 50426 39268 50428 39320
rect 50490 39268 50502 39320
rect 50564 39268 50566 39320
rect 50404 39266 50428 39268
rect 50484 39266 50508 39268
rect 50564 39266 50588 39268
rect 50348 39246 50644 39266
rect 50348 37990 50644 38010
rect 50404 37988 50428 37990
rect 50484 37988 50508 37990
rect 50564 37988 50588 37990
rect 50426 37936 50428 37988
rect 50490 37936 50502 37988
rect 50564 37936 50566 37988
rect 50404 37934 50428 37936
rect 50484 37934 50508 37936
rect 50564 37934 50588 37936
rect 50348 37914 50644 37934
rect 50348 36658 50644 36678
rect 50404 36656 50428 36658
rect 50484 36656 50508 36658
rect 50564 36656 50588 36658
rect 50426 36604 50428 36656
rect 50490 36604 50502 36656
rect 50564 36604 50566 36656
rect 50404 36602 50428 36604
rect 50484 36602 50508 36604
rect 50564 36602 50588 36604
rect 50348 36582 50644 36602
rect 50348 35326 50644 35346
rect 50404 35324 50428 35326
rect 50484 35324 50508 35326
rect 50564 35324 50588 35326
rect 50426 35272 50428 35324
rect 50490 35272 50502 35324
rect 50564 35272 50566 35324
rect 50404 35270 50428 35272
rect 50484 35270 50508 35272
rect 50564 35270 50588 35272
rect 50348 35250 50644 35270
rect 50348 33994 50644 34014
rect 50404 33992 50428 33994
rect 50484 33992 50508 33994
rect 50564 33992 50588 33994
rect 50426 33940 50428 33992
rect 50490 33940 50502 33992
rect 50564 33940 50566 33992
rect 50404 33938 50428 33940
rect 50484 33938 50508 33940
rect 50564 33938 50588 33940
rect 50348 33918 50644 33938
rect 50348 32662 50644 32682
rect 50404 32660 50428 32662
rect 50484 32660 50508 32662
rect 50564 32660 50588 32662
rect 50426 32608 50428 32660
rect 50490 32608 50502 32660
rect 50564 32608 50566 32660
rect 50404 32606 50428 32608
rect 50484 32606 50508 32608
rect 50564 32606 50588 32608
rect 50348 32586 50644 32606
rect 50348 31330 50644 31350
rect 50404 31328 50428 31330
rect 50484 31328 50508 31330
rect 50564 31328 50588 31330
rect 50426 31276 50428 31328
rect 50490 31276 50502 31328
rect 50564 31276 50566 31328
rect 50404 31274 50428 31276
rect 50484 31274 50508 31276
rect 50564 31274 50588 31276
rect 50348 31254 50644 31274
rect 50348 29998 50644 30018
rect 50404 29996 50428 29998
rect 50484 29996 50508 29998
rect 50564 29996 50588 29998
rect 50426 29944 50428 29996
rect 50490 29944 50502 29996
rect 50564 29944 50566 29996
rect 50404 29942 50428 29944
rect 50484 29942 50508 29944
rect 50564 29942 50588 29944
rect 50348 29922 50644 29942
rect 50614 29441 50666 29447
rect 50614 29383 50666 29389
rect 50626 29225 50654 29383
rect 50614 29219 50666 29225
rect 50614 29161 50666 29167
rect 50348 28666 50644 28686
rect 50404 28664 50428 28666
rect 50484 28664 50508 28666
rect 50564 28664 50588 28666
rect 50426 28612 50428 28664
rect 50490 28612 50502 28664
rect 50564 28612 50566 28664
rect 50404 28610 50428 28612
rect 50484 28610 50508 28612
rect 50564 28610 50588 28612
rect 50348 28590 50644 28610
rect 50348 27334 50644 27354
rect 50404 27332 50428 27334
rect 50484 27332 50508 27334
rect 50564 27332 50588 27334
rect 50426 27280 50428 27332
rect 50490 27280 50502 27332
rect 50564 27280 50566 27332
rect 50404 27278 50428 27280
rect 50484 27278 50508 27280
rect 50564 27278 50588 27280
rect 50348 27258 50644 27278
rect 50348 26002 50644 26022
rect 50404 26000 50428 26002
rect 50484 26000 50508 26002
rect 50564 26000 50588 26002
rect 50426 25948 50428 26000
rect 50490 25948 50502 26000
rect 50564 25948 50566 26000
rect 50404 25946 50428 25948
rect 50484 25946 50508 25948
rect 50564 25946 50588 25948
rect 50348 25926 50644 25946
rect 50348 24670 50644 24690
rect 50404 24668 50428 24670
rect 50484 24668 50508 24670
rect 50564 24668 50588 24670
rect 50426 24616 50428 24668
rect 50490 24616 50502 24668
rect 50564 24616 50566 24668
rect 50404 24614 50428 24616
rect 50484 24614 50508 24616
rect 50564 24614 50588 24616
rect 50348 24594 50644 24614
rect 50348 23338 50644 23358
rect 50404 23336 50428 23338
rect 50484 23336 50508 23338
rect 50564 23336 50588 23338
rect 50426 23284 50428 23336
rect 50490 23284 50502 23336
rect 50564 23284 50566 23336
rect 50404 23282 50428 23284
rect 50484 23282 50508 23284
rect 50564 23282 50588 23284
rect 50348 23262 50644 23282
rect 50348 22006 50644 22026
rect 50404 22004 50428 22006
rect 50484 22004 50508 22006
rect 50564 22004 50588 22006
rect 50426 21952 50428 22004
rect 50490 21952 50502 22004
rect 50564 21952 50566 22004
rect 50404 21950 50428 21952
rect 50484 21950 50508 21952
rect 50564 21950 50588 21952
rect 50348 21930 50644 21950
rect 50348 20674 50644 20694
rect 50404 20672 50428 20674
rect 50484 20672 50508 20674
rect 50564 20672 50588 20674
rect 50426 20620 50428 20672
rect 50490 20620 50502 20672
rect 50564 20620 50566 20672
rect 50404 20618 50428 20620
rect 50484 20618 50508 20620
rect 50564 20618 50588 20620
rect 50348 20598 50644 20618
rect 50348 19342 50644 19362
rect 50404 19340 50428 19342
rect 50484 19340 50508 19342
rect 50564 19340 50588 19342
rect 50426 19288 50428 19340
rect 50490 19288 50502 19340
rect 50564 19288 50566 19340
rect 50404 19286 50428 19288
rect 50484 19286 50508 19288
rect 50564 19286 50588 19288
rect 50348 19266 50644 19286
rect 50818 19235 50846 56689
rect 51298 56531 51326 57586
rect 51286 56525 51338 56531
rect 51286 56467 51338 56473
rect 51778 55717 51806 59200
rect 52054 57043 52106 57049
rect 52054 56985 52106 56991
rect 52066 56309 52094 56985
rect 52258 56975 52286 59200
rect 52246 56969 52298 56975
rect 52246 56911 52298 56917
rect 52834 56531 52862 59200
rect 53314 56531 53342 59200
rect 53890 56901 53918 59200
rect 53878 56895 53930 56901
rect 53878 56837 53930 56843
rect 53974 56747 54026 56753
rect 53974 56689 54026 56695
rect 52822 56525 52874 56531
rect 52822 56467 52874 56473
rect 53302 56525 53354 56531
rect 53302 56467 53354 56473
rect 52054 56303 52106 56309
rect 52054 56245 52106 56251
rect 52630 56229 52682 56235
rect 52630 56171 52682 56177
rect 53686 56229 53738 56235
rect 53686 56171 53738 56177
rect 51766 55711 51818 55717
rect 51766 55653 51818 55659
rect 51670 52899 51722 52905
rect 51670 52841 51722 52847
rect 51574 45425 51626 45431
rect 51574 45367 51626 45373
rect 51586 45135 51614 45367
rect 51574 45129 51626 45135
rect 51574 45071 51626 45077
rect 51286 37433 51338 37439
rect 51286 37375 51338 37381
rect 50806 19229 50858 19235
rect 50806 19171 50858 19177
rect 50348 18010 50644 18030
rect 50404 18008 50428 18010
rect 50484 18008 50508 18010
rect 50564 18008 50588 18010
rect 50426 17956 50428 18008
rect 50490 17956 50502 18008
rect 50564 17956 50566 18008
rect 50404 17954 50428 17956
rect 50484 17954 50508 17956
rect 50564 17954 50588 17956
rect 50348 17934 50644 17954
rect 50348 16678 50644 16698
rect 50404 16676 50428 16678
rect 50484 16676 50508 16678
rect 50564 16676 50588 16678
rect 50426 16624 50428 16676
rect 50490 16624 50502 16676
rect 50564 16624 50566 16676
rect 50404 16622 50428 16624
rect 50484 16622 50508 16624
rect 50564 16622 50588 16624
rect 50348 16602 50644 16622
rect 50348 15346 50644 15366
rect 50404 15344 50428 15346
rect 50484 15344 50508 15346
rect 50564 15344 50588 15346
rect 50426 15292 50428 15344
rect 50490 15292 50502 15344
rect 50564 15292 50566 15344
rect 50404 15290 50428 15292
rect 50484 15290 50508 15292
rect 50564 15290 50588 15292
rect 50348 15270 50644 15290
rect 51190 14271 51242 14277
rect 51190 14213 51242 14219
rect 50348 14014 50644 14034
rect 50404 14012 50428 14014
rect 50484 14012 50508 14014
rect 50564 14012 50588 14014
rect 50426 13960 50428 14012
rect 50490 13960 50502 14012
rect 50564 13960 50566 14012
rect 50404 13958 50428 13960
rect 50484 13958 50508 13960
rect 50564 13958 50588 13960
rect 50348 13938 50644 13958
rect 50348 12682 50644 12702
rect 50404 12680 50428 12682
rect 50484 12680 50508 12682
rect 50564 12680 50588 12682
rect 50426 12628 50428 12680
rect 50490 12628 50502 12680
rect 50564 12628 50566 12680
rect 50404 12626 50428 12628
rect 50484 12626 50508 12628
rect 50564 12626 50588 12628
rect 50348 12606 50644 12626
rect 50348 11350 50644 11370
rect 50404 11348 50428 11350
rect 50484 11348 50508 11350
rect 50564 11348 50588 11350
rect 50426 11296 50428 11348
rect 50490 11296 50502 11348
rect 50564 11296 50566 11348
rect 50404 11294 50428 11296
rect 50484 11294 50508 11296
rect 50564 11294 50588 11296
rect 50348 11274 50644 11294
rect 50348 10018 50644 10038
rect 50404 10016 50428 10018
rect 50484 10016 50508 10018
rect 50564 10016 50588 10018
rect 50426 9964 50428 10016
rect 50490 9964 50502 10016
rect 50564 9964 50566 10016
rect 50404 9962 50428 9964
rect 50484 9962 50508 9964
rect 50564 9962 50588 9964
rect 50348 9942 50644 9962
rect 50348 8686 50644 8706
rect 50404 8684 50428 8686
rect 50484 8684 50508 8686
rect 50564 8684 50588 8686
rect 50426 8632 50428 8684
rect 50490 8632 50502 8684
rect 50564 8632 50566 8684
rect 50404 8630 50428 8632
rect 50484 8630 50508 8632
rect 50564 8630 50588 8632
rect 50348 8610 50644 8630
rect 51202 7913 51230 14213
rect 51190 7907 51242 7913
rect 51190 7849 51242 7855
rect 50348 7354 50644 7374
rect 50404 7352 50428 7354
rect 50484 7352 50508 7354
rect 50564 7352 50588 7354
rect 50426 7300 50428 7352
rect 50490 7300 50502 7352
rect 50564 7300 50566 7352
rect 50404 7298 50428 7300
rect 50484 7298 50508 7300
rect 50564 7298 50588 7300
rect 50348 7278 50644 7298
rect 50230 7093 50282 7099
rect 50230 7035 50282 7041
rect 50134 6871 50186 6877
rect 50134 6813 50186 6819
rect 50422 6871 50474 6877
rect 50422 6813 50474 6819
rect 50038 3541 50090 3547
rect 50038 3483 50090 3489
rect 50038 2875 50090 2881
rect 50038 2817 50090 2823
rect 50050 800 50078 2817
rect 50146 800 50174 6813
rect 50434 6433 50462 6813
rect 51298 6581 51326 37375
rect 51682 7173 51710 52841
rect 52438 49421 52490 49427
rect 52438 49363 52490 49369
rect 51766 48903 51818 48909
rect 51766 48845 51818 48851
rect 51778 7765 51806 48845
rect 52246 48089 52298 48095
rect 52246 48031 52298 48037
rect 52258 17294 52286 48031
rect 52342 41429 52394 41435
rect 52342 41371 52394 41377
rect 52162 17266 52286 17294
rect 51862 7907 51914 7913
rect 51862 7849 51914 7855
rect 51766 7759 51818 7765
rect 51766 7701 51818 7707
rect 51874 7617 51902 7849
rect 51862 7611 51914 7617
rect 51862 7553 51914 7559
rect 52162 7511 52190 17266
rect 52354 12974 52382 41371
rect 52258 12946 52382 12974
rect 52148 7502 52204 7511
rect 51766 7463 51818 7469
rect 52148 7437 52204 7446
rect 51766 7405 51818 7411
rect 51670 7167 51722 7173
rect 51670 7109 51722 7115
rect 51478 6945 51530 6951
rect 51478 6887 51530 6893
rect 51286 6575 51338 6581
rect 51286 6517 51338 6523
rect 50422 6427 50474 6433
rect 50422 6369 50474 6375
rect 51094 6131 51146 6137
rect 51094 6073 51146 6079
rect 50348 6022 50644 6042
rect 50404 6020 50428 6022
rect 50484 6020 50508 6022
rect 50564 6020 50588 6022
rect 50426 5968 50428 6020
rect 50490 5968 50502 6020
rect 50564 5968 50566 6020
rect 50404 5966 50428 5968
rect 50484 5966 50508 5968
rect 50564 5966 50588 5968
rect 50348 5946 50644 5966
rect 50710 5687 50762 5693
rect 50710 5629 50762 5635
rect 50422 5021 50474 5027
rect 50422 4963 50474 4969
rect 50434 4824 50462 4963
rect 50242 4796 50462 4824
rect 50242 2604 50270 4796
rect 50348 4690 50644 4710
rect 50404 4688 50428 4690
rect 50484 4688 50508 4690
rect 50564 4688 50588 4690
rect 50426 4636 50428 4688
rect 50490 4636 50502 4688
rect 50564 4636 50566 4688
rect 50404 4634 50428 4636
rect 50484 4634 50508 4636
rect 50564 4634 50588 4636
rect 50348 4614 50644 4634
rect 50722 4139 50750 5629
rect 50902 5021 50954 5027
rect 50902 4963 50954 4969
rect 50710 4133 50762 4139
rect 50710 4075 50762 4081
rect 50710 3689 50762 3695
rect 50710 3631 50762 3637
rect 50806 3689 50858 3695
rect 50806 3631 50858 3637
rect 50348 3358 50644 3378
rect 50404 3356 50428 3358
rect 50484 3356 50508 3358
rect 50564 3356 50588 3358
rect 50426 3304 50428 3356
rect 50490 3304 50502 3356
rect 50564 3304 50566 3356
rect 50404 3302 50428 3304
rect 50484 3302 50508 3304
rect 50564 3302 50588 3304
rect 50348 3282 50644 3302
rect 50242 2576 50366 2604
rect 50338 800 50366 2576
rect 50722 1864 50750 3631
rect 50434 1836 50750 1864
rect 50434 800 50462 1836
rect 50518 1765 50570 1771
rect 50518 1707 50570 1713
rect 50530 800 50558 1707
rect 50710 1691 50762 1697
rect 50710 1633 50762 1639
rect 50722 800 50750 1633
rect 50818 800 50846 3631
rect 50914 1697 50942 4963
rect 50998 4281 51050 4287
rect 50998 4223 51050 4229
rect 50902 1691 50954 1697
rect 50902 1633 50954 1639
rect 50902 1543 50954 1549
rect 50902 1485 50954 1491
rect 50914 800 50942 1485
rect 51010 800 51038 4223
rect 51106 1771 51134 6073
rect 51382 3911 51434 3917
rect 51382 3853 51434 3859
rect 51286 3689 51338 3695
rect 51202 3649 51286 3677
rect 51094 1765 51146 1771
rect 51094 1707 51146 1713
rect 51202 800 51230 3649
rect 51286 3631 51338 3637
rect 51286 3541 51338 3547
rect 51286 3483 51338 3489
rect 51298 800 51326 3483
rect 51394 800 51422 3853
rect 51490 3547 51518 6887
rect 51574 6205 51626 6211
rect 51574 6147 51626 6153
rect 51478 3541 51530 3547
rect 51478 3483 51530 3489
rect 51478 3023 51530 3029
rect 51478 2965 51530 2971
rect 51490 800 51518 2965
rect 51586 1549 51614 6147
rect 51778 5120 51806 7405
rect 52258 6433 52286 12946
rect 52342 8573 52394 8579
rect 52450 8547 52478 49363
rect 52534 24927 52586 24933
rect 52534 24869 52586 24875
rect 52342 8515 52394 8521
rect 52436 8538 52492 8547
rect 52354 8376 52382 8515
rect 52436 8473 52492 8482
rect 52546 8376 52574 24869
rect 52642 12974 52670 56171
rect 53590 50753 53642 50759
rect 53590 50695 53642 50701
rect 53206 39209 53258 39215
rect 53206 39151 53258 39157
rect 53014 20117 53066 20123
rect 53014 20059 53066 20065
rect 52642 12946 52766 12974
rect 52630 9461 52682 9467
rect 52630 9403 52682 9409
rect 52642 9245 52670 9403
rect 52630 9239 52682 9245
rect 52630 9181 52682 9187
rect 52354 8348 52574 8376
rect 52342 7463 52394 7469
rect 52342 7405 52394 7411
rect 52246 6427 52298 6433
rect 52246 6369 52298 6375
rect 52246 6279 52298 6285
rect 52246 6221 52298 6227
rect 52150 5687 52202 5693
rect 52150 5629 52202 5635
rect 51682 5092 51806 5120
rect 51574 1543 51626 1549
rect 51574 1485 51626 1491
rect 51682 800 51710 5092
rect 51862 5021 51914 5027
rect 51862 4963 51914 4969
rect 51958 5021 52010 5027
rect 51958 4963 52010 4969
rect 51874 3917 51902 4963
rect 51862 3911 51914 3917
rect 51862 3853 51914 3859
rect 51970 3788 51998 4963
rect 51778 3760 51998 3788
rect 51778 800 51806 3760
rect 52054 3689 52106 3695
rect 51970 3649 52054 3677
rect 51970 1864 51998 3649
rect 52054 3631 52106 3637
rect 52054 3541 52106 3547
rect 52054 3483 52106 3489
rect 51874 1836 51998 1864
rect 51874 800 51902 1836
rect 52066 800 52094 3483
rect 52162 800 52190 5629
rect 52258 3103 52286 6221
rect 52246 3097 52298 3103
rect 52246 3039 52298 3045
rect 52246 2949 52298 2955
rect 52246 2891 52298 2897
rect 52258 800 52286 2891
rect 52354 800 52382 7405
rect 52738 7215 52766 12946
rect 52916 8390 52972 8399
rect 52916 8325 52918 8334
rect 52970 8325 52972 8334
rect 52918 8293 52970 8299
rect 53026 7913 53054 20059
rect 53110 8203 53162 8209
rect 53110 8145 53162 8151
rect 53014 7907 53066 7913
rect 53014 7849 53066 7855
rect 52822 7759 52874 7765
rect 52822 7701 52874 7707
rect 52724 7206 52780 7215
rect 52724 7141 52780 7150
rect 52726 6945 52778 6951
rect 52726 6887 52778 6893
rect 52534 5687 52586 5693
rect 52534 5629 52586 5635
rect 52546 800 52574 5629
rect 52630 4355 52682 4361
rect 52630 4297 52682 4303
rect 52642 800 52670 4297
rect 52738 3547 52766 6887
rect 52726 3541 52778 3547
rect 52726 3483 52778 3489
rect 52834 2894 52862 7701
rect 53014 4281 53066 4287
rect 53014 4223 53066 4229
rect 52738 2866 52862 2894
rect 52918 2949 52970 2955
rect 52918 2891 52970 2897
rect 52738 800 52766 2866
rect 52930 800 52958 2891
rect 53026 800 53054 4223
rect 53122 800 53150 8145
rect 53218 7691 53246 39151
rect 53398 14493 53450 14499
rect 53398 14435 53450 14441
rect 53410 9023 53438 14435
rect 53398 9017 53450 9023
rect 53398 8959 53450 8965
rect 53494 8277 53546 8283
rect 53494 8219 53546 8225
rect 53206 7685 53258 7691
rect 53206 7627 53258 7633
rect 53302 5021 53354 5027
rect 53302 4963 53354 4969
rect 53314 2900 53342 4963
rect 53398 3689 53450 3695
rect 53398 3631 53450 3637
rect 53218 2872 53342 2900
rect 53218 800 53246 2872
rect 53410 800 53438 3631
rect 53506 800 53534 8219
rect 53602 6919 53630 50695
rect 53698 19827 53726 56171
rect 53878 42761 53930 42767
rect 53878 42703 53930 42709
rect 53890 42545 53918 42703
rect 53878 42539 53930 42545
rect 53878 42481 53930 42487
rect 53986 20567 54014 56689
rect 54370 56531 54398 59200
rect 54550 57413 54602 57419
rect 54550 57355 54602 57361
rect 54358 56525 54410 56531
rect 54358 56467 54410 56473
rect 54562 56309 54590 57355
rect 54946 56531 54974 59200
rect 55426 56901 55454 59200
rect 55414 56895 55466 56901
rect 55414 56837 55466 56843
rect 55318 56821 55370 56827
rect 55318 56763 55370 56769
rect 54934 56525 54986 56531
rect 54934 56467 54986 56473
rect 55126 56451 55178 56457
rect 55126 56393 55178 56399
rect 54550 56303 54602 56309
rect 54550 56245 54602 56251
rect 55030 56303 55082 56309
rect 55030 56245 55082 56251
rect 54646 29441 54698 29447
rect 54646 29383 54698 29389
rect 53974 20561 54026 20567
rect 53974 20503 54026 20509
rect 53686 19821 53738 19827
rect 53686 19763 53738 19769
rect 54262 9609 54314 9615
rect 54262 9551 54314 9557
rect 54454 9609 54506 9615
rect 54454 9551 54506 9557
rect 53878 8795 53930 8801
rect 53878 8737 53930 8743
rect 53588 6910 53644 6919
rect 53588 6845 53644 6854
rect 53686 5687 53738 5693
rect 53686 5629 53738 5635
rect 53590 5613 53642 5619
rect 53590 5555 53642 5561
rect 53602 800 53630 5555
rect 53698 2955 53726 5629
rect 53782 3023 53834 3029
rect 53782 2965 53834 2971
rect 53686 2949 53738 2955
rect 53686 2891 53738 2897
rect 53794 1568 53822 2965
rect 53698 1540 53822 1568
rect 53698 800 53726 1540
rect 53890 800 53918 8737
rect 54070 8277 54122 8283
rect 54070 8219 54122 8225
rect 54082 7247 54110 8219
rect 54070 7241 54122 7247
rect 54070 7183 54122 7189
rect 53974 6353 54026 6359
rect 53974 6295 54026 6301
rect 53986 800 54014 6295
rect 54070 4355 54122 4361
rect 54070 4297 54122 4303
rect 54082 800 54110 4297
rect 54274 800 54302 9551
rect 54466 9171 54494 9551
rect 54454 9165 54506 9171
rect 54454 9107 54506 9113
rect 54658 9097 54686 29383
rect 54742 11607 54794 11613
rect 54742 11549 54794 11555
rect 54646 9091 54698 9097
rect 54646 9033 54698 9039
rect 54550 9017 54602 9023
rect 54550 8959 54602 8965
rect 54358 6279 54410 6285
rect 54358 6221 54410 6227
rect 54370 800 54398 6221
rect 54454 3541 54506 3547
rect 54454 3483 54506 3489
rect 54466 800 54494 3483
rect 54562 800 54590 8959
rect 54754 8135 54782 11549
rect 54934 9905 54986 9911
rect 54934 9847 54986 9853
rect 54742 8129 54794 8135
rect 54742 8071 54794 8077
rect 54742 7019 54794 7025
rect 54742 6961 54794 6967
rect 54754 800 54782 6961
rect 54838 2949 54890 2955
rect 54838 2891 54890 2897
rect 54850 800 54878 2891
rect 54946 800 54974 9847
rect 55042 5915 55070 56245
rect 55138 25895 55166 56393
rect 55330 56235 55358 56763
rect 55510 56747 55562 56753
rect 55510 56689 55562 56695
rect 55522 56383 55550 56689
rect 56002 56531 56030 59200
rect 55990 56525 56042 56531
rect 55990 56467 56042 56473
rect 55510 56377 55562 56383
rect 55510 56319 55562 56325
rect 55318 56229 55370 56235
rect 55318 56171 55370 56177
rect 56482 55717 56510 59200
rect 57058 56901 57086 59200
rect 57046 56895 57098 56901
rect 57046 56837 57098 56843
rect 56950 56229 57002 56235
rect 56950 56171 57002 56177
rect 56470 55711 56522 55717
rect 56470 55653 56522 55659
rect 56566 55563 56618 55569
rect 56566 55505 56618 55511
rect 55606 55045 55658 55051
rect 55606 54987 55658 54993
rect 55510 29663 55562 29669
rect 55510 29605 55562 29611
rect 55522 29225 55550 29605
rect 55510 29219 55562 29225
rect 55510 29161 55562 29167
rect 55126 25889 55178 25895
rect 55126 25831 55178 25837
rect 55318 9905 55370 9911
rect 55318 9847 55370 9853
rect 55126 6205 55178 6211
rect 55126 6147 55178 6153
rect 55030 5909 55082 5915
rect 55030 5851 55082 5857
rect 55138 3196 55166 6147
rect 55222 3467 55274 3473
rect 55222 3409 55274 3415
rect 55042 3168 55166 3196
rect 55042 800 55070 3168
rect 55234 800 55262 3409
rect 55330 800 55358 9847
rect 55618 9837 55646 54987
rect 56374 54083 56426 54089
rect 56374 54025 56426 54031
rect 55894 37433 55946 37439
rect 55894 37375 55946 37381
rect 55702 29441 55754 29447
rect 55702 29383 55754 29389
rect 55714 10355 55742 29383
rect 55906 10429 55934 37375
rect 56278 13013 56330 13019
rect 56278 12955 56330 12961
rect 55894 10423 55946 10429
rect 55894 10365 55946 10371
rect 55702 10349 55754 10355
rect 55702 10291 55754 10297
rect 55702 10127 55754 10133
rect 55702 10069 55754 10075
rect 56086 10127 56138 10133
rect 56086 10069 56138 10075
rect 55606 9831 55658 9837
rect 55606 9773 55658 9779
rect 55414 7019 55466 7025
rect 55414 6961 55466 6967
rect 55426 800 55454 6961
rect 55606 4355 55658 4361
rect 55606 4297 55658 4303
rect 55618 800 55646 4297
rect 55714 800 55742 10069
rect 55990 8869 56042 8875
rect 55990 8811 56042 8817
rect 55798 7685 55850 7691
rect 55798 7627 55850 7633
rect 55810 800 55838 7627
rect 56002 4213 56030 8811
rect 55990 4207 56042 4213
rect 55990 4149 56042 4155
rect 55894 3763 55946 3769
rect 55894 3705 55946 3711
rect 55906 800 55934 3705
rect 56098 800 56126 10069
rect 56182 7685 56234 7691
rect 56182 7627 56234 7633
rect 56194 800 56222 7627
rect 56290 7617 56318 12955
rect 56386 7807 56414 54025
rect 56470 38765 56522 38771
rect 56470 38707 56522 38713
rect 56482 10577 56510 38707
rect 56578 33221 56606 55505
rect 56566 33215 56618 33221
rect 56566 33157 56618 33163
rect 56962 13241 56990 56171
rect 57538 55717 57566 59200
rect 57526 55711 57578 55717
rect 57526 55653 57578 55659
rect 57430 55563 57482 55569
rect 57430 55505 57482 55511
rect 57334 42095 57386 42101
rect 57334 42037 57386 42043
rect 56950 13235 57002 13241
rect 56950 13177 57002 13183
rect 57346 12575 57374 42037
rect 57334 12569 57386 12575
rect 57334 12511 57386 12517
rect 57442 12279 57470 55505
rect 58114 54385 58142 59200
rect 58594 56309 58622 59200
rect 58582 56303 58634 56309
rect 58582 56245 58634 56251
rect 59170 55199 59198 59200
rect 59158 55193 59210 55199
rect 59158 55135 59210 55141
rect 58102 54379 58154 54385
rect 58102 54321 58154 54327
rect 57814 54231 57866 54237
rect 57814 54173 57866 54179
rect 57718 53417 57770 53423
rect 57718 53359 57770 53365
rect 57622 50087 57674 50093
rect 57622 50029 57674 50035
rect 57634 49871 57662 50029
rect 57622 49865 57674 49871
rect 57622 49807 57674 49813
rect 57730 21159 57758 53359
rect 57718 21153 57770 21159
rect 57718 21095 57770 21101
rect 57430 12273 57482 12279
rect 57430 12215 57482 12221
rect 57526 12199 57578 12205
rect 57526 12141 57578 12147
rect 57142 11459 57194 11465
rect 57142 11401 57194 11407
rect 56758 10941 56810 10947
rect 56758 10883 56810 10889
rect 56566 10867 56618 10873
rect 56566 10809 56618 10815
rect 56470 10571 56522 10577
rect 56470 10513 56522 10519
rect 56470 10275 56522 10281
rect 56470 10217 56522 10223
rect 56372 7798 56428 7807
rect 56372 7733 56428 7742
rect 56278 7611 56330 7617
rect 56278 7553 56330 7559
rect 56278 6945 56330 6951
rect 56278 6887 56330 6893
rect 56290 3917 56318 6887
rect 56374 6427 56426 6433
rect 56374 6369 56426 6375
rect 56278 3911 56330 3917
rect 56278 3853 56330 3859
rect 56278 3541 56330 3547
rect 56278 3483 56330 3489
rect 56290 800 56318 3483
rect 56386 3251 56414 6369
rect 56374 3245 56426 3251
rect 56374 3187 56426 3193
rect 56374 3097 56426 3103
rect 56372 3062 56374 3071
rect 56426 3062 56428 3071
rect 56372 2997 56428 3006
rect 56482 800 56510 10217
rect 56578 4995 56606 10809
rect 56564 4986 56620 4995
rect 56564 4921 56620 4930
rect 56770 4824 56798 10883
rect 56950 8351 57002 8357
rect 56950 8293 57002 8299
rect 56854 7685 56906 7691
rect 56854 7627 56906 7633
rect 56578 4796 56798 4824
rect 56578 4287 56606 4796
rect 56660 4690 56716 4699
rect 56660 4625 56716 4634
rect 56566 4281 56618 4287
rect 56566 4223 56618 4229
rect 56674 3640 56702 4625
rect 56758 4503 56810 4509
rect 56758 4445 56810 4451
rect 56770 3843 56798 4445
rect 56758 3837 56810 3843
rect 56758 3779 56810 3785
rect 56566 3615 56618 3621
rect 56674 3612 56798 3640
rect 56866 3621 56894 7627
rect 56566 3557 56618 3563
rect 56578 800 56606 3557
rect 56662 3023 56714 3029
rect 56662 2965 56714 2971
rect 56674 800 56702 2965
rect 56770 800 56798 3612
rect 56854 3615 56906 3621
rect 56854 3557 56906 3563
rect 56962 800 56990 8293
rect 57046 5021 57098 5027
rect 57046 4963 57098 4969
rect 57058 800 57086 4963
rect 57154 800 57182 11401
rect 57238 9017 57290 9023
rect 57238 8959 57290 8965
rect 57250 800 57278 8959
rect 57334 8943 57386 8949
rect 57334 8885 57386 8891
rect 57346 4509 57374 8885
rect 57430 5687 57482 5693
rect 57430 5629 57482 5635
rect 57334 4503 57386 4509
rect 57334 4445 57386 4451
rect 57334 4355 57386 4361
rect 57334 4297 57386 4303
rect 57346 3029 57374 4297
rect 57334 3023 57386 3029
rect 57334 2965 57386 2971
rect 57442 800 57470 5629
rect 57538 800 57566 12141
rect 57622 9683 57674 9689
rect 57622 9625 57674 9631
rect 57634 800 57662 9625
rect 57826 9541 57854 54173
rect 59650 53867 59678 59200
rect 59638 53861 59690 53867
rect 59638 53803 59690 53809
rect 58198 11607 58250 11613
rect 58198 11549 58250 11555
rect 57814 9535 57866 9541
rect 57814 9477 57866 9483
rect 58102 6353 58154 6359
rect 58102 6295 58154 6301
rect 57814 4947 57866 4953
rect 57814 4889 57866 4895
rect 57826 800 57854 4889
rect 57910 4207 57962 4213
rect 57910 4149 57962 4155
rect 57922 800 57950 4149
rect 58006 3245 58058 3251
rect 58006 3187 58058 3193
rect 58018 800 58046 3187
rect 58114 800 58142 6295
rect 58210 3695 58238 11549
rect 58582 10201 58634 10207
rect 58582 10143 58634 10149
rect 58390 8277 58442 8283
rect 58390 8219 58442 8225
rect 58294 4281 58346 4287
rect 58294 4223 58346 4229
rect 58198 3689 58250 3695
rect 58198 3631 58250 3637
rect 58306 800 58334 4223
rect 58402 800 58430 8219
rect 58486 7019 58538 7025
rect 58486 6961 58538 6967
rect 58498 800 58526 6961
rect 58594 800 58622 10143
rect 58966 8573 59018 8579
rect 58966 8515 59018 8521
rect 58774 7759 58826 7765
rect 58774 7701 58826 7707
rect 58786 800 58814 7701
rect 58870 6279 58922 6285
rect 58870 6221 58922 6227
rect 58882 800 58910 6221
rect 58978 800 59006 8515
rect 59830 8203 59882 8209
rect 59830 8145 59882 8151
rect 59350 7833 59402 7839
rect 59350 7775 59402 7781
rect 59254 4873 59306 4879
rect 59254 4815 59306 4821
rect 59158 3763 59210 3769
rect 59158 3705 59210 3711
rect 59170 800 59198 3705
rect 59266 800 59294 4815
rect 59362 800 59390 7775
rect 59638 5613 59690 5619
rect 59638 5555 59690 5561
rect 59446 3837 59498 3843
rect 59446 3779 59498 3785
rect 59458 800 59486 3779
rect 59650 800 59678 5555
rect 59734 3689 59786 3695
rect 59734 3631 59786 3637
rect 59746 800 59774 3631
rect 59842 800 59870 8145
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1364 0 1420 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2708 0 2764 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3188 0 3244 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 4052 0 4108 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4532 0 4588 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4916 0 4972 800
rect 5012 0 5068 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5396 0 5452 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5876 0 5932 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6260 0 6316 800
rect 6356 0 6412 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6740 0 6796 800
rect 6836 0 6892 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7220 0 7276 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7604 0 7660 800
rect 7700 0 7756 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 8084 0 8140 800
rect 8180 0 8236 800
rect 8276 0 8332 800
rect 8468 0 8524 800
rect 8564 0 8620 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8948 0 9004 800
rect 9044 0 9100 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9428 0 9484 800
rect 9524 0 9580 800
rect 9620 0 9676 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10004 0 10060 800
rect 10100 0 10156 800
rect 10292 0 10348 800
rect 10388 0 10444 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10772 0 10828 800
rect 10868 0 10924 800
rect 10964 0 11020 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11348 0 11404 800
rect 11444 0 11500 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11828 0 11884 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12212 0 12268 800
rect 12308 0 12364 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12692 0 12748 800
rect 12788 0 12844 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13172 0 13228 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13652 0 13708 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14036 0 14092 800
rect 14132 0 14188 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14516 0 14572 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 14996 0 15052 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15380 0 15436 800
rect 15476 0 15532 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15860 0 15916 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16340 0 16396 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17204 0 17260 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17684 0 17740 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19028 0 19084 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20468 0 20524 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21812 0 21868 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22292 0 22348 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23156 0 23212 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23636 0 23692 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 24020 0 24076 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24500 0 24556 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24980 0 25036 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25364 0 25420 800
rect 25460 0 25516 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25844 0 25900 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26324 0 26380 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26708 0 26764 800
rect 26804 0 26860 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27188 0 27244 800
rect 27284 0 27340 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27668 0 27724 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 28052 0 28108 800
rect 28148 0 28204 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28532 0 28588 800
rect 28628 0 28684 800
rect 28724 0 28780 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29108 0 29164 800
rect 29204 0 29260 800
rect 29396 0 29452 800
rect 29492 0 29548 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29876 0 29932 800
rect 29972 0 30028 800
rect 30068 0 30124 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30452 0 30508 800
rect 30548 0 30604 800
rect 30740 0 30796 800
rect 30836 0 30892 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31220 0 31276 800
rect 31316 0 31372 800
rect 31412 0 31468 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31796 0 31852 800
rect 31892 0 31948 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32276 0 32332 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32660 0 32716 800
rect 32756 0 32812 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33140 0 33196 800
rect 33236 0 33292 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33620 0 33676 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34100 0 34156 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34484 0 34540 800
rect 34580 0 34636 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 34964 0 35020 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35444 0 35500 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36308 0 36364 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36788 0 36844 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37652 0 37708 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38132 0 38188 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39476 0 39532 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40916 0 40972 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42260 0 42316 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42740 0 42796 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43604 0 43660 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 44084 0 44140 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44468 0 44524 800
rect 44564 0 44620 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44948 0 45004 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45428 0 45484 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45812 0 45868 800
rect 45908 0 45964 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46292 0 46348 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46772 0 46828 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47156 0 47212 800
rect 47252 0 47308 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47636 0 47692 800
rect 47732 0 47788 800
rect 47828 0 47884 800
rect 48020 0 48076 800
rect 48116 0 48172 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48500 0 48556 800
rect 48596 0 48652 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48980 0 49036 800
rect 49076 0 49132 800
rect 49172 0 49228 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49556 0 49612 800
rect 49652 0 49708 800
rect 49844 0 49900 800
rect 49940 0 49996 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50324 0 50380 800
rect 50420 0 50476 800
rect 50516 0 50572 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50900 0 50956 800
rect 50996 0 51052 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51380 0 51436 800
rect 51476 0 51532 800
rect 51668 0 51724 800
rect 51764 0 51820 800
rect 51860 0 51916 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52244 0 52300 800
rect 52340 0 52396 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52724 0 52780 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53108 0 53164 800
rect 53204 0 53260 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53588 0 53644 800
rect 53684 0 53740 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54068 0 54124 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54548 0 54604 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 54932 0 54988 800
rect 55028 0 55084 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55412 0 55468 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55892 0 55948 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56756 0 56812 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57236 0 57292 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58580 0 58636 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< via2 >>
rect 2228 8186 2284 8242
rect 2516 7611 2572 7650
rect 2516 7594 2518 7611
rect 2518 7594 2570 7611
rect 2570 7594 2572 7611
rect 4268 57302 4324 57304
rect 4348 57302 4404 57304
rect 4428 57302 4484 57304
rect 4508 57302 4564 57304
rect 4268 57250 4294 57302
rect 4294 57250 4324 57302
rect 4348 57250 4358 57302
rect 4358 57250 4404 57302
rect 4428 57250 4474 57302
rect 4474 57250 4484 57302
rect 4508 57250 4538 57302
rect 4538 57250 4564 57302
rect 4268 57248 4324 57250
rect 4348 57248 4404 57250
rect 4428 57248 4484 57250
rect 4508 57248 4564 57250
rect 4268 55970 4324 55972
rect 4348 55970 4404 55972
rect 4428 55970 4484 55972
rect 4508 55970 4564 55972
rect 4268 55918 4294 55970
rect 4294 55918 4324 55970
rect 4348 55918 4358 55970
rect 4358 55918 4404 55970
rect 4428 55918 4474 55970
rect 4474 55918 4484 55970
rect 4508 55918 4538 55970
rect 4538 55918 4564 55970
rect 4268 55916 4324 55918
rect 4348 55916 4404 55918
rect 4428 55916 4484 55918
rect 4508 55916 4564 55918
rect 4268 54638 4324 54640
rect 4348 54638 4404 54640
rect 4428 54638 4484 54640
rect 4508 54638 4564 54640
rect 4268 54586 4294 54638
rect 4294 54586 4324 54638
rect 4348 54586 4358 54638
rect 4358 54586 4404 54638
rect 4428 54586 4474 54638
rect 4474 54586 4484 54638
rect 4508 54586 4538 54638
rect 4538 54586 4564 54638
rect 4268 54584 4324 54586
rect 4348 54584 4404 54586
rect 4428 54584 4484 54586
rect 4508 54584 4564 54586
rect 4268 53306 4324 53308
rect 4348 53306 4404 53308
rect 4428 53306 4484 53308
rect 4508 53306 4564 53308
rect 4268 53254 4294 53306
rect 4294 53254 4324 53306
rect 4348 53254 4358 53306
rect 4358 53254 4404 53306
rect 4428 53254 4474 53306
rect 4474 53254 4484 53306
rect 4508 53254 4538 53306
rect 4538 53254 4564 53306
rect 4268 53252 4324 53254
rect 4348 53252 4404 53254
rect 4428 53252 4484 53254
rect 4508 53252 4564 53254
rect 4268 51974 4324 51976
rect 4348 51974 4404 51976
rect 4428 51974 4484 51976
rect 4508 51974 4564 51976
rect 4268 51922 4294 51974
rect 4294 51922 4324 51974
rect 4348 51922 4358 51974
rect 4358 51922 4404 51974
rect 4428 51922 4474 51974
rect 4474 51922 4484 51974
rect 4508 51922 4538 51974
rect 4538 51922 4564 51974
rect 4268 51920 4324 51922
rect 4348 51920 4404 51922
rect 4428 51920 4484 51922
rect 4508 51920 4564 51922
rect 4268 50642 4324 50644
rect 4348 50642 4404 50644
rect 4428 50642 4484 50644
rect 4508 50642 4564 50644
rect 4268 50590 4294 50642
rect 4294 50590 4324 50642
rect 4348 50590 4358 50642
rect 4358 50590 4404 50642
rect 4428 50590 4474 50642
rect 4474 50590 4484 50642
rect 4508 50590 4538 50642
rect 4538 50590 4564 50642
rect 4268 50588 4324 50590
rect 4348 50588 4404 50590
rect 4428 50588 4484 50590
rect 4508 50588 4564 50590
rect 4268 49310 4324 49312
rect 4348 49310 4404 49312
rect 4428 49310 4484 49312
rect 4508 49310 4564 49312
rect 4268 49258 4294 49310
rect 4294 49258 4324 49310
rect 4348 49258 4358 49310
rect 4358 49258 4404 49310
rect 4428 49258 4474 49310
rect 4474 49258 4484 49310
rect 4508 49258 4538 49310
rect 4538 49258 4564 49310
rect 4268 49256 4324 49258
rect 4348 49256 4404 49258
rect 4428 49256 4484 49258
rect 4508 49256 4564 49258
rect 4268 47978 4324 47980
rect 4348 47978 4404 47980
rect 4428 47978 4484 47980
rect 4508 47978 4564 47980
rect 4268 47926 4294 47978
rect 4294 47926 4324 47978
rect 4348 47926 4358 47978
rect 4358 47926 4404 47978
rect 4428 47926 4474 47978
rect 4474 47926 4484 47978
rect 4508 47926 4538 47978
rect 4538 47926 4564 47978
rect 4268 47924 4324 47926
rect 4348 47924 4404 47926
rect 4428 47924 4484 47926
rect 4508 47924 4564 47926
rect 4268 46646 4324 46648
rect 4348 46646 4404 46648
rect 4428 46646 4484 46648
rect 4508 46646 4564 46648
rect 4268 46594 4294 46646
rect 4294 46594 4324 46646
rect 4348 46594 4358 46646
rect 4358 46594 4404 46646
rect 4428 46594 4474 46646
rect 4474 46594 4484 46646
rect 4508 46594 4538 46646
rect 4538 46594 4564 46646
rect 4268 46592 4324 46594
rect 4348 46592 4404 46594
rect 4428 46592 4484 46594
rect 4508 46592 4564 46594
rect 4268 45314 4324 45316
rect 4348 45314 4404 45316
rect 4428 45314 4484 45316
rect 4508 45314 4564 45316
rect 4268 45262 4294 45314
rect 4294 45262 4324 45314
rect 4348 45262 4358 45314
rect 4358 45262 4404 45314
rect 4428 45262 4474 45314
rect 4474 45262 4484 45314
rect 4508 45262 4538 45314
rect 4538 45262 4564 45314
rect 4268 45260 4324 45262
rect 4348 45260 4404 45262
rect 4428 45260 4484 45262
rect 4508 45260 4564 45262
rect 4268 43982 4324 43984
rect 4348 43982 4404 43984
rect 4428 43982 4484 43984
rect 4508 43982 4564 43984
rect 4268 43930 4294 43982
rect 4294 43930 4324 43982
rect 4348 43930 4358 43982
rect 4358 43930 4404 43982
rect 4428 43930 4474 43982
rect 4474 43930 4484 43982
rect 4508 43930 4538 43982
rect 4538 43930 4564 43982
rect 4268 43928 4324 43930
rect 4348 43928 4404 43930
rect 4428 43928 4484 43930
rect 4508 43928 4564 43930
rect 4268 42650 4324 42652
rect 4348 42650 4404 42652
rect 4428 42650 4484 42652
rect 4508 42650 4564 42652
rect 4268 42598 4294 42650
rect 4294 42598 4324 42650
rect 4348 42598 4358 42650
rect 4358 42598 4404 42650
rect 4428 42598 4474 42650
rect 4474 42598 4484 42650
rect 4508 42598 4538 42650
rect 4538 42598 4564 42650
rect 4268 42596 4324 42598
rect 4348 42596 4404 42598
rect 4428 42596 4484 42598
rect 4508 42596 4564 42598
rect 4268 41318 4324 41320
rect 4348 41318 4404 41320
rect 4428 41318 4484 41320
rect 4508 41318 4564 41320
rect 4268 41266 4294 41318
rect 4294 41266 4324 41318
rect 4348 41266 4358 41318
rect 4358 41266 4404 41318
rect 4428 41266 4474 41318
rect 4474 41266 4484 41318
rect 4508 41266 4538 41318
rect 4538 41266 4564 41318
rect 4268 41264 4324 41266
rect 4348 41264 4404 41266
rect 4428 41264 4484 41266
rect 4508 41264 4564 41266
rect 4268 39986 4324 39988
rect 4348 39986 4404 39988
rect 4428 39986 4484 39988
rect 4508 39986 4564 39988
rect 4268 39934 4294 39986
rect 4294 39934 4324 39986
rect 4348 39934 4358 39986
rect 4358 39934 4404 39986
rect 4428 39934 4474 39986
rect 4474 39934 4484 39986
rect 4508 39934 4538 39986
rect 4538 39934 4564 39986
rect 4268 39932 4324 39934
rect 4348 39932 4404 39934
rect 4428 39932 4484 39934
rect 4508 39932 4564 39934
rect 4268 38654 4324 38656
rect 4348 38654 4404 38656
rect 4428 38654 4484 38656
rect 4508 38654 4564 38656
rect 4268 38602 4294 38654
rect 4294 38602 4324 38654
rect 4348 38602 4358 38654
rect 4358 38602 4404 38654
rect 4428 38602 4474 38654
rect 4474 38602 4484 38654
rect 4508 38602 4538 38654
rect 4538 38602 4564 38654
rect 4268 38600 4324 38602
rect 4348 38600 4404 38602
rect 4428 38600 4484 38602
rect 4508 38600 4564 38602
rect 4268 37322 4324 37324
rect 4348 37322 4404 37324
rect 4428 37322 4484 37324
rect 4508 37322 4564 37324
rect 4268 37270 4294 37322
rect 4294 37270 4324 37322
rect 4348 37270 4358 37322
rect 4358 37270 4404 37322
rect 4428 37270 4474 37322
rect 4474 37270 4484 37322
rect 4508 37270 4538 37322
rect 4538 37270 4564 37322
rect 4268 37268 4324 37270
rect 4348 37268 4404 37270
rect 4428 37268 4484 37270
rect 4508 37268 4564 37270
rect 4268 35990 4324 35992
rect 4348 35990 4404 35992
rect 4428 35990 4484 35992
rect 4508 35990 4564 35992
rect 4268 35938 4294 35990
rect 4294 35938 4324 35990
rect 4348 35938 4358 35990
rect 4358 35938 4404 35990
rect 4428 35938 4474 35990
rect 4474 35938 4484 35990
rect 4508 35938 4538 35990
rect 4538 35938 4564 35990
rect 4268 35936 4324 35938
rect 4348 35936 4404 35938
rect 4428 35936 4484 35938
rect 4508 35936 4564 35938
rect 4268 34658 4324 34660
rect 4348 34658 4404 34660
rect 4428 34658 4484 34660
rect 4508 34658 4564 34660
rect 4268 34606 4294 34658
rect 4294 34606 4324 34658
rect 4348 34606 4358 34658
rect 4358 34606 4404 34658
rect 4428 34606 4474 34658
rect 4474 34606 4484 34658
rect 4508 34606 4538 34658
rect 4538 34606 4564 34658
rect 4268 34604 4324 34606
rect 4348 34604 4404 34606
rect 4428 34604 4484 34606
rect 4508 34604 4564 34606
rect 4268 33326 4324 33328
rect 4348 33326 4404 33328
rect 4428 33326 4484 33328
rect 4508 33326 4564 33328
rect 4268 33274 4294 33326
rect 4294 33274 4324 33326
rect 4348 33274 4358 33326
rect 4358 33274 4404 33326
rect 4428 33274 4474 33326
rect 4474 33274 4484 33326
rect 4508 33274 4538 33326
rect 4538 33274 4564 33326
rect 4268 33272 4324 33274
rect 4348 33272 4404 33274
rect 4428 33272 4484 33274
rect 4508 33272 4564 33274
rect 4268 31994 4324 31996
rect 4348 31994 4404 31996
rect 4428 31994 4484 31996
rect 4508 31994 4564 31996
rect 4268 31942 4294 31994
rect 4294 31942 4324 31994
rect 4348 31942 4358 31994
rect 4358 31942 4404 31994
rect 4428 31942 4474 31994
rect 4474 31942 4484 31994
rect 4508 31942 4538 31994
rect 4538 31942 4564 31994
rect 4268 31940 4324 31942
rect 4348 31940 4404 31942
rect 4428 31940 4484 31942
rect 4508 31940 4564 31942
rect 4268 30662 4324 30664
rect 4348 30662 4404 30664
rect 4428 30662 4484 30664
rect 4508 30662 4564 30664
rect 4268 30610 4294 30662
rect 4294 30610 4324 30662
rect 4348 30610 4358 30662
rect 4358 30610 4404 30662
rect 4428 30610 4474 30662
rect 4474 30610 4484 30662
rect 4508 30610 4538 30662
rect 4538 30610 4564 30662
rect 4268 30608 4324 30610
rect 4348 30608 4404 30610
rect 4428 30608 4484 30610
rect 4508 30608 4564 30610
rect 4268 29330 4324 29332
rect 4348 29330 4404 29332
rect 4428 29330 4484 29332
rect 4508 29330 4564 29332
rect 4268 29278 4294 29330
rect 4294 29278 4324 29330
rect 4348 29278 4358 29330
rect 4358 29278 4404 29330
rect 4428 29278 4474 29330
rect 4474 29278 4484 29330
rect 4508 29278 4538 29330
rect 4538 29278 4564 29330
rect 4268 29276 4324 29278
rect 4348 29276 4404 29278
rect 4428 29276 4484 29278
rect 4508 29276 4564 29278
rect 4268 27998 4324 28000
rect 4348 27998 4404 28000
rect 4428 27998 4484 28000
rect 4508 27998 4564 28000
rect 4268 27946 4294 27998
rect 4294 27946 4324 27998
rect 4348 27946 4358 27998
rect 4358 27946 4404 27998
rect 4428 27946 4474 27998
rect 4474 27946 4484 27998
rect 4508 27946 4538 27998
rect 4538 27946 4564 27998
rect 4268 27944 4324 27946
rect 4348 27944 4404 27946
rect 4428 27944 4484 27946
rect 4508 27944 4564 27946
rect 4268 26666 4324 26668
rect 4348 26666 4404 26668
rect 4428 26666 4484 26668
rect 4508 26666 4564 26668
rect 4268 26614 4294 26666
rect 4294 26614 4324 26666
rect 4348 26614 4358 26666
rect 4358 26614 4404 26666
rect 4428 26614 4474 26666
rect 4474 26614 4484 26666
rect 4508 26614 4538 26666
rect 4538 26614 4564 26666
rect 4268 26612 4324 26614
rect 4348 26612 4404 26614
rect 4428 26612 4484 26614
rect 4508 26612 4564 26614
rect 4268 25334 4324 25336
rect 4348 25334 4404 25336
rect 4428 25334 4484 25336
rect 4508 25334 4564 25336
rect 4268 25282 4294 25334
rect 4294 25282 4324 25334
rect 4348 25282 4358 25334
rect 4358 25282 4404 25334
rect 4428 25282 4474 25334
rect 4474 25282 4484 25334
rect 4508 25282 4538 25334
rect 4538 25282 4564 25334
rect 4268 25280 4324 25282
rect 4348 25280 4404 25282
rect 4428 25280 4484 25282
rect 4508 25280 4564 25282
rect 4268 24002 4324 24004
rect 4348 24002 4404 24004
rect 4428 24002 4484 24004
rect 4508 24002 4564 24004
rect 4268 23950 4294 24002
rect 4294 23950 4324 24002
rect 4348 23950 4358 24002
rect 4358 23950 4404 24002
rect 4428 23950 4474 24002
rect 4474 23950 4484 24002
rect 4508 23950 4538 24002
rect 4538 23950 4564 24002
rect 4268 23948 4324 23950
rect 4348 23948 4404 23950
rect 4428 23948 4484 23950
rect 4508 23948 4564 23950
rect 4268 22670 4324 22672
rect 4348 22670 4404 22672
rect 4428 22670 4484 22672
rect 4508 22670 4564 22672
rect 4268 22618 4294 22670
rect 4294 22618 4324 22670
rect 4348 22618 4358 22670
rect 4358 22618 4404 22670
rect 4428 22618 4474 22670
rect 4474 22618 4484 22670
rect 4508 22618 4538 22670
rect 4538 22618 4564 22670
rect 4268 22616 4324 22618
rect 4348 22616 4404 22618
rect 4428 22616 4484 22618
rect 4508 22616 4564 22618
rect 4268 21338 4324 21340
rect 4348 21338 4404 21340
rect 4428 21338 4484 21340
rect 4508 21338 4564 21340
rect 4268 21286 4294 21338
rect 4294 21286 4324 21338
rect 4348 21286 4358 21338
rect 4358 21286 4404 21338
rect 4428 21286 4474 21338
rect 4474 21286 4484 21338
rect 4508 21286 4538 21338
rect 4538 21286 4564 21338
rect 4268 21284 4324 21286
rect 4348 21284 4404 21286
rect 4428 21284 4484 21286
rect 4508 21284 4564 21286
rect 4268 20006 4324 20008
rect 4348 20006 4404 20008
rect 4428 20006 4484 20008
rect 4508 20006 4564 20008
rect 4268 19954 4294 20006
rect 4294 19954 4324 20006
rect 4348 19954 4358 20006
rect 4358 19954 4404 20006
rect 4428 19954 4474 20006
rect 4474 19954 4484 20006
rect 4508 19954 4538 20006
rect 4538 19954 4564 20006
rect 4268 19952 4324 19954
rect 4348 19952 4404 19954
rect 4428 19952 4484 19954
rect 4508 19952 4564 19954
rect 4268 18674 4324 18676
rect 4348 18674 4404 18676
rect 4428 18674 4484 18676
rect 4508 18674 4564 18676
rect 4268 18622 4294 18674
rect 4294 18622 4324 18674
rect 4348 18622 4358 18674
rect 4358 18622 4404 18674
rect 4428 18622 4474 18674
rect 4474 18622 4484 18674
rect 4508 18622 4538 18674
rect 4538 18622 4564 18674
rect 4268 18620 4324 18622
rect 4348 18620 4404 18622
rect 4428 18620 4484 18622
rect 4508 18620 4564 18622
rect 4268 17342 4324 17344
rect 4348 17342 4404 17344
rect 4428 17342 4484 17344
rect 4508 17342 4564 17344
rect 4268 17290 4294 17342
rect 4294 17290 4324 17342
rect 4348 17290 4358 17342
rect 4358 17290 4404 17342
rect 4428 17290 4474 17342
rect 4474 17290 4484 17342
rect 4508 17290 4538 17342
rect 4538 17290 4564 17342
rect 4268 17288 4324 17290
rect 4348 17288 4404 17290
rect 4428 17288 4484 17290
rect 4508 17288 4564 17290
rect 4268 16010 4324 16012
rect 4348 16010 4404 16012
rect 4428 16010 4484 16012
rect 4508 16010 4564 16012
rect 4268 15958 4294 16010
rect 4294 15958 4324 16010
rect 4348 15958 4358 16010
rect 4358 15958 4404 16010
rect 4428 15958 4474 16010
rect 4474 15958 4484 16010
rect 4508 15958 4538 16010
rect 4538 15958 4564 16010
rect 4268 15956 4324 15958
rect 4348 15956 4404 15958
rect 4428 15956 4484 15958
rect 4508 15956 4564 15958
rect 4268 14678 4324 14680
rect 4348 14678 4404 14680
rect 4428 14678 4484 14680
rect 4508 14678 4564 14680
rect 4268 14626 4294 14678
rect 4294 14626 4324 14678
rect 4348 14626 4358 14678
rect 4358 14626 4404 14678
rect 4428 14626 4474 14678
rect 4474 14626 4484 14678
rect 4508 14626 4538 14678
rect 4538 14626 4564 14678
rect 4268 14624 4324 14626
rect 4348 14624 4404 14626
rect 4428 14624 4484 14626
rect 4508 14624 4564 14626
rect 4268 13346 4324 13348
rect 4348 13346 4404 13348
rect 4428 13346 4484 13348
rect 4508 13346 4564 13348
rect 4268 13294 4294 13346
rect 4294 13294 4324 13346
rect 4348 13294 4358 13346
rect 4358 13294 4404 13346
rect 4428 13294 4474 13346
rect 4474 13294 4484 13346
rect 4508 13294 4538 13346
rect 4538 13294 4564 13346
rect 4268 13292 4324 13294
rect 4348 13292 4404 13294
rect 4428 13292 4484 13294
rect 4508 13292 4564 13294
rect 4268 12014 4324 12016
rect 4348 12014 4404 12016
rect 4428 12014 4484 12016
rect 4508 12014 4564 12016
rect 4268 11962 4294 12014
rect 4294 11962 4324 12014
rect 4348 11962 4358 12014
rect 4358 11962 4404 12014
rect 4428 11962 4474 12014
rect 4474 11962 4484 12014
rect 4508 11962 4538 12014
rect 4538 11962 4564 12014
rect 4268 11960 4324 11962
rect 4348 11960 4404 11962
rect 4428 11960 4484 11962
rect 4508 11960 4564 11962
rect 4268 10682 4324 10684
rect 4348 10682 4404 10684
rect 4428 10682 4484 10684
rect 4508 10682 4564 10684
rect 4268 10630 4294 10682
rect 4294 10630 4324 10682
rect 4348 10630 4358 10682
rect 4358 10630 4404 10682
rect 4428 10630 4474 10682
rect 4474 10630 4484 10682
rect 4508 10630 4538 10682
rect 4538 10630 4564 10682
rect 4268 10628 4324 10630
rect 4348 10628 4404 10630
rect 4428 10628 4484 10630
rect 4508 10628 4564 10630
rect 4268 9350 4324 9352
rect 4348 9350 4404 9352
rect 4428 9350 4484 9352
rect 4508 9350 4564 9352
rect 4268 9298 4294 9350
rect 4294 9298 4324 9350
rect 4348 9298 4358 9350
rect 4358 9298 4404 9350
rect 4428 9298 4474 9350
rect 4474 9298 4484 9350
rect 4508 9298 4538 9350
rect 4538 9298 4564 9350
rect 4268 9296 4324 9298
rect 4348 9296 4404 9298
rect 4428 9296 4484 9298
rect 4508 9296 4564 9298
rect 4268 8018 4324 8020
rect 4348 8018 4404 8020
rect 4428 8018 4484 8020
rect 4508 8018 4564 8020
rect 4268 7966 4294 8018
rect 4294 7966 4324 8018
rect 4348 7966 4358 8018
rect 4358 7966 4404 8018
rect 4428 7966 4474 8018
rect 4474 7966 4484 8018
rect 4508 7966 4538 8018
rect 4538 7966 4564 8018
rect 4268 7964 4324 7966
rect 4348 7964 4404 7966
rect 4428 7964 4484 7966
rect 4508 7964 4564 7966
rect 4532 6893 4534 6910
rect 4534 6893 4586 6910
rect 4586 6893 4588 6910
rect 4532 6854 4588 6893
rect 4268 6686 4324 6688
rect 4348 6686 4404 6688
rect 4428 6686 4484 6688
rect 4508 6686 4564 6688
rect 4268 6634 4294 6686
rect 4294 6634 4324 6686
rect 4348 6634 4358 6686
rect 4358 6634 4404 6686
rect 4428 6634 4474 6686
rect 4474 6634 4484 6686
rect 4508 6634 4538 6686
rect 4538 6634 4564 6686
rect 4268 6632 4324 6634
rect 4348 6632 4404 6634
rect 4428 6632 4484 6634
rect 4508 6632 4564 6634
rect 4268 5354 4324 5356
rect 4348 5354 4404 5356
rect 4428 5354 4484 5356
rect 4508 5354 4564 5356
rect 4268 5302 4294 5354
rect 4294 5302 4324 5354
rect 4348 5302 4358 5354
rect 4358 5302 4404 5354
rect 4428 5302 4474 5354
rect 4474 5302 4484 5354
rect 4508 5302 4538 5354
rect 4538 5302 4564 5354
rect 4268 5300 4324 5302
rect 4348 5300 4404 5302
rect 4428 5300 4484 5302
rect 4508 5300 4564 5302
rect 4268 4022 4324 4024
rect 4348 4022 4404 4024
rect 4428 4022 4484 4024
rect 4508 4022 4564 4024
rect 4268 3970 4294 4022
rect 4294 3970 4324 4022
rect 4348 3970 4358 4022
rect 4358 3970 4404 4022
rect 4428 3970 4474 4022
rect 4474 3970 4484 4022
rect 4508 3970 4538 4022
rect 4538 3970 4564 4022
rect 4268 3968 4324 3970
rect 4348 3968 4404 3970
rect 4428 3968 4484 3970
rect 4508 3968 4564 3970
rect 4268 2690 4324 2692
rect 4348 2690 4404 2692
rect 4428 2690 4484 2692
rect 4508 2690 4564 2692
rect 4268 2638 4294 2690
rect 4294 2638 4324 2690
rect 4348 2638 4358 2690
rect 4358 2638 4404 2690
rect 4428 2638 4474 2690
rect 4474 2638 4484 2690
rect 4508 2638 4538 2690
rect 4538 2638 4564 2690
rect 4268 2636 4324 2638
rect 4348 2636 4404 2638
rect 4428 2636 4484 2638
rect 4508 2636 4564 2638
rect 7220 56177 7222 56194
rect 7222 56177 7274 56194
rect 7274 56177 7276 56194
rect 7220 56138 7276 56177
rect 5396 7041 5398 7058
rect 5398 7041 5450 7058
rect 5450 7041 5452 7058
rect 5396 7002 5452 7041
rect 6740 7298 6796 7354
rect 8372 28906 8428 28962
rect 7220 24910 7276 24966
rect 8372 26094 8428 26150
rect 8228 24927 8284 24966
rect 8228 24910 8230 24927
rect 8230 24910 8282 24927
rect 8282 24910 8284 24927
rect 7412 17231 7468 17270
rect 7412 17214 7414 17231
rect 7414 17214 7466 17231
rect 7466 17214 7468 17231
rect 7316 7150 7372 7206
rect 7508 8482 7564 8538
rect 7796 13366 7852 13422
rect 7988 13366 8044 13422
rect 7604 7742 7660 7798
rect 7892 8482 7948 8538
rect 7988 8334 8044 8390
rect 7892 7150 7948 7206
rect 8084 4338 8140 4394
rect 7988 4190 8044 4246
rect 8372 9666 8428 9722
rect 8660 9074 8716 9130
rect 8564 8926 8620 8982
rect 8756 8926 8812 8982
rect 8564 8225 8566 8242
rect 8566 8225 8618 8242
rect 8618 8225 8620 8242
rect 8564 8186 8620 8225
rect 8564 7890 8620 7946
rect 8468 7446 8524 7502
rect 8756 7742 8812 7798
rect 8756 7485 8758 7502
rect 8758 7485 8810 7502
rect 8810 7485 8812 7502
rect 8756 7446 8812 7485
rect 9044 17231 9100 17270
rect 9044 17214 9046 17231
rect 9046 17214 9098 17231
rect 9098 17214 9100 17231
rect 9044 8965 9046 8982
rect 9046 8965 9098 8982
rect 9098 8965 9100 8982
rect 9044 8926 9100 8965
rect 9044 7890 9100 7946
rect 8564 3746 8620 3802
rect 9428 7890 9484 7946
rect 10196 7759 10252 7798
rect 10196 7742 10198 7759
rect 10198 7742 10250 7759
rect 10250 7742 10252 7759
rect 9908 7485 9910 7502
rect 9910 7485 9962 7502
rect 9962 7485 9964 7502
rect 9908 7446 9964 7485
rect 10004 6871 10060 6910
rect 10004 6854 10006 6871
rect 10006 6854 10058 6871
rect 10058 6854 10060 6871
rect 9716 4486 9772 4542
rect 9908 3894 9964 3950
rect 10580 6893 10582 6910
rect 10582 6893 10634 6910
rect 10634 6893 10636 6910
rect 10580 6854 10636 6893
rect 10868 8778 10924 8834
rect 10868 6706 10924 6762
rect 11060 8630 11116 8686
rect 12212 7150 12268 7206
rect 12404 8334 12460 8390
rect 12980 8482 13036 8538
rect 13652 8482 13708 8538
rect 12788 7298 12844 7354
rect 13940 7446 13996 7502
rect 13268 7298 13324 7354
rect 12980 6706 13036 6762
rect 13748 3746 13804 3802
rect 16436 8778 16492 8834
rect 16340 8630 16396 8686
rect 17588 6114 17644 6170
rect 17780 5818 17836 5874
rect 18356 6558 18412 6614
rect 18932 7298 18988 7354
rect 19628 56636 19684 56638
rect 19708 56636 19764 56638
rect 19788 56636 19844 56638
rect 19868 56636 19924 56638
rect 19628 56584 19654 56636
rect 19654 56584 19684 56636
rect 19708 56584 19718 56636
rect 19718 56584 19764 56636
rect 19788 56584 19834 56636
rect 19834 56584 19844 56636
rect 19868 56584 19898 56636
rect 19898 56584 19924 56636
rect 19628 56582 19684 56584
rect 19708 56582 19764 56584
rect 19788 56582 19844 56584
rect 19868 56582 19924 56584
rect 19628 55304 19684 55306
rect 19708 55304 19764 55306
rect 19788 55304 19844 55306
rect 19868 55304 19924 55306
rect 19628 55252 19654 55304
rect 19654 55252 19684 55304
rect 19708 55252 19718 55304
rect 19718 55252 19764 55304
rect 19788 55252 19834 55304
rect 19834 55252 19844 55304
rect 19868 55252 19898 55304
rect 19898 55252 19924 55304
rect 19628 55250 19684 55252
rect 19708 55250 19764 55252
rect 19788 55250 19844 55252
rect 19868 55250 19924 55252
rect 19628 53972 19684 53974
rect 19708 53972 19764 53974
rect 19788 53972 19844 53974
rect 19868 53972 19924 53974
rect 19628 53920 19654 53972
rect 19654 53920 19684 53972
rect 19708 53920 19718 53972
rect 19718 53920 19764 53972
rect 19788 53920 19834 53972
rect 19834 53920 19844 53972
rect 19868 53920 19898 53972
rect 19898 53920 19924 53972
rect 19628 53918 19684 53920
rect 19708 53918 19764 53920
rect 19788 53918 19844 53920
rect 19868 53918 19924 53920
rect 19628 52640 19684 52642
rect 19708 52640 19764 52642
rect 19788 52640 19844 52642
rect 19868 52640 19924 52642
rect 19628 52588 19654 52640
rect 19654 52588 19684 52640
rect 19708 52588 19718 52640
rect 19718 52588 19764 52640
rect 19788 52588 19834 52640
rect 19834 52588 19844 52640
rect 19868 52588 19898 52640
rect 19898 52588 19924 52640
rect 19628 52586 19684 52588
rect 19708 52586 19764 52588
rect 19788 52586 19844 52588
rect 19868 52586 19924 52588
rect 19628 51308 19684 51310
rect 19708 51308 19764 51310
rect 19788 51308 19844 51310
rect 19868 51308 19924 51310
rect 19628 51256 19654 51308
rect 19654 51256 19684 51308
rect 19708 51256 19718 51308
rect 19718 51256 19764 51308
rect 19788 51256 19834 51308
rect 19834 51256 19844 51308
rect 19868 51256 19898 51308
rect 19898 51256 19924 51308
rect 19628 51254 19684 51256
rect 19708 51254 19764 51256
rect 19788 51254 19844 51256
rect 19868 51254 19924 51256
rect 19628 49976 19684 49978
rect 19708 49976 19764 49978
rect 19788 49976 19844 49978
rect 19868 49976 19924 49978
rect 19628 49924 19654 49976
rect 19654 49924 19684 49976
rect 19708 49924 19718 49976
rect 19718 49924 19764 49976
rect 19788 49924 19834 49976
rect 19834 49924 19844 49976
rect 19868 49924 19898 49976
rect 19898 49924 19924 49976
rect 19628 49922 19684 49924
rect 19708 49922 19764 49924
rect 19788 49922 19844 49924
rect 19868 49922 19924 49924
rect 19628 48644 19684 48646
rect 19708 48644 19764 48646
rect 19788 48644 19844 48646
rect 19868 48644 19924 48646
rect 19628 48592 19654 48644
rect 19654 48592 19684 48644
rect 19708 48592 19718 48644
rect 19718 48592 19764 48644
rect 19788 48592 19834 48644
rect 19834 48592 19844 48644
rect 19868 48592 19898 48644
rect 19898 48592 19924 48644
rect 19628 48590 19684 48592
rect 19708 48590 19764 48592
rect 19788 48590 19844 48592
rect 19868 48590 19924 48592
rect 19628 47312 19684 47314
rect 19708 47312 19764 47314
rect 19788 47312 19844 47314
rect 19868 47312 19924 47314
rect 19628 47260 19654 47312
rect 19654 47260 19684 47312
rect 19708 47260 19718 47312
rect 19718 47260 19764 47312
rect 19788 47260 19834 47312
rect 19834 47260 19844 47312
rect 19868 47260 19898 47312
rect 19898 47260 19924 47312
rect 19628 47258 19684 47260
rect 19708 47258 19764 47260
rect 19788 47258 19844 47260
rect 19868 47258 19924 47260
rect 19628 45980 19684 45982
rect 19708 45980 19764 45982
rect 19788 45980 19844 45982
rect 19868 45980 19924 45982
rect 19628 45928 19654 45980
rect 19654 45928 19684 45980
rect 19708 45928 19718 45980
rect 19718 45928 19764 45980
rect 19788 45928 19834 45980
rect 19834 45928 19844 45980
rect 19868 45928 19898 45980
rect 19898 45928 19924 45980
rect 19628 45926 19684 45928
rect 19708 45926 19764 45928
rect 19788 45926 19844 45928
rect 19868 45926 19924 45928
rect 19628 44648 19684 44650
rect 19708 44648 19764 44650
rect 19788 44648 19844 44650
rect 19868 44648 19924 44650
rect 19628 44596 19654 44648
rect 19654 44596 19684 44648
rect 19708 44596 19718 44648
rect 19718 44596 19764 44648
rect 19788 44596 19834 44648
rect 19834 44596 19844 44648
rect 19868 44596 19898 44648
rect 19898 44596 19924 44648
rect 19628 44594 19684 44596
rect 19708 44594 19764 44596
rect 19788 44594 19844 44596
rect 19868 44594 19924 44596
rect 19628 43316 19684 43318
rect 19708 43316 19764 43318
rect 19788 43316 19844 43318
rect 19868 43316 19924 43318
rect 19628 43264 19654 43316
rect 19654 43264 19684 43316
rect 19708 43264 19718 43316
rect 19718 43264 19764 43316
rect 19788 43264 19834 43316
rect 19834 43264 19844 43316
rect 19868 43264 19898 43316
rect 19898 43264 19924 43316
rect 19628 43262 19684 43264
rect 19708 43262 19764 43264
rect 19788 43262 19844 43264
rect 19868 43262 19924 43264
rect 19628 41984 19684 41986
rect 19708 41984 19764 41986
rect 19788 41984 19844 41986
rect 19868 41984 19924 41986
rect 19628 41932 19654 41984
rect 19654 41932 19684 41984
rect 19708 41932 19718 41984
rect 19718 41932 19764 41984
rect 19788 41932 19834 41984
rect 19834 41932 19844 41984
rect 19868 41932 19898 41984
rect 19898 41932 19924 41984
rect 19628 41930 19684 41932
rect 19708 41930 19764 41932
rect 19788 41930 19844 41932
rect 19868 41930 19924 41932
rect 19628 40652 19684 40654
rect 19708 40652 19764 40654
rect 19788 40652 19844 40654
rect 19868 40652 19924 40654
rect 19628 40600 19654 40652
rect 19654 40600 19684 40652
rect 19708 40600 19718 40652
rect 19718 40600 19764 40652
rect 19788 40600 19834 40652
rect 19834 40600 19844 40652
rect 19868 40600 19898 40652
rect 19898 40600 19924 40652
rect 19628 40598 19684 40600
rect 19708 40598 19764 40600
rect 19788 40598 19844 40600
rect 19868 40598 19924 40600
rect 19628 39320 19684 39322
rect 19708 39320 19764 39322
rect 19788 39320 19844 39322
rect 19868 39320 19924 39322
rect 19628 39268 19654 39320
rect 19654 39268 19684 39320
rect 19708 39268 19718 39320
rect 19718 39268 19764 39320
rect 19788 39268 19834 39320
rect 19834 39268 19844 39320
rect 19868 39268 19898 39320
rect 19898 39268 19924 39320
rect 19628 39266 19684 39268
rect 19708 39266 19764 39268
rect 19788 39266 19844 39268
rect 19868 39266 19924 39268
rect 19628 37988 19684 37990
rect 19708 37988 19764 37990
rect 19788 37988 19844 37990
rect 19868 37988 19924 37990
rect 19628 37936 19654 37988
rect 19654 37936 19684 37988
rect 19708 37936 19718 37988
rect 19718 37936 19764 37988
rect 19788 37936 19834 37988
rect 19834 37936 19844 37988
rect 19868 37936 19898 37988
rect 19898 37936 19924 37988
rect 19628 37934 19684 37936
rect 19708 37934 19764 37936
rect 19788 37934 19844 37936
rect 19868 37934 19924 37936
rect 19628 36656 19684 36658
rect 19708 36656 19764 36658
rect 19788 36656 19844 36658
rect 19868 36656 19924 36658
rect 19628 36604 19654 36656
rect 19654 36604 19684 36656
rect 19708 36604 19718 36656
rect 19718 36604 19764 36656
rect 19788 36604 19834 36656
rect 19834 36604 19844 36656
rect 19868 36604 19898 36656
rect 19898 36604 19924 36656
rect 19628 36602 19684 36604
rect 19708 36602 19764 36604
rect 19788 36602 19844 36604
rect 19868 36602 19924 36604
rect 19628 35324 19684 35326
rect 19708 35324 19764 35326
rect 19788 35324 19844 35326
rect 19868 35324 19924 35326
rect 19628 35272 19654 35324
rect 19654 35272 19684 35324
rect 19708 35272 19718 35324
rect 19718 35272 19764 35324
rect 19788 35272 19834 35324
rect 19834 35272 19844 35324
rect 19868 35272 19898 35324
rect 19898 35272 19924 35324
rect 19628 35270 19684 35272
rect 19708 35270 19764 35272
rect 19788 35270 19844 35272
rect 19868 35270 19924 35272
rect 19628 33992 19684 33994
rect 19708 33992 19764 33994
rect 19788 33992 19844 33994
rect 19868 33992 19924 33994
rect 19628 33940 19654 33992
rect 19654 33940 19684 33992
rect 19708 33940 19718 33992
rect 19718 33940 19764 33992
rect 19788 33940 19834 33992
rect 19834 33940 19844 33992
rect 19868 33940 19898 33992
rect 19898 33940 19924 33992
rect 19628 33938 19684 33940
rect 19708 33938 19764 33940
rect 19788 33938 19844 33940
rect 19868 33938 19924 33940
rect 19628 32660 19684 32662
rect 19708 32660 19764 32662
rect 19788 32660 19844 32662
rect 19868 32660 19924 32662
rect 19628 32608 19654 32660
rect 19654 32608 19684 32660
rect 19708 32608 19718 32660
rect 19718 32608 19764 32660
rect 19788 32608 19834 32660
rect 19834 32608 19844 32660
rect 19868 32608 19898 32660
rect 19898 32608 19924 32660
rect 19628 32606 19684 32608
rect 19708 32606 19764 32608
rect 19788 32606 19844 32608
rect 19868 32606 19924 32608
rect 19628 31328 19684 31330
rect 19708 31328 19764 31330
rect 19788 31328 19844 31330
rect 19868 31328 19924 31330
rect 19628 31276 19654 31328
rect 19654 31276 19684 31328
rect 19708 31276 19718 31328
rect 19718 31276 19764 31328
rect 19788 31276 19834 31328
rect 19834 31276 19844 31328
rect 19868 31276 19898 31328
rect 19898 31276 19924 31328
rect 19628 31274 19684 31276
rect 19708 31274 19764 31276
rect 19788 31274 19844 31276
rect 19868 31274 19924 31276
rect 19628 29996 19684 29998
rect 19708 29996 19764 29998
rect 19788 29996 19844 29998
rect 19868 29996 19924 29998
rect 19628 29944 19654 29996
rect 19654 29944 19684 29996
rect 19708 29944 19718 29996
rect 19718 29944 19764 29996
rect 19788 29944 19834 29996
rect 19834 29944 19844 29996
rect 19868 29944 19898 29996
rect 19898 29944 19924 29996
rect 19628 29942 19684 29944
rect 19708 29942 19764 29944
rect 19788 29942 19844 29944
rect 19868 29942 19924 29944
rect 19628 28664 19684 28666
rect 19708 28664 19764 28666
rect 19788 28664 19844 28666
rect 19868 28664 19924 28666
rect 19628 28612 19654 28664
rect 19654 28612 19684 28664
rect 19708 28612 19718 28664
rect 19718 28612 19764 28664
rect 19788 28612 19834 28664
rect 19834 28612 19844 28664
rect 19868 28612 19898 28664
rect 19898 28612 19924 28664
rect 19628 28610 19684 28612
rect 19708 28610 19764 28612
rect 19788 28610 19844 28612
rect 19868 28610 19924 28612
rect 19628 27332 19684 27334
rect 19708 27332 19764 27334
rect 19788 27332 19844 27334
rect 19868 27332 19924 27334
rect 19628 27280 19654 27332
rect 19654 27280 19684 27332
rect 19708 27280 19718 27332
rect 19718 27280 19764 27332
rect 19788 27280 19834 27332
rect 19834 27280 19844 27332
rect 19868 27280 19898 27332
rect 19898 27280 19924 27332
rect 19628 27278 19684 27280
rect 19708 27278 19764 27280
rect 19788 27278 19844 27280
rect 19868 27278 19924 27280
rect 19628 26000 19684 26002
rect 19708 26000 19764 26002
rect 19788 26000 19844 26002
rect 19868 26000 19924 26002
rect 19628 25948 19654 26000
rect 19654 25948 19684 26000
rect 19708 25948 19718 26000
rect 19718 25948 19764 26000
rect 19788 25948 19834 26000
rect 19834 25948 19844 26000
rect 19868 25948 19898 26000
rect 19898 25948 19924 26000
rect 19628 25946 19684 25948
rect 19708 25946 19764 25948
rect 19788 25946 19844 25948
rect 19868 25946 19924 25948
rect 19628 24668 19684 24670
rect 19708 24668 19764 24670
rect 19788 24668 19844 24670
rect 19868 24668 19924 24670
rect 19628 24616 19654 24668
rect 19654 24616 19684 24668
rect 19708 24616 19718 24668
rect 19718 24616 19764 24668
rect 19788 24616 19834 24668
rect 19834 24616 19844 24668
rect 19868 24616 19898 24668
rect 19898 24616 19924 24668
rect 19628 24614 19684 24616
rect 19708 24614 19764 24616
rect 19788 24614 19844 24616
rect 19868 24614 19924 24616
rect 19628 23336 19684 23338
rect 19708 23336 19764 23338
rect 19788 23336 19844 23338
rect 19868 23336 19924 23338
rect 19628 23284 19654 23336
rect 19654 23284 19684 23336
rect 19708 23284 19718 23336
rect 19718 23284 19764 23336
rect 19788 23284 19834 23336
rect 19834 23284 19844 23336
rect 19868 23284 19898 23336
rect 19898 23284 19924 23336
rect 19628 23282 19684 23284
rect 19708 23282 19764 23284
rect 19788 23282 19844 23284
rect 19868 23282 19924 23284
rect 19628 22004 19684 22006
rect 19708 22004 19764 22006
rect 19788 22004 19844 22006
rect 19868 22004 19924 22006
rect 19628 21952 19654 22004
rect 19654 21952 19684 22004
rect 19708 21952 19718 22004
rect 19718 21952 19764 22004
rect 19788 21952 19834 22004
rect 19834 21952 19844 22004
rect 19868 21952 19898 22004
rect 19898 21952 19924 22004
rect 19628 21950 19684 21952
rect 19708 21950 19764 21952
rect 19788 21950 19844 21952
rect 19868 21950 19924 21952
rect 19628 20672 19684 20674
rect 19708 20672 19764 20674
rect 19788 20672 19844 20674
rect 19868 20672 19924 20674
rect 19628 20620 19654 20672
rect 19654 20620 19684 20672
rect 19708 20620 19718 20672
rect 19718 20620 19764 20672
rect 19788 20620 19834 20672
rect 19834 20620 19844 20672
rect 19868 20620 19898 20672
rect 19898 20620 19924 20672
rect 19628 20618 19684 20620
rect 19708 20618 19764 20620
rect 19788 20618 19844 20620
rect 19868 20618 19924 20620
rect 19628 19340 19684 19342
rect 19708 19340 19764 19342
rect 19788 19340 19844 19342
rect 19868 19340 19924 19342
rect 19628 19288 19654 19340
rect 19654 19288 19684 19340
rect 19708 19288 19718 19340
rect 19718 19288 19764 19340
rect 19788 19288 19834 19340
rect 19834 19288 19844 19340
rect 19868 19288 19898 19340
rect 19898 19288 19924 19340
rect 19628 19286 19684 19288
rect 19708 19286 19764 19288
rect 19788 19286 19844 19288
rect 19868 19286 19924 19288
rect 19628 18008 19684 18010
rect 19708 18008 19764 18010
rect 19788 18008 19844 18010
rect 19868 18008 19924 18010
rect 19628 17956 19654 18008
rect 19654 17956 19684 18008
rect 19708 17956 19718 18008
rect 19718 17956 19764 18008
rect 19788 17956 19834 18008
rect 19834 17956 19844 18008
rect 19868 17956 19898 18008
rect 19898 17956 19924 18008
rect 19628 17954 19684 17956
rect 19708 17954 19764 17956
rect 19788 17954 19844 17956
rect 19868 17954 19924 17956
rect 19628 16676 19684 16678
rect 19708 16676 19764 16678
rect 19788 16676 19844 16678
rect 19868 16676 19924 16678
rect 19628 16624 19654 16676
rect 19654 16624 19684 16676
rect 19708 16624 19718 16676
rect 19718 16624 19764 16676
rect 19788 16624 19834 16676
rect 19834 16624 19844 16676
rect 19868 16624 19898 16676
rect 19898 16624 19924 16676
rect 19628 16622 19684 16624
rect 19708 16622 19764 16624
rect 19788 16622 19844 16624
rect 19868 16622 19924 16624
rect 19628 15344 19684 15346
rect 19708 15344 19764 15346
rect 19788 15344 19844 15346
rect 19868 15344 19924 15346
rect 19628 15292 19654 15344
rect 19654 15292 19684 15344
rect 19708 15292 19718 15344
rect 19718 15292 19764 15344
rect 19788 15292 19834 15344
rect 19834 15292 19844 15344
rect 19868 15292 19898 15344
rect 19898 15292 19924 15344
rect 19628 15290 19684 15292
rect 19708 15290 19764 15292
rect 19788 15290 19844 15292
rect 19868 15290 19924 15292
rect 19628 14012 19684 14014
rect 19708 14012 19764 14014
rect 19788 14012 19844 14014
rect 19868 14012 19924 14014
rect 19628 13960 19654 14012
rect 19654 13960 19684 14012
rect 19708 13960 19718 14012
rect 19718 13960 19764 14012
rect 19788 13960 19834 14012
rect 19834 13960 19844 14012
rect 19868 13960 19898 14012
rect 19898 13960 19924 14012
rect 19628 13958 19684 13960
rect 19708 13958 19764 13960
rect 19788 13958 19844 13960
rect 19868 13958 19924 13960
rect 19628 12680 19684 12682
rect 19708 12680 19764 12682
rect 19788 12680 19844 12682
rect 19868 12680 19924 12682
rect 19628 12628 19654 12680
rect 19654 12628 19684 12680
rect 19708 12628 19718 12680
rect 19718 12628 19764 12680
rect 19788 12628 19834 12680
rect 19834 12628 19844 12680
rect 19868 12628 19898 12680
rect 19898 12628 19924 12680
rect 19628 12626 19684 12628
rect 19708 12626 19764 12628
rect 19788 12626 19844 12628
rect 19868 12626 19924 12628
rect 19628 11348 19684 11350
rect 19708 11348 19764 11350
rect 19788 11348 19844 11350
rect 19868 11348 19924 11350
rect 19628 11296 19654 11348
rect 19654 11296 19684 11348
rect 19708 11296 19718 11348
rect 19718 11296 19764 11348
rect 19788 11296 19834 11348
rect 19834 11296 19844 11348
rect 19868 11296 19898 11348
rect 19898 11296 19924 11348
rect 19628 11294 19684 11296
rect 19708 11294 19764 11296
rect 19788 11294 19844 11296
rect 19868 11294 19924 11296
rect 19628 10016 19684 10018
rect 19708 10016 19764 10018
rect 19788 10016 19844 10018
rect 19868 10016 19924 10018
rect 19628 9964 19654 10016
rect 19654 9964 19684 10016
rect 19708 9964 19718 10016
rect 19718 9964 19764 10016
rect 19788 9964 19834 10016
rect 19834 9964 19844 10016
rect 19868 9964 19898 10016
rect 19898 9964 19924 10016
rect 19628 9962 19684 9964
rect 19708 9962 19764 9964
rect 19788 9962 19844 9964
rect 19868 9962 19924 9964
rect 19628 8684 19684 8686
rect 19708 8684 19764 8686
rect 19788 8684 19844 8686
rect 19868 8684 19924 8686
rect 19628 8632 19654 8684
rect 19654 8632 19684 8684
rect 19708 8632 19718 8684
rect 19718 8632 19764 8684
rect 19788 8632 19834 8684
rect 19834 8632 19844 8684
rect 19868 8632 19898 8684
rect 19898 8632 19924 8684
rect 19628 8630 19684 8632
rect 19708 8630 19764 8632
rect 19788 8630 19844 8632
rect 19868 8630 19924 8632
rect 19628 7352 19684 7354
rect 19708 7352 19764 7354
rect 19788 7352 19844 7354
rect 19868 7352 19924 7354
rect 19628 7300 19654 7352
rect 19654 7300 19684 7352
rect 19708 7300 19718 7352
rect 19718 7300 19764 7352
rect 19788 7300 19834 7352
rect 19834 7300 19844 7352
rect 19868 7300 19898 7352
rect 19898 7300 19924 7352
rect 19628 7298 19684 7300
rect 19708 7298 19764 7300
rect 19788 7298 19844 7300
rect 19868 7298 19924 7300
rect 19604 6427 19660 6466
rect 20468 7298 20524 7354
rect 19604 6410 19606 6427
rect 19606 6410 19658 6427
rect 19658 6410 19660 6427
rect 19220 4190 19276 4246
rect 19628 6020 19684 6022
rect 19708 6020 19764 6022
rect 19788 6020 19844 6022
rect 19868 6020 19924 6022
rect 19628 5968 19654 6020
rect 19654 5968 19684 6020
rect 19708 5968 19718 6020
rect 19718 5968 19764 6020
rect 19788 5968 19834 6020
rect 19834 5968 19844 6020
rect 19868 5968 19898 6020
rect 19898 5968 19924 6020
rect 19628 5966 19684 5968
rect 19708 5966 19764 5968
rect 19788 5966 19844 5968
rect 19868 5966 19924 5968
rect 19628 4688 19684 4690
rect 19708 4688 19764 4690
rect 19788 4688 19844 4690
rect 19868 4688 19924 4690
rect 19628 4636 19654 4688
rect 19654 4636 19684 4688
rect 19708 4636 19718 4688
rect 19718 4636 19764 4688
rect 19788 4636 19834 4688
rect 19834 4636 19844 4688
rect 19868 4636 19898 4688
rect 19898 4636 19924 4688
rect 19628 4634 19684 4636
rect 19708 4634 19764 4636
rect 19788 4634 19844 4636
rect 19868 4634 19924 4636
rect 19628 3356 19684 3358
rect 19708 3356 19764 3358
rect 19788 3356 19844 3358
rect 19868 3356 19924 3358
rect 19628 3304 19654 3356
rect 19654 3304 19684 3356
rect 19708 3304 19718 3356
rect 19718 3304 19764 3356
rect 19788 3304 19834 3356
rect 19834 3304 19844 3356
rect 19868 3304 19898 3356
rect 19898 3304 19924 3356
rect 19628 3302 19684 3304
rect 19708 3302 19764 3304
rect 19788 3302 19844 3304
rect 19868 3302 19924 3304
rect 21332 5966 21388 6022
rect 20852 3467 20908 3506
rect 20852 3450 20854 3467
rect 20854 3450 20906 3467
rect 20906 3450 20908 3467
rect 21140 3171 21196 3210
rect 21140 3154 21142 3171
rect 21142 3154 21194 3171
rect 21194 3154 21196 3171
rect 21140 2897 21142 2914
rect 21142 2897 21194 2914
rect 21194 2897 21196 2914
rect 21140 2858 21196 2897
rect 22676 6410 22732 6466
rect 22676 5670 22732 5726
rect 23156 7298 23212 7354
rect 23636 6558 23692 6614
rect 23828 7298 23884 7354
rect 24020 6262 24076 6318
rect 28052 7890 28108 7946
rect 27284 7298 27340 7354
rect 28052 7298 28108 7354
rect 28436 6558 28492 6614
rect 30836 8038 30892 8094
rect 30068 5670 30124 5726
rect 34988 57302 35044 57304
rect 35068 57302 35124 57304
rect 35148 57302 35204 57304
rect 35228 57302 35284 57304
rect 34988 57250 35014 57302
rect 35014 57250 35044 57302
rect 35068 57250 35078 57302
rect 35078 57250 35124 57302
rect 35148 57250 35194 57302
rect 35194 57250 35204 57302
rect 35228 57250 35258 57302
rect 35258 57250 35284 57302
rect 34988 57248 35044 57250
rect 35068 57248 35124 57250
rect 35148 57248 35204 57250
rect 35228 57248 35284 57250
rect 32852 6558 32908 6614
rect 32756 6262 32812 6318
rect 33044 6706 33100 6762
rect 33140 6558 33196 6614
rect 34988 55970 35044 55972
rect 35068 55970 35124 55972
rect 35148 55970 35204 55972
rect 35228 55970 35284 55972
rect 34988 55918 35014 55970
rect 35014 55918 35044 55970
rect 35068 55918 35078 55970
rect 35078 55918 35124 55970
rect 35148 55918 35194 55970
rect 35194 55918 35204 55970
rect 35228 55918 35258 55970
rect 35258 55918 35284 55970
rect 34988 55916 35044 55918
rect 35068 55916 35124 55918
rect 35148 55916 35204 55918
rect 35228 55916 35284 55918
rect 34988 54638 35044 54640
rect 35068 54638 35124 54640
rect 35148 54638 35204 54640
rect 35228 54638 35284 54640
rect 34988 54586 35014 54638
rect 35014 54586 35044 54638
rect 35068 54586 35078 54638
rect 35078 54586 35124 54638
rect 35148 54586 35194 54638
rect 35194 54586 35204 54638
rect 35228 54586 35258 54638
rect 35258 54586 35284 54638
rect 34988 54584 35044 54586
rect 35068 54584 35124 54586
rect 35148 54584 35204 54586
rect 35228 54584 35284 54586
rect 34988 53306 35044 53308
rect 35068 53306 35124 53308
rect 35148 53306 35204 53308
rect 35228 53306 35284 53308
rect 34988 53254 35014 53306
rect 35014 53254 35044 53306
rect 35068 53254 35078 53306
rect 35078 53254 35124 53306
rect 35148 53254 35194 53306
rect 35194 53254 35204 53306
rect 35228 53254 35258 53306
rect 35258 53254 35284 53306
rect 34988 53252 35044 53254
rect 35068 53252 35124 53254
rect 35148 53252 35204 53254
rect 35228 53252 35284 53254
rect 34988 51974 35044 51976
rect 35068 51974 35124 51976
rect 35148 51974 35204 51976
rect 35228 51974 35284 51976
rect 34988 51922 35014 51974
rect 35014 51922 35044 51974
rect 35068 51922 35078 51974
rect 35078 51922 35124 51974
rect 35148 51922 35194 51974
rect 35194 51922 35204 51974
rect 35228 51922 35258 51974
rect 35258 51922 35284 51974
rect 34988 51920 35044 51922
rect 35068 51920 35124 51922
rect 35148 51920 35204 51922
rect 35228 51920 35284 51922
rect 34988 50642 35044 50644
rect 35068 50642 35124 50644
rect 35148 50642 35204 50644
rect 35228 50642 35284 50644
rect 34988 50590 35014 50642
rect 35014 50590 35044 50642
rect 35068 50590 35078 50642
rect 35078 50590 35124 50642
rect 35148 50590 35194 50642
rect 35194 50590 35204 50642
rect 35228 50590 35258 50642
rect 35258 50590 35284 50642
rect 34988 50588 35044 50590
rect 35068 50588 35124 50590
rect 35148 50588 35204 50590
rect 35228 50588 35284 50590
rect 34988 49310 35044 49312
rect 35068 49310 35124 49312
rect 35148 49310 35204 49312
rect 35228 49310 35284 49312
rect 34988 49258 35014 49310
rect 35014 49258 35044 49310
rect 35068 49258 35078 49310
rect 35078 49258 35124 49310
rect 35148 49258 35194 49310
rect 35194 49258 35204 49310
rect 35228 49258 35258 49310
rect 35258 49258 35284 49310
rect 34988 49256 35044 49258
rect 35068 49256 35124 49258
rect 35148 49256 35204 49258
rect 35228 49256 35284 49258
rect 34988 47978 35044 47980
rect 35068 47978 35124 47980
rect 35148 47978 35204 47980
rect 35228 47978 35284 47980
rect 34988 47926 35014 47978
rect 35014 47926 35044 47978
rect 35068 47926 35078 47978
rect 35078 47926 35124 47978
rect 35148 47926 35194 47978
rect 35194 47926 35204 47978
rect 35228 47926 35258 47978
rect 35258 47926 35284 47978
rect 34988 47924 35044 47926
rect 35068 47924 35124 47926
rect 35148 47924 35204 47926
rect 35228 47924 35284 47926
rect 33044 6262 33100 6318
rect 33812 6706 33868 6762
rect 34988 46646 35044 46648
rect 35068 46646 35124 46648
rect 35148 46646 35204 46648
rect 35228 46646 35284 46648
rect 34988 46594 35014 46646
rect 35014 46594 35044 46646
rect 35068 46594 35078 46646
rect 35078 46594 35124 46646
rect 35148 46594 35194 46646
rect 35194 46594 35204 46646
rect 35228 46594 35258 46646
rect 35258 46594 35284 46646
rect 34988 46592 35044 46594
rect 35068 46592 35124 46594
rect 35148 46592 35204 46594
rect 35228 46592 35284 46594
rect 34988 45314 35044 45316
rect 35068 45314 35124 45316
rect 35148 45314 35204 45316
rect 35228 45314 35284 45316
rect 34988 45262 35014 45314
rect 35014 45262 35044 45314
rect 35068 45262 35078 45314
rect 35078 45262 35124 45314
rect 35148 45262 35194 45314
rect 35194 45262 35204 45314
rect 35228 45262 35258 45314
rect 35258 45262 35284 45314
rect 34988 45260 35044 45262
rect 35068 45260 35124 45262
rect 35148 45260 35204 45262
rect 35228 45260 35284 45262
rect 34988 43982 35044 43984
rect 35068 43982 35124 43984
rect 35148 43982 35204 43984
rect 35228 43982 35284 43984
rect 34988 43930 35014 43982
rect 35014 43930 35044 43982
rect 35068 43930 35078 43982
rect 35078 43930 35124 43982
rect 35148 43930 35194 43982
rect 35194 43930 35204 43982
rect 35228 43930 35258 43982
rect 35258 43930 35284 43982
rect 34988 43928 35044 43930
rect 35068 43928 35124 43930
rect 35148 43928 35204 43930
rect 35228 43928 35284 43930
rect 34988 42650 35044 42652
rect 35068 42650 35124 42652
rect 35148 42650 35204 42652
rect 35228 42650 35284 42652
rect 34988 42598 35014 42650
rect 35014 42598 35044 42650
rect 35068 42598 35078 42650
rect 35078 42598 35124 42650
rect 35148 42598 35194 42650
rect 35194 42598 35204 42650
rect 35228 42598 35258 42650
rect 35258 42598 35284 42650
rect 34988 42596 35044 42598
rect 35068 42596 35124 42598
rect 35148 42596 35204 42598
rect 35228 42596 35284 42598
rect 34988 41318 35044 41320
rect 35068 41318 35124 41320
rect 35148 41318 35204 41320
rect 35228 41318 35284 41320
rect 34988 41266 35014 41318
rect 35014 41266 35044 41318
rect 35068 41266 35078 41318
rect 35078 41266 35124 41318
rect 35148 41266 35194 41318
rect 35194 41266 35204 41318
rect 35228 41266 35258 41318
rect 35258 41266 35284 41318
rect 34988 41264 35044 41266
rect 35068 41264 35124 41266
rect 35148 41264 35204 41266
rect 35228 41264 35284 41266
rect 34988 39986 35044 39988
rect 35068 39986 35124 39988
rect 35148 39986 35204 39988
rect 35228 39986 35284 39988
rect 34988 39934 35014 39986
rect 35014 39934 35044 39986
rect 35068 39934 35078 39986
rect 35078 39934 35124 39986
rect 35148 39934 35194 39986
rect 35194 39934 35204 39986
rect 35228 39934 35258 39986
rect 35258 39934 35284 39986
rect 34988 39932 35044 39934
rect 35068 39932 35124 39934
rect 35148 39932 35204 39934
rect 35228 39932 35284 39934
rect 34988 38654 35044 38656
rect 35068 38654 35124 38656
rect 35148 38654 35204 38656
rect 35228 38654 35284 38656
rect 34988 38602 35014 38654
rect 35014 38602 35044 38654
rect 35068 38602 35078 38654
rect 35078 38602 35124 38654
rect 35148 38602 35194 38654
rect 35194 38602 35204 38654
rect 35228 38602 35258 38654
rect 35258 38602 35284 38654
rect 34988 38600 35044 38602
rect 35068 38600 35124 38602
rect 35148 38600 35204 38602
rect 35228 38600 35284 38602
rect 34988 37322 35044 37324
rect 35068 37322 35124 37324
rect 35148 37322 35204 37324
rect 35228 37322 35284 37324
rect 34988 37270 35014 37322
rect 35014 37270 35044 37322
rect 35068 37270 35078 37322
rect 35078 37270 35124 37322
rect 35148 37270 35194 37322
rect 35194 37270 35204 37322
rect 35228 37270 35258 37322
rect 35258 37270 35284 37322
rect 34988 37268 35044 37270
rect 35068 37268 35124 37270
rect 35148 37268 35204 37270
rect 35228 37268 35284 37270
rect 34988 35990 35044 35992
rect 35068 35990 35124 35992
rect 35148 35990 35204 35992
rect 35228 35990 35284 35992
rect 34988 35938 35014 35990
rect 35014 35938 35044 35990
rect 35068 35938 35078 35990
rect 35078 35938 35124 35990
rect 35148 35938 35194 35990
rect 35194 35938 35204 35990
rect 35228 35938 35258 35990
rect 35258 35938 35284 35990
rect 34988 35936 35044 35938
rect 35068 35936 35124 35938
rect 35148 35936 35204 35938
rect 35228 35936 35284 35938
rect 34988 34658 35044 34660
rect 35068 34658 35124 34660
rect 35148 34658 35204 34660
rect 35228 34658 35284 34660
rect 34988 34606 35014 34658
rect 35014 34606 35044 34658
rect 35068 34606 35078 34658
rect 35078 34606 35124 34658
rect 35148 34606 35194 34658
rect 35194 34606 35204 34658
rect 35228 34606 35258 34658
rect 35258 34606 35284 34658
rect 34988 34604 35044 34606
rect 35068 34604 35124 34606
rect 35148 34604 35204 34606
rect 35228 34604 35284 34606
rect 34988 33326 35044 33328
rect 35068 33326 35124 33328
rect 35148 33326 35204 33328
rect 35228 33326 35284 33328
rect 34988 33274 35014 33326
rect 35014 33274 35044 33326
rect 35068 33274 35078 33326
rect 35078 33274 35124 33326
rect 35148 33274 35194 33326
rect 35194 33274 35204 33326
rect 35228 33274 35258 33326
rect 35258 33274 35284 33326
rect 34988 33272 35044 33274
rect 35068 33272 35124 33274
rect 35148 33272 35204 33274
rect 35228 33272 35284 33274
rect 33716 3302 33772 3358
rect 34292 3746 34348 3802
rect 34988 31994 35044 31996
rect 35068 31994 35124 31996
rect 35148 31994 35204 31996
rect 35228 31994 35284 31996
rect 34988 31942 35014 31994
rect 35014 31942 35044 31994
rect 35068 31942 35078 31994
rect 35078 31942 35124 31994
rect 35148 31942 35194 31994
rect 35194 31942 35204 31994
rect 35228 31942 35258 31994
rect 35258 31942 35284 31994
rect 34988 31940 35044 31942
rect 35068 31940 35124 31942
rect 35148 31940 35204 31942
rect 35228 31940 35284 31942
rect 34988 30662 35044 30664
rect 35068 30662 35124 30664
rect 35148 30662 35204 30664
rect 35228 30662 35284 30664
rect 34988 30610 35014 30662
rect 35014 30610 35044 30662
rect 35068 30610 35078 30662
rect 35078 30610 35124 30662
rect 35148 30610 35194 30662
rect 35194 30610 35204 30662
rect 35228 30610 35258 30662
rect 35258 30610 35284 30662
rect 34988 30608 35044 30610
rect 35068 30608 35124 30610
rect 35148 30608 35204 30610
rect 35228 30608 35284 30610
rect 34988 29330 35044 29332
rect 35068 29330 35124 29332
rect 35148 29330 35204 29332
rect 35228 29330 35284 29332
rect 34988 29278 35014 29330
rect 35014 29278 35044 29330
rect 35068 29278 35078 29330
rect 35078 29278 35124 29330
rect 35148 29278 35194 29330
rect 35194 29278 35204 29330
rect 35228 29278 35258 29330
rect 35258 29278 35284 29330
rect 34988 29276 35044 29278
rect 35068 29276 35124 29278
rect 35148 29276 35204 29278
rect 35228 29276 35284 29278
rect 34988 27998 35044 28000
rect 35068 27998 35124 28000
rect 35148 27998 35204 28000
rect 35228 27998 35284 28000
rect 34988 27946 35014 27998
rect 35014 27946 35044 27998
rect 35068 27946 35078 27998
rect 35078 27946 35124 27998
rect 35148 27946 35194 27998
rect 35194 27946 35204 27998
rect 35228 27946 35258 27998
rect 35258 27946 35284 27998
rect 34988 27944 35044 27946
rect 35068 27944 35124 27946
rect 35148 27944 35204 27946
rect 35228 27944 35284 27946
rect 34988 26666 35044 26668
rect 35068 26666 35124 26668
rect 35148 26666 35204 26668
rect 35228 26666 35284 26668
rect 34988 26614 35014 26666
rect 35014 26614 35044 26666
rect 35068 26614 35078 26666
rect 35078 26614 35124 26666
rect 35148 26614 35194 26666
rect 35194 26614 35204 26666
rect 35228 26614 35258 26666
rect 35258 26614 35284 26666
rect 34988 26612 35044 26614
rect 35068 26612 35124 26614
rect 35148 26612 35204 26614
rect 35228 26612 35284 26614
rect 34988 25334 35044 25336
rect 35068 25334 35124 25336
rect 35148 25334 35204 25336
rect 35228 25334 35284 25336
rect 34988 25282 35014 25334
rect 35014 25282 35044 25334
rect 35068 25282 35078 25334
rect 35078 25282 35124 25334
rect 35148 25282 35194 25334
rect 35194 25282 35204 25334
rect 35228 25282 35258 25334
rect 35258 25282 35284 25334
rect 34988 25280 35044 25282
rect 35068 25280 35124 25282
rect 35148 25280 35204 25282
rect 35228 25280 35284 25282
rect 34988 24002 35044 24004
rect 35068 24002 35124 24004
rect 35148 24002 35204 24004
rect 35228 24002 35284 24004
rect 34988 23950 35014 24002
rect 35014 23950 35044 24002
rect 35068 23950 35078 24002
rect 35078 23950 35124 24002
rect 35148 23950 35194 24002
rect 35194 23950 35204 24002
rect 35228 23950 35258 24002
rect 35258 23950 35284 24002
rect 34988 23948 35044 23950
rect 35068 23948 35124 23950
rect 35148 23948 35204 23950
rect 35228 23948 35284 23950
rect 34988 22670 35044 22672
rect 35068 22670 35124 22672
rect 35148 22670 35204 22672
rect 35228 22670 35284 22672
rect 34988 22618 35014 22670
rect 35014 22618 35044 22670
rect 35068 22618 35078 22670
rect 35078 22618 35124 22670
rect 35148 22618 35194 22670
rect 35194 22618 35204 22670
rect 35228 22618 35258 22670
rect 35258 22618 35284 22670
rect 34988 22616 35044 22618
rect 35068 22616 35124 22618
rect 35148 22616 35204 22618
rect 35228 22616 35284 22618
rect 34988 21338 35044 21340
rect 35068 21338 35124 21340
rect 35148 21338 35204 21340
rect 35228 21338 35284 21340
rect 34988 21286 35014 21338
rect 35014 21286 35044 21338
rect 35068 21286 35078 21338
rect 35078 21286 35124 21338
rect 35148 21286 35194 21338
rect 35194 21286 35204 21338
rect 35228 21286 35258 21338
rect 35258 21286 35284 21338
rect 34988 21284 35044 21286
rect 35068 21284 35124 21286
rect 35148 21284 35204 21286
rect 35228 21284 35284 21286
rect 34988 20006 35044 20008
rect 35068 20006 35124 20008
rect 35148 20006 35204 20008
rect 35228 20006 35284 20008
rect 34988 19954 35014 20006
rect 35014 19954 35044 20006
rect 35068 19954 35078 20006
rect 35078 19954 35124 20006
rect 35148 19954 35194 20006
rect 35194 19954 35204 20006
rect 35228 19954 35258 20006
rect 35258 19954 35284 20006
rect 34988 19952 35044 19954
rect 35068 19952 35124 19954
rect 35148 19952 35204 19954
rect 35228 19952 35284 19954
rect 34988 18674 35044 18676
rect 35068 18674 35124 18676
rect 35148 18674 35204 18676
rect 35228 18674 35284 18676
rect 34988 18622 35014 18674
rect 35014 18622 35044 18674
rect 35068 18622 35078 18674
rect 35078 18622 35124 18674
rect 35148 18622 35194 18674
rect 35194 18622 35204 18674
rect 35228 18622 35258 18674
rect 35258 18622 35284 18674
rect 34988 18620 35044 18622
rect 35068 18620 35124 18622
rect 35148 18620 35204 18622
rect 35228 18620 35284 18622
rect 34988 17342 35044 17344
rect 35068 17342 35124 17344
rect 35148 17342 35204 17344
rect 35228 17342 35284 17344
rect 34988 17290 35014 17342
rect 35014 17290 35044 17342
rect 35068 17290 35078 17342
rect 35078 17290 35124 17342
rect 35148 17290 35194 17342
rect 35194 17290 35204 17342
rect 35228 17290 35258 17342
rect 35258 17290 35284 17342
rect 34988 17288 35044 17290
rect 35068 17288 35124 17290
rect 35148 17288 35204 17290
rect 35228 17288 35284 17290
rect 34988 16010 35044 16012
rect 35068 16010 35124 16012
rect 35148 16010 35204 16012
rect 35228 16010 35284 16012
rect 34988 15958 35014 16010
rect 35014 15958 35044 16010
rect 35068 15958 35078 16010
rect 35078 15958 35124 16010
rect 35148 15958 35194 16010
rect 35194 15958 35204 16010
rect 35228 15958 35258 16010
rect 35258 15958 35284 16010
rect 34988 15956 35044 15958
rect 35068 15956 35124 15958
rect 35148 15956 35204 15958
rect 35228 15956 35284 15958
rect 34988 14678 35044 14680
rect 35068 14678 35124 14680
rect 35148 14678 35204 14680
rect 35228 14678 35284 14680
rect 34988 14626 35014 14678
rect 35014 14626 35044 14678
rect 35068 14626 35078 14678
rect 35078 14626 35124 14678
rect 35148 14626 35194 14678
rect 35194 14626 35204 14678
rect 35228 14626 35258 14678
rect 35258 14626 35284 14678
rect 34988 14624 35044 14626
rect 35068 14624 35124 14626
rect 35148 14624 35204 14626
rect 35228 14624 35284 14626
rect 34988 13346 35044 13348
rect 35068 13346 35124 13348
rect 35148 13346 35204 13348
rect 35228 13346 35284 13348
rect 34988 13294 35014 13346
rect 35014 13294 35044 13346
rect 35068 13294 35078 13346
rect 35078 13294 35124 13346
rect 35148 13294 35194 13346
rect 35194 13294 35204 13346
rect 35228 13294 35258 13346
rect 35258 13294 35284 13346
rect 34988 13292 35044 13294
rect 35068 13292 35124 13294
rect 35148 13292 35204 13294
rect 35228 13292 35284 13294
rect 34988 12014 35044 12016
rect 35068 12014 35124 12016
rect 35148 12014 35204 12016
rect 35228 12014 35284 12016
rect 34988 11962 35014 12014
rect 35014 11962 35044 12014
rect 35068 11962 35078 12014
rect 35078 11962 35124 12014
rect 35148 11962 35194 12014
rect 35194 11962 35204 12014
rect 35228 11962 35258 12014
rect 35258 11962 35284 12014
rect 34988 11960 35044 11962
rect 35068 11960 35124 11962
rect 35148 11960 35204 11962
rect 35228 11960 35284 11962
rect 34988 10682 35044 10684
rect 35068 10682 35124 10684
rect 35148 10682 35204 10684
rect 35228 10682 35284 10684
rect 34988 10630 35014 10682
rect 35014 10630 35044 10682
rect 35068 10630 35078 10682
rect 35078 10630 35124 10682
rect 35148 10630 35194 10682
rect 35194 10630 35204 10682
rect 35228 10630 35258 10682
rect 35258 10630 35284 10682
rect 34988 10628 35044 10630
rect 35068 10628 35124 10630
rect 35148 10628 35204 10630
rect 35228 10628 35284 10630
rect 34988 9350 35044 9352
rect 35068 9350 35124 9352
rect 35148 9350 35204 9352
rect 35228 9350 35284 9352
rect 34988 9298 35014 9350
rect 35014 9298 35044 9350
rect 35068 9298 35078 9350
rect 35078 9298 35124 9350
rect 35148 9298 35194 9350
rect 35194 9298 35204 9350
rect 35228 9298 35258 9350
rect 35258 9298 35284 9350
rect 34988 9296 35044 9298
rect 35068 9296 35124 9298
rect 35148 9296 35204 9298
rect 35228 9296 35284 9298
rect 34988 8018 35044 8020
rect 35068 8018 35124 8020
rect 35148 8018 35204 8020
rect 35228 8018 35284 8020
rect 34988 7966 35014 8018
rect 35014 7966 35044 8018
rect 35068 7966 35078 8018
rect 35078 7966 35124 8018
rect 35148 7966 35194 8018
rect 35194 7966 35204 8018
rect 35228 7966 35258 8018
rect 35258 7966 35284 8018
rect 34988 7964 35044 7966
rect 35068 7964 35124 7966
rect 35148 7964 35204 7966
rect 35228 7964 35284 7966
rect 34580 6706 34636 6762
rect 34676 6427 34732 6466
rect 34676 6410 34678 6427
rect 34678 6410 34730 6427
rect 34730 6410 34732 6427
rect 35444 6745 35446 6762
rect 35446 6745 35498 6762
rect 35498 6745 35500 6762
rect 35444 6706 35500 6745
rect 34988 6686 35044 6688
rect 35068 6686 35124 6688
rect 35148 6686 35204 6688
rect 35228 6686 35284 6688
rect 34988 6634 35014 6686
rect 35014 6634 35044 6686
rect 35068 6634 35078 6686
rect 35078 6634 35124 6686
rect 35148 6634 35194 6686
rect 35194 6634 35204 6686
rect 35228 6634 35258 6686
rect 35258 6634 35284 6686
rect 34988 6632 35044 6634
rect 35068 6632 35124 6634
rect 35148 6632 35204 6634
rect 35228 6632 35284 6634
rect 34988 5354 35044 5356
rect 35068 5354 35124 5356
rect 35148 5354 35204 5356
rect 35228 5354 35284 5356
rect 34988 5302 35014 5354
rect 35014 5302 35044 5354
rect 35068 5302 35078 5354
rect 35078 5302 35124 5354
rect 35148 5302 35194 5354
rect 35194 5302 35204 5354
rect 35228 5302 35258 5354
rect 35258 5302 35284 5354
rect 34988 5300 35044 5302
rect 35068 5300 35124 5302
rect 35148 5300 35204 5302
rect 35228 5300 35284 5302
rect 34988 4022 35044 4024
rect 35068 4022 35124 4024
rect 35148 4022 35204 4024
rect 35228 4022 35284 4024
rect 34988 3970 35014 4022
rect 35014 3970 35044 4022
rect 35068 3970 35078 4022
rect 35078 3970 35124 4022
rect 35148 3970 35194 4022
rect 35194 3970 35204 4022
rect 35228 3970 35258 4022
rect 35258 3970 35284 4022
rect 34988 3968 35044 3970
rect 35068 3968 35124 3970
rect 35148 3968 35204 3970
rect 35228 3968 35284 3970
rect 34988 2690 35044 2692
rect 35068 2690 35124 2692
rect 35148 2690 35204 2692
rect 35228 2690 35284 2692
rect 34988 2638 35014 2690
rect 35014 2638 35044 2690
rect 35068 2638 35078 2690
rect 35078 2638 35124 2690
rect 35148 2638 35194 2690
rect 35194 2638 35204 2690
rect 35228 2638 35258 2690
rect 35258 2638 35284 2690
rect 34988 2636 35044 2638
rect 35068 2636 35124 2638
rect 35148 2636 35204 2638
rect 35228 2636 35284 2638
rect 38132 7890 38188 7946
rect 38132 7594 38188 7650
rect 39380 7298 39436 7354
rect 39284 6706 39340 6762
rect 40340 8186 40396 8242
rect 40724 5818 40780 5874
rect 41876 6410 41932 6466
rect 42356 6745 42358 6762
rect 42358 6745 42410 6762
rect 42410 6745 42412 6762
rect 42356 6706 42412 6745
rect 42356 6114 42412 6170
rect 43700 6279 43756 6318
rect 43700 6262 43702 6279
rect 43702 6262 43754 6279
rect 43754 6262 43756 6279
rect 44180 8038 44236 8094
rect 46100 8186 46156 8242
rect 50348 56636 50404 56638
rect 50428 56636 50484 56638
rect 50508 56636 50564 56638
rect 50588 56636 50644 56638
rect 50348 56584 50374 56636
rect 50374 56584 50404 56636
rect 50428 56584 50438 56636
rect 50438 56584 50484 56636
rect 50508 56584 50554 56636
rect 50554 56584 50564 56636
rect 50588 56584 50618 56636
rect 50618 56584 50644 56636
rect 50348 56582 50404 56584
rect 50428 56582 50484 56584
rect 50508 56582 50564 56584
rect 50588 56582 50644 56584
rect 46484 8186 46540 8242
rect 47924 8038 47980 8094
rect 46292 7002 46348 7058
rect 46388 5966 46444 6022
rect 50348 55304 50404 55306
rect 50428 55304 50484 55306
rect 50508 55304 50564 55306
rect 50588 55304 50644 55306
rect 50348 55252 50374 55304
rect 50374 55252 50404 55304
rect 50428 55252 50438 55304
rect 50438 55252 50484 55304
rect 50508 55252 50554 55304
rect 50554 55252 50564 55304
rect 50588 55252 50618 55304
rect 50618 55252 50644 55304
rect 50348 55250 50404 55252
rect 50428 55250 50484 55252
rect 50508 55250 50564 55252
rect 50588 55250 50644 55252
rect 48500 6706 48556 6762
rect 50036 7890 50092 7946
rect 50348 53972 50404 53974
rect 50428 53972 50484 53974
rect 50508 53972 50564 53974
rect 50588 53972 50644 53974
rect 50348 53920 50374 53972
rect 50374 53920 50404 53972
rect 50428 53920 50438 53972
rect 50438 53920 50484 53972
rect 50508 53920 50554 53972
rect 50554 53920 50564 53972
rect 50588 53920 50618 53972
rect 50618 53920 50644 53972
rect 50348 53918 50404 53920
rect 50428 53918 50484 53920
rect 50508 53918 50564 53920
rect 50588 53918 50644 53920
rect 50348 52640 50404 52642
rect 50428 52640 50484 52642
rect 50508 52640 50564 52642
rect 50588 52640 50644 52642
rect 50348 52588 50374 52640
rect 50374 52588 50404 52640
rect 50428 52588 50438 52640
rect 50438 52588 50484 52640
rect 50508 52588 50554 52640
rect 50554 52588 50564 52640
rect 50588 52588 50618 52640
rect 50618 52588 50644 52640
rect 50348 52586 50404 52588
rect 50428 52586 50484 52588
rect 50508 52586 50564 52588
rect 50588 52586 50644 52588
rect 50348 51308 50404 51310
rect 50428 51308 50484 51310
rect 50508 51308 50564 51310
rect 50588 51308 50644 51310
rect 50348 51256 50374 51308
rect 50374 51256 50404 51308
rect 50428 51256 50438 51308
rect 50438 51256 50484 51308
rect 50508 51256 50554 51308
rect 50554 51256 50564 51308
rect 50588 51256 50618 51308
rect 50618 51256 50644 51308
rect 50348 51254 50404 51256
rect 50428 51254 50484 51256
rect 50508 51254 50564 51256
rect 50588 51254 50644 51256
rect 50348 49976 50404 49978
rect 50428 49976 50484 49978
rect 50508 49976 50564 49978
rect 50588 49976 50644 49978
rect 50348 49924 50374 49976
rect 50374 49924 50404 49976
rect 50428 49924 50438 49976
rect 50438 49924 50484 49976
rect 50508 49924 50554 49976
rect 50554 49924 50564 49976
rect 50588 49924 50618 49976
rect 50618 49924 50644 49976
rect 50348 49922 50404 49924
rect 50428 49922 50484 49924
rect 50508 49922 50564 49924
rect 50588 49922 50644 49924
rect 50348 48644 50404 48646
rect 50428 48644 50484 48646
rect 50508 48644 50564 48646
rect 50588 48644 50644 48646
rect 50348 48592 50374 48644
rect 50374 48592 50404 48644
rect 50428 48592 50438 48644
rect 50438 48592 50484 48644
rect 50508 48592 50554 48644
rect 50554 48592 50564 48644
rect 50588 48592 50618 48644
rect 50618 48592 50644 48644
rect 50348 48590 50404 48592
rect 50428 48590 50484 48592
rect 50508 48590 50564 48592
rect 50588 48590 50644 48592
rect 50348 47312 50404 47314
rect 50428 47312 50484 47314
rect 50508 47312 50564 47314
rect 50588 47312 50644 47314
rect 50348 47260 50374 47312
rect 50374 47260 50404 47312
rect 50428 47260 50438 47312
rect 50438 47260 50484 47312
rect 50508 47260 50554 47312
rect 50554 47260 50564 47312
rect 50588 47260 50618 47312
rect 50618 47260 50644 47312
rect 50348 47258 50404 47260
rect 50428 47258 50484 47260
rect 50508 47258 50564 47260
rect 50588 47258 50644 47260
rect 50348 45980 50404 45982
rect 50428 45980 50484 45982
rect 50508 45980 50564 45982
rect 50588 45980 50644 45982
rect 50348 45928 50374 45980
rect 50374 45928 50404 45980
rect 50428 45928 50438 45980
rect 50438 45928 50484 45980
rect 50508 45928 50554 45980
rect 50554 45928 50564 45980
rect 50588 45928 50618 45980
rect 50618 45928 50644 45980
rect 50348 45926 50404 45928
rect 50428 45926 50484 45928
rect 50508 45926 50564 45928
rect 50588 45926 50644 45928
rect 50348 44648 50404 44650
rect 50428 44648 50484 44650
rect 50508 44648 50564 44650
rect 50588 44648 50644 44650
rect 50348 44596 50374 44648
rect 50374 44596 50404 44648
rect 50428 44596 50438 44648
rect 50438 44596 50484 44648
rect 50508 44596 50554 44648
rect 50554 44596 50564 44648
rect 50588 44596 50618 44648
rect 50618 44596 50644 44648
rect 50348 44594 50404 44596
rect 50428 44594 50484 44596
rect 50508 44594 50564 44596
rect 50588 44594 50644 44596
rect 50348 43316 50404 43318
rect 50428 43316 50484 43318
rect 50508 43316 50564 43318
rect 50588 43316 50644 43318
rect 50348 43264 50374 43316
rect 50374 43264 50404 43316
rect 50428 43264 50438 43316
rect 50438 43264 50484 43316
rect 50508 43264 50554 43316
rect 50554 43264 50564 43316
rect 50588 43264 50618 43316
rect 50618 43264 50644 43316
rect 50348 43262 50404 43264
rect 50428 43262 50484 43264
rect 50508 43262 50564 43264
rect 50588 43262 50644 43264
rect 50348 41984 50404 41986
rect 50428 41984 50484 41986
rect 50508 41984 50564 41986
rect 50588 41984 50644 41986
rect 50348 41932 50374 41984
rect 50374 41932 50404 41984
rect 50428 41932 50438 41984
rect 50438 41932 50484 41984
rect 50508 41932 50554 41984
rect 50554 41932 50564 41984
rect 50588 41932 50618 41984
rect 50618 41932 50644 41984
rect 50348 41930 50404 41932
rect 50428 41930 50484 41932
rect 50508 41930 50564 41932
rect 50588 41930 50644 41932
rect 50348 40652 50404 40654
rect 50428 40652 50484 40654
rect 50508 40652 50564 40654
rect 50588 40652 50644 40654
rect 50348 40600 50374 40652
rect 50374 40600 50404 40652
rect 50428 40600 50438 40652
rect 50438 40600 50484 40652
rect 50508 40600 50554 40652
rect 50554 40600 50564 40652
rect 50588 40600 50618 40652
rect 50618 40600 50644 40652
rect 50348 40598 50404 40600
rect 50428 40598 50484 40600
rect 50508 40598 50564 40600
rect 50588 40598 50644 40600
rect 50348 39320 50404 39322
rect 50428 39320 50484 39322
rect 50508 39320 50564 39322
rect 50588 39320 50644 39322
rect 50348 39268 50374 39320
rect 50374 39268 50404 39320
rect 50428 39268 50438 39320
rect 50438 39268 50484 39320
rect 50508 39268 50554 39320
rect 50554 39268 50564 39320
rect 50588 39268 50618 39320
rect 50618 39268 50644 39320
rect 50348 39266 50404 39268
rect 50428 39266 50484 39268
rect 50508 39266 50564 39268
rect 50588 39266 50644 39268
rect 50348 37988 50404 37990
rect 50428 37988 50484 37990
rect 50508 37988 50564 37990
rect 50588 37988 50644 37990
rect 50348 37936 50374 37988
rect 50374 37936 50404 37988
rect 50428 37936 50438 37988
rect 50438 37936 50484 37988
rect 50508 37936 50554 37988
rect 50554 37936 50564 37988
rect 50588 37936 50618 37988
rect 50618 37936 50644 37988
rect 50348 37934 50404 37936
rect 50428 37934 50484 37936
rect 50508 37934 50564 37936
rect 50588 37934 50644 37936
rect 50348 36656 50404 36658
rect 50428 36656 50484 36658
rect 50508 36656 50564 36658
rect 50588 36656 50644 36658
rect 50348 36604 50374 36656
rect 50374 36604 50404 36656
rect 50428 36604 50438 36656
rect 50438 36604 50484 36656
rect 50508 36604 50554 36656
rect 50554 36604 50564 36656
rect 50588 36604 50618 36656
rect 50618 36604 50644 36656
rect 50348 36602 50404 36604
rect 50428 36602 50484 36604
rect 50508 36602 50564 36604
rect 50588 36602 50644 36604
rect 50348 35324 50404 35326
rect 50428 35324 50484 35326
rect 50508 35324 50564 35326
rect 50588 35324 50644 35326
rect 50348 35272 50374 35324
rect 50374 35272 50404 35324
rect 50428 35272 50438 35324
rect 50438 35272 50484 35324
rect 50508 35272 50554 35324
rect 50554 35272 50564 35324
rect 50588 35272 50618 35324
rect 50618 35272 50644 35324
rect 50348 35270 50404 35272
rect 50428 35270 50484 35272
rect 50508 35270 50564 35272
rect 50588 35270 50644 35272
rect 50348 33992 50404 33994
rect 50428 33992 50484 33994
rect 50508 33992 50564 33994
rect 50588 33992 50644 33994
rect 50348 33940 50374 33992
rect 50374 33940 50404 33992
rect 50428 33940 50438 33992
rect 50438 33940 50484 33992
rect 50508 33940 50554 33992
rect 50554 33940 50564 33992
rect 50588 33940 50618 33992
rect 50618 33940 50644 33992
rect 50348 33938 50404 33940
rect 50428 33938 50484 33940
rect 50508 33938 50564 33940
rect 50588 33938 50644 33940
rect 50348 32660 50404 32662
rect 50428 32660 50484 32662
rect 50508 32660 50564 32662
rect 50588 32660 50644 32662
rect 50348 32608 50374 32660
rect 50374 32608 50404 32660
rect 50428 32608 50438 32660
rect 50438 32608 50484 32660
rect 50508 32608 50554 32660
rect 50554 32608 50564 32660
rect 50588 32608 50618 32660
rect 50618 32608 50644 32660
rect 50348 32606 50404 32608
rect 50428 32606 50484 32608
rect 50508 32606 50564 32608
rect 50588 32606 50644 32608
rect 50348 31328 50404 31330
rect 50428 31328 50484 31330
rect 50508 31328 50564 31330
rect 50588 31328 50644 31330
rect 50348 31276 50374 31328
rect 50374 31276 50404 31328
rect 50428 31276 50438 31328
rect 50438 31276 50484 31328
rect 50508 31276 50554 31328
rect 50554 31276 50564 31328
rect 50588 31276 50618 31328
rect 50618 31276 50644 31328
rect 50348 31274 50404 31276
rect 50428 31274 50484 31276
rect 50508 31274 50564 31276
rect 50588 31274 50644 31276
rect 50348 29996 50404 29998
rect 50428 29996 50484 29998
rect 50508 29996 50564 29998
rect 50588 29996 50644 29998
rect 50348 29944 50374 29996
rect 50374 29944 50404 29996
rect 50428 29944 50438 29996
rect 50438 29944 50484 29996
rect 50508 29944 50554 29996
rect 50554 29944 50564 29996
rect 50588 29944 50618 29996
rect 50618 29944 50644 29996
rect 50348 29942 50404 29944
rect 50428 29942 50484 29944
rect 50508 29942 50564 29944
rect 50588 29942 50644 29944
rect 50348 28664 50404 28666
rect 50428 28664 50484 28666
rect 50508 28664 50564 28666
rect 50588 28664 50644 28666
rect 50348 28612 50374 28664
rect 50374 28612 50404 28664
rect 50428 28612 50438 28664
rect 50438 28612 50484 28664
rect 50508 28612 50554 28664
rect 50554 28612 50564 28664
rect 50588 28612 50618 28664
rect 50618 28612 50644 28664
rect 50348 28610 50404 28612
rect 50428 28610 50484 28612
rect 50508 28610 50564 28612
rect 50588 28610 50644 28612
rect 50348 27332 50404 27334
rect 50428 27332 50484 27334
rect 50508 27332 50564 27334
rect 50588 27332 50644 27334
rect 50348 27280 50374 27332
rect 50374 27280 50404 27332
rect 50428 27280 50438 27332
rect 50438 27280 50484 27332
rect 50508 27280 50554 27332
rect 50554 27280 50564 27332
rect 50588 27280 50618 27332
rect 50618 27280 50644 27332
rect 50348 27278 50404 27280
rect 50428 27278 50484 27280
rect 50508 27278 50564 27280
rect 50588 27278 50644 27280
rect 50348 26000 50404 26002
rect 50428 26000 50484 26002
rect 50508 26000 50564 26002
rect 50588 26000 50644 26002
rect 50348 25948 50374 26000
rect 50374 25948 50404 26000
rect 50428 25948 50438 26000
rect 50438 25948 50484 26000
rect 50508 25948 50554 26000
rect 50554 25948 50564 26000
rect 50588 25948 50618 26000
rect 50618 25948 50644 26000
rect 50348 25946 50404 25948
rect 50428 25946 50484 25948
rect 50508 25946 50564 25948
rect 50588 25946 50644 25948
rect 50348 24668 50404 24670
rect 50428 24668 50484 24670
rect 50508 24668 50564 24670
rect 50588 24668 50644 24670
rect 50348 24616 50374 24668
rect 50374 24616 50404 24668
rect 50428 24616 50438 24668
rect 50438 24616 50484 24668
rect 50508 24616 50554 24668
rect 50554 24616 50564 24668
rect 50588 24616 50618 24668
rect 50618 24616 50644 24668
rect 50348 24614 50404 24616
rect 50428 24614 50484 24616
rect 50508 24614 50564 24616
rect 50588 24614 50644 24616
rect 50348 23336 50404 23338
rect 50428 23336 50484 23338
rect 50508 23336 50564 23338
rect 50588 23336 50644 23338
rect 50348 23284 50374 23336
rect 50374 23284 50404 23336
rect 50428 23284 50438 23336
rect 50438 23284 50484 23336
rect 50508 23284 50554 23336
rect 50554 23284 50564 23336
rect 50588 23284 50618 23336
rect 50618 23284 50644 23336
rect 50348 23282 50404 23284
rect 50428 23282 50484 23284
rect 50508 23282 50564 23284
rect 50588 23282 50644 23284
rect 50348 22004 50404 22006
rect 50428 22004 50484 22006
rect 50508 22004 50564 22006
rect 50588 22004 50644 22006
rect 50348 21952 50374 22004
rect 50374 21952 50404 22004
rect 50428 21952 50438 22004
rect 50438 21952 50484 22004
rect 50508 21952 50554 22004
rect 50554 21952 50564 22004
rect 50588 21952 50618 22004
rect 50618 21952 50644 22004
rect 50348 21950 50404 21952
rect 50428 21950 50484 21952
rect 50508 21950 50564 21952
rect 50588 21950 50644 21952
rect 50348 20672 50404 20674
rect 50428 20672 50484 20674
rect 50508 20672 50564 20674
rect 50588 20672 50644 20674
rect 50348 20620 50374 20672
rect 50374 20620 50404 20672
rect 50428 20620 50438 20672
rect 50438 20620 50484 20672
rect 50508 20620 50554 20672
rect 50554 20620 50564 20672
rect 50588 20620 50618 20672
rect 50618 20620 50644 20672
rect 50348 20618 50404 20620
rect 50428 20618 50484 20620
rect 50508 20618 50564 20620
rect 50588 20618 50644 20620
rect 50348 19340 50404 19342
rect 50428 19340 50484 19342
rect 50508 19340 50564 19342
rect 50588 19340 50644 19342
rect 50348 19288 50374 19340
rect 50374 19288 50404 19340
rect 50428 19288 50438 19340
rect 50438 19288 50484 19340
rect 50508 19288 50554 19340
rect 50554 19288 50564 19340
rect 50588 19288 50618 19340
rect 50618 19288 50644 19340
rect 50348 19286 50404 19288
rect 50428 19286 50484 19288
rect 50508 19286 50564 19288
rect 50588 19286 50644 19288
rect 50348 18008 50404 18010
rect 50428 18008 50484 18010
rect 50508 18008 50564 18010
rect 50588 18008 50644 18010
rect 50348 17956 50374 18008
rect 50374 17956 50404 18008
rect 50428 17956 50438 18008
rect 50438 17956 50484 18008
rect 50508 17956 50554 18008
rect 50554 17956 50564 18008
rect 50588 17956 50618 18008
rect 50618 17956 50644 18008
rect 50348 17954 50404 17956
rect 50428 17954 50484 17956
rect 50508 17954 50564 17956
rect 50588 17954 50644 17956
rect 50348 16676 50404 16678
rect 50428 16676 50484 16678
rect 50508 16676 50564 16678
rect 50588 16676 50644 16678
rect 50348 16624 50374 16676
rect 50374 16624 50404 16676
rect 50428 16624 50438 16676
rect 50438 16624 50484 16676
rect 50508 16624 50554 16676
rect 50554 16624 50564 16676
rect 50588 16624 50618 16676
rect 50618 16624 50644 16676
rect 50348 16622 50404 16624
rect 50428 16622 50484 16624
rect 50508 16622 50564 16624
rect 50588 16622 50644 16624
rect 50348 15344 50404 15346
rect 50428 15344 50484 15346
rect 50508 15344 50564 15346
rect 50588 15344 50644 15346
rect 50348 15292 50374 15344
rect 50374 15292 50404 15344
rect 50428 15292 50438 15344
rect 50438 15292 50484 15344
rect 50508 15292 50554 15344
rect 50554 15292 50564 15344
rect 50588 15292 50618 15344
rect 50618 15292 50644 15344
rect 50348 15290 50404 15292
rect 50428 15290 50484 15292
rect 50508 15290 50564 15292
rect 50588 15290 50644 15292
rect 50348 14012 50404 14014
rect 50428 14012 50484 14014
rect 50508 14012 50564 14014
rect 50588 14012 50644 14014
rect 50348 13960 50374 14012
rect 50374 13960 50404 14012
rect 50428 13960 50438 14012
rect 50438 13960 50484 14012
rect 50508 13960 50554 14012
rect 50554 13960 50564 14012
rect 50588 13960 50618 14012
rect 50618 13960 50644 14012
rect 50348 13958 50404 13960
rect 50428 13958 50484 13960
rect 50508 13958 50564 13960
rect 50588 13958 50644 13960
rect 50348 12680 50404 12682
rect 50428 12680 50484 12682
rect 50508 12680 50564 12682
rect 50588 12680 50644 12682
rect 50348 12628 50374 12680
rect 50374 12628 50404 12680
rect 50428 12628 50438 12680
rect 50438 12628 50484 12680
rect 50508 12628 50554 12680
rect 50554 12628 50564 12680
rect 50588 12628 50618 12680
rect 50618 12628 50644 12680
rect 50348 12626 50404 12628
rect 50428 12626 50484 12628
rect 50508 12626 50564 12628
rect 50588 12626 50644 12628
rect 50348 11348 50404 11350
rect 50428 11348 50484 11350
rect 50508 11348 50564 11350
rect 50588 11348 50644 11350
rect 50348 11296 50374 11348
rect 50374 11296 50404 11348
rect 50428 11296 50438 11348
rect 50438 11296 50484 11348
rect 50508 11296 50554 11348
rect 50554 11296 50564 11348
rect 50588 11296 50618 11348
rect 50618 11296 50644 11348
rect 50348 11294 50404 11296
rect 50428 11294 50484 11296
rect 50508 11294 50564 11296
rect 50588 11294 50644 11296
rect 50348 10016 50404 10018
rect 50428 10016 50484 10018
rect 50508 10016 50564 10018
rect 50588 10016 50644 10018
rect 50348 9964 50374 10016
rect 50374 9964 50404 10016
rect 50428 9964 50438 10016
rect 50438 9964 50484 10016
rect 50508 9964 50554 10016
rect 50554 9964 50564 10016
rect 50588 9964 50618 10016
rect 50618 9964 50644 10016
rect 50348 9962 50404 9964
rect 50428 9962 50484 9964
rect 50508 9962 50564 9964
rect 50588 9962 50644 9964
rect 50348 8684 50404 8686
rect 50428 8684 50484 8686
rect 50508 8684 50564 8686
rect 50588 8684 50644 8686
rect 50348 8632 50374 8684
rect 50374 8632 50404 8684
rect 50428 8632 50438 8684
rect 50438 8632 50484 8684
rect 50508 8632 50554 8684
rect 50554 8632 50564 8684
rect 50588 8632 50618 8684
rect 50618 8632 50644 8684
rect 50348 8630 50404 8632
rect 50428 8630 50484 8632
rect 50508 8630 50564 8632
rect 50588 8630 50644 8632
rect 50348 7352 50404 7354
rect 50428 7352 50484 7354
rect 50508 7352 50564 7354
rect 50588 7352 50644 7354
rect 50348 7300 50374 7352
rect 50374 7300 50404 7352
rect 50428 7300 50438 7352
rect 50438 7300 50484 7352
rect 50508 7300 50554 7352
rect 50554 7300 50564 7352
rect 50588 7300 50618 7352
rect 50618 7300 50644 7352
rect 50348 7298 50404 7300
rect 50428 7298 50484 7300
rect 50508 7298 50564 7300
rect 50588 7298 50644 7300
rect 52148 7446 52204 7502
rect 50348 6020 50404 6022
rect 50428 6020 50484 6022
rect 50508 6020 50564 6022
rect 50588 6020 50644 6022
rect 50348 5968 50374 6020
rect 50374 5968 50404 6020
rect 50428 5968 50438 6020
rect 50438 5968 50484 6020
rect 50508 5968 50554 6020
rect 50554 5968 50564 6020
rect 50588 5968 50618 6020
rect 50618 5968 50644 6020
rect 50348 5966 50404 5968
rect 50428 5966 50484 5968
rect 50508 5966 50564 5968
rect 50588 5966 50644 5968
rect 50348 4688 50404 4690
rect 50428 4688 50484 4690
rect 50508 4688 50564 4690
rect 50588 4688 50644 4690
rect 50348 4636 50374 4688
rect 50374 4636 50404 4688
rect 50428 4636 50438 4688
rect 50438 4636 50484 4688
rect 50508 4636 50554 4688
rect 50554 4636 50564 4688
rect 50588 4636 50618 4688
rect 50618 4636 50644 4688
rect 50348 4634 50404 4636
rect 50428 4634 50484 4636
rect 50508 4634 50564 4636
rect 50588 4634 50644 4636
rect 50348 3356 50404 3358
rect 50428 3356 50484 3358
rect 50508 3356 50564 3358
rect 50588 3356 50644 3358
rect 50348 3304 50374 3356
rect 50374 3304 50404 3356
rect 50428 3304 50438 3356
rect 50438 3304 50484 3356
rect 50508 3304 50554 3356
rect 50554 3304 50564 3356
rect 50588 3304 50618 3356
rect 50618 3304 50644 3356
rect 50348 3302 50404 3304
rect 50428 3302 50484 3304
rect 50508 3302 50564 3304
rect 50588 3302 50644 3304
rect 52436 8482 52492 8538
rect 52916 8351 52972 8390
rect 52916 8334 52918 8351
rect 52918 8334 52970 8351
rect 52970 8334 52972 8351
rect 52724 7150 52780 7206
rect 53588 6854 53644 6910
rect 56372 7742 56428 7798
rect 56372 3045 56374 3062
rect 56374 3045 56426 3062
rect 56426 3045 56428 3062
rect 56372 3006 56428 3045
rect 56564 4930 56620 4986
rect 56660 4634 56716 4690
<< metal3 >>
rect 4256 57308 4576 57309
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 57243 4576 57244
rect 34976 57308 35296 57309
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 57243 35296 57244
rect 19616 56642 19936 56643
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 56577 19936 56578
rect 50336 56642 50656 56643
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 56577 50656 56578
rect 7215 56196 7281 56199
rect 7354 56196 7360 56198
rect 7215 56194 7360 56196
rect 7215 56138 7220 56194
rect 7276 56138 7360 56194
rect 7215 56136 7360 56138
rect 7215 56133 7281 56136
rect 7354 56134 7360 56136
rect 7424 56134 7430 56198
rect 4256 55976 4576 55977
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 55911 4576 55912
rect 34976 55976 35296 55977
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 55911 35296 55912
rect 19616 55310 19936 55311
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 55245 19936 55246
rect 50336 55310 50656 55311
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 55245 50656 55246
rect 4256 54644 4576 54645
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 54579 4576 54580
rect 34976 54644 35296 54645
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 54579 35296 54580
rect 19616 53978 19936 53979
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 53913 19936 53914
rect 50336 53978 50656 53979
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 53913 50656 53914
rect 4256 53312 4576 53313
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 53247 4576 53248
rect 34976 53312 35296 53313
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 53247 35296 53248
rect 19616 52646 19936 52647
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 52581 19936 52582
rect 50336 52646 50656 52647
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 52581 50656 52582
rect 4256 51980 4576 51981
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 51915 4576 51916
rect 34976 51980 35296 51981
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 51915 35296 51916
rect 19616 51314 19936 51315
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 51249 19936 51250
rect 50336 51314 50656 51315
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 51249 50656 51250
rect 4256 50648 4576 50649
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 50583 4576 50584
rect 34976 50648 35296 50649
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 50583 35296 50584
rect 19616 49982 19936 49983
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 49917 19936 49918
rect 50336 49982 50656 49983
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 49917 50656 49918
rect 4256 49316 4576 49317
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 49251 4576 49252
rect 34976 49316 35296 49317
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 49251 35296 49252
rect 19616 48650 19936 48651
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 48585 19936 48586
rect 50336 48650 50656 48651
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 48585 50656 48586
rect 4256 47984 4576 47985
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 47919 4576 47920
rect 34976 47984 35296 47985
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 47919 35296 47920
rect 19616 47318 19936 47319
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 47253 19936 47254
rect 50336 47318 50656 47319
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 47253 50656 47254
rect 4256 46652 4576 46653
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 46587 4576 46588
rect 34976 46652 35296 46653
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 46587 35296 46588
rect 19616 45986 19936 45987
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 45921 19936 45922
rect 50336 45986 50656 45987
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 45921 50656 45922
rect 4256 45320 4576 45321
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 45255 4576 45256
rect 34976 45320 35296 45321
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 45255 35296 45256
rect 19616 44654 19936 44655
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 44589 19936 44590
rect 50336 44654 50656 44655
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 44589 50656 44590
rect 4256 43988 4576 43989
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 43923 4576 43924
rect 34976 43988 35296 43989
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 43923 35296 43924
rect 19616 43322 19936 43323
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 43257 19936 43258
rect 50336 43322 50656 43323
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 43257 50656 43258
rect 4256 42656 4576 42657
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 42591 4576 42592
rect 34976 42656 35296 42657
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 42591 35296 42592
rect 19616 41990 19936 41991
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 41925 19936 41926
rect 50336 41990 50656 41991
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 41925 50656 41926
rect 4256 41324 4576 41325
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 41259 4576 41260
rect 34976 41324 35296 41325
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 41259 35296 41260
rect 19616 40658 19936 40659
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 40593 19936 40594
rect 50336 40658 50656 40659
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 40593 50656 40594
rect 4256 39992 4576 39993
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 39927 4576 39928
rect 34976 39992 35296 39993
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 39927 35296 39928
rect 19616 39326 19936 39327
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 39261 19936 39262
rect 50336 39326 50656 39327
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 39261 50656 39262
rect 4256 38660 4576 38661
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 38595 4576 38596
rect 34976 38660 35296 38661
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 38595 35296 38596
rect 19616 37994 19936 37995
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 37929 19936 37930
rect 50336 37994 50656 37995
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 37929 50656 37930
rect 4256 37328 4576 37329
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 37263 4576 37264
rect 34976 37328 35296 37329
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 37263 35296 37264
rect 19616 36662 19936 36663
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 36597 19936 36598
rect 50336 36662 50656 36663
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 36597 50656 36598
rect 4256 35996 4576 35997
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 35931 4576 35932
rect 34976 35996 35296 35997
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 35931 35296 35932
rect 19616 35330 19936 35331
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 35265 19936 35266
rect 50336 35330 50656 35331
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 35265 50656 35266
rect 4256 34664 4576 34665
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 34599 4576 34600
rect 34976 34664 35296 34665
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 34599 35296 34600
rect 19616 33998 19936 33999
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 33933 19936 33934
rect 50336 33998 50656 33999
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 33933 50656 33934
rect 4256 33332 4576 33333
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 33267 4576 33268
rect 34976 33332 35296 33333
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 33267 35296 33268
rect 19616 32666 19936 32667
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 32601 19936 32602
rect 50336 32666 50656 32667
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 32601 50656 32602
rect 4256 32000 4576 32001
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 31935 4576 31936
rect 34976 32000 35296 32001
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 31935 35296 31936
rect 19616 31334 19936 31335
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 31269 19936 31270
rect 50336 31334 50656 31335
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 31269 50656 31270
rect 4256 30668 4576 30669
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 30603 4576 30604
rect 34976 30668 35296 30669
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 30603 35296 30604
rect 19616 30002 19936 30003
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 29937 19936 29938
rect 50336 30002 50656 30003
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 29937 50656 29938
rect 4256 29336 4576 29337
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 29271 4576 29272
rect 34976 29336 35296 29337
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 29271 35296 29272
rect 8122 28902 8128 28966
rect 8192 28964 8198 28966
rect 8367 28964 8433 28967
rect 8192 28962 8433 28964
rect 8192 28906 8372 28962
rect 8428 28906 8433 28962
rect 8192 28904 8433 28906
rect 8192 28902 8198 28904
rect 8367 28901 8433 28904
rect 19616 28670 19936 28671
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 28605 19936 28606
rect 50336 28670 50656 28671
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 28605 50656 28606
rect 4256 28004 4576 28005
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 27939 4576 27940
rect 34976 28004 35296 28005
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 27939 35296 27940
rect 19616 27338 19936 27339
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 27273 19936 27274
rect 50336 27338 50656 27339
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 27273 50656 27274
rect 4256 26672 4576 26673
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 26607 4576 26608
rect 34976 26672 35296 26673
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 26607 35296 26608
rect 8367 26154 8433 26155
rect 8314 26152 8320 26154
rect 8276 26092 8320 26152
rect 8384 26150 8433 26154
rect 8428 26094 8433 26150
rect 8314 26090 8320 26092
rect 8384 26090 8433 26094
rect 8367 26089 8433 26090
rect 19616 26006 19936 26007
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 25941 19936 25942
rect 50336 26006 50656 26007
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 25941 50656 25942
rect 4256 25340 4576 25341
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 25275 4576 25276
rect 34976 25340 35296 25341
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 25275 35296 25276
rect 7215 24968 7281 24971
rect 8223 24968 8289 24971
rect 7215 24966 8289 24968
rect 7215 24910 7220 24966
rect 7276 24910 8228 24966
rect 8284 24910 8289 24966
rect 7215 24908 8289 24910
rect 7215 24905 7281 24908
rect 8223 24905 8289 24908
rect 19616 24674 19936 24675
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 24609 19936 24610
rect 50336 24674 50656 24675
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 24609 50656 24610
rect 4256 24008 4576 24009
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 23943 4576 23944
rect 34976 24008 35296 24009
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 23943 35296 23944
rect 19616 23342 19936 23343
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 23277 19936 23278
rect 50336 23342 50656 23343
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 23277 50656 23278
rect 4256 22676 4576 22677
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 22611 4576 22612
rect 34976 22676 35296 22677
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 22611 35296 22612
rect 19616 22010 19936 22011
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 21945 19936 21946
rect 50336 22010 50656 22011
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 21945 50656 21946
rect 4256 21344 4576 21345
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 21279 4576 21280
rect 34976 21344 35296 21345
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 21279 35296 21280
rect 19616 20678 19936 20679
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 20613 19936 20614
rect 50336 20678 50656 20679
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 20613 50656 20614
rect 4256 20012 4576 20013
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 19947 4576 19948
rect 34976 20012 35296 20013
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 19947 35296 19948
rect 19616 19346 19936 19347
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 19281 19936 19282
rect 50336 19346 50656 19347
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 19281 50656 19282
rect 4256 18680 4576 18681
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 18615 4576 18616
rect 34976 18680 35296 18681
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 18615 35296 18616
rect 19616 18014 19936 18015
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 17949 19936 17950
rect 50336 18014 50656 18015
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 17949 50656 17950
rect 4256 17348 4576 17349
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 17283 4576 17284
rect 34976 17348 35296 17349
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 17283 35296 17284
rect 7407 17272 7473 17275
rect 9039 17272 9105 17275
rect 7407 17270 9105 17272
rect 7407 17214 7412 17270
rect 7468 17214 9044 17270
rect 9100 17214 9105 17270
rect 7407 17212 9105 17214
rect 7407 17209 7473 17212
rect 9039 17209 9105 17212
rect 19616 16682 19936 16683
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 16617 19936 16618
rect 50336 16682 50656 16683
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 16617 50656 16618
rect 4256 16016 4576 16017
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 15951 4576 15952
rect 34976 16016 35296 16017
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 15951 35296 15952
rect 19616 15350 19936 15351
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 15285 19936 15286
rect 50336 15350 50656 15351
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 15285 50656 15286
rect 4256 14684 4576 14685
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 14619 4576 14620
rect 34976 14684 35296 14685
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 14619 35296 14620
rect 19616 14018 19936 14019
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 13953 19936 13954
rect 50336 14018 50656 14019
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 13953 50656 13954
rect 7791 13424 7857 13427
rect 7983 13424 8049 13427
rect 7791 13422 8049 13424
rect 7791 13366 7796 13422
rect 7852 13366 7988 13422
rect 8044 13366 8049 13422
rect 7791 13364 8049 13366
rect 7791 13361 7857 13364
rect 7983 13361 8049 13364
rect 4256 13352 4576 13353
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 13287 4576 13288
rect 34976 13352 35296 13353
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 13287 35296 13288
rect 19616 12686 19936 12687
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 12621 19936 12622
rect 50336 12686 50656 12687
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 12621 50656 12622
rect 4256 12020 4576 12021
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 11955 4576 11956
rect 34976 12020 35296 12021
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 11955 35296 11956
rect 19616 11354 19936 11355
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 11289 19936 11290
rect 50336 11354 50656 11355
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 11289 50656 11290
rect 4256 10688 4576 10689
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 10623 4576 10624
rect 34976 10688 35296 10689
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 10623 35296 10624
rect 19616 10022 19936 10023
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 9957 19936 9958
rect 50336 10022 50656 10023
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 9957 50656 9958
rect 8367 9724 8433 9727
rect 8367 9722 8574 9724
rect 8367 9666 8372 9722
rect 8428 9666 8574 9722
rect 8367 9664 8574 9666
rect 8367 9661 8433 9664
rect 4256 9356 4576 9357
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 9291 4576 9292
rect 8514 8987 8574 9664
rect 34976 9356 35296 9357
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 9291 35296 9292
rect 8655 9132 8721 9135
rect 10042 9132 10048 9134
rect 8655 9130 10048 9132
rect 8655 9074 8660 9130
rect 8716 9074 10048 9130
rect 8655 9072 10048 9074
rect 8655 9069 8721 9072
rect 10042 9070 10048 9072
rect 10112 9070 10118 9134
rect 8514 8982 8625 8987
rect 8514 8926 8564 8982
rect 8620 8926 8625 8982
rect 8514 8924 8625 8926
rect 8559 8921 8625 8924
rect 8751 8984 8817 8987
rect 9039 8984 9105 8987
rect 8751 8982 9105 8984
rect 8751 8926 8756 8982
rect 8812 8926 9044 8982
rect 9100 8926 9105 8982
rect 8751 8924 9105 8926
rect 8751 8921 8817 8924
rect 9039 8921 9105 8924
rect 10863 8836 10929 8839
rect 16431 8836 16497 8839
rect 10863 8834 16497 8836
rect 10863 8778 10868 8834
rect 10924 8778 16436 8834
rect 16492 8778 16497 8834
rect 10863 8776 16497 8778
rect 10863 8773 10929 8776
rect 16431 8773 16497 8776
rect 11055 8688 11121 8691
rect 16335 8688 16401 8691
rect 11055 8686 16401 8688
rect 11055 8630 11060 8686
rect 11116 8630 16340 8686
rect 16396 8630 16401 8686
rect 11055 8628 16401 8630
rect 11055 8625 11121 8628
rect 16335 8625 16401 8628
rect 19616 8690 19936 8691
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 8625 19936 8626
rect 50336 8690 50656 8691
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 8625 50656 8626
rect 7503 8540 7569 8543
rect 7887 8540 7953 8543
rect 12975 8540 13041 8543
rect 7503 8538 7614 8540
rect 7503 8482 7508 8538
rect 7564 8482 7614 8538
rect 7503 8477 7614 8482
rect 7887 8538 13041 8540
rect 7887 8482 7892 8538
rect 7948 8482 12980 8538
rect 13036 8482 13041 8538
rect 7887 8480 13041 8482
rect 7887 8477 7953 8480
rect 12975 8477 13041 8480
rect 13647 8540 13713 8543
rect 52431 8540 52497 8543
rect 13647 8538 52497 8540
rect 13647 8482 13652 8538
rect 13708 8482 52436 8538
rect 52492 8482 52497 8538
rect 13647 8480 52497 8482
rect 13647 8477 13713 8480
rect 52431 8477 52497 8480
rect 7554 8392 7614 8477
rect 7983 8392 8049 8395
rect 7554 8390 8049 8392
rect 7554 8334 7988 8390
rect 8044 8334 8049 8390
rect 7554 8332 8049 8334
rect 7983 8329 8049 8332
rect 12399 8392 12465 8395
rect 52911 8392 52977 8395
rect 12399 8390 52977 8392
rect 12399 8334 12404 8390
rect 12460 8334 52916 8390
rect 52972 8334 52977 8390
rect 12399 8332 52977 8334
rect 12399 8329 12465 8332
rect 52911 8329 52977 8332
rect 2223 8244 2289 8247
rect 8559 8244 8625 8247
rect 40335 8244 40401 8247
rect 2223 8242 7998 8244
rect 2223 8186 2228 8242
rect 2284 8186 7998 8242
rect 2223 8184 7998 8186
rect 2223 8181 2289 8184
rect 7938 8096 7998 8184
rect 8559 8242 40401 8244
rect 8559 8186 8564 8242
rect 8620 8186 40340 8242
rect 40396 8186 40401 8242
rect 8559 8184 40401 8186
rect 8559 8181 8625 8184
rect 40335 8181 40401 8184
rect 46095 8244 46161 8247
rect 46479 8244 46545 8247
rect 46095 8242 46545 8244
rect 46095 8186 46100 8242
rect 46156 8186 46484 8242
rect 46540 8186 46545 8242
rect 46095 8184 46545 8186
rect 46095 8181 46161 8184
rect 46479 8181 46545 8184
rect 30831 8096 30897 8099
rect 7938 8094 30897 8096
rect 7938 8038 30836 8094
rect 30892 8038 30897 8094
rect 7938 8036 30897 8038
rect 30831 8033 30897 8036
rect 44175 8096 44241 8099
rect 47919 8096 47985 8099
rect 44175 8094 47985 8096
rect 44175 8038 44180 8094
rect 44236 8038 47924 8094
rect 47980 8038 47985 8094
rect 44175 8036 47985 8038
rect 44175 8033 44241 8036
rect 47919 8033 47985 8036
rect 4256 8024 4576 8025
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 7959 4576 7960
rect 34976 8024 35296 8025
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 7959 35296 7960
rect 8559 7948 8625 7951
rect 9039 7948 9105 7951
rect 8559 7946 9105 7948
rect 8559 7890 8564 7946
rect 8620 7890 9044 7946
rect 9100 7890 9105 7946
rect 8559 7888 9105 7890
rect 8559 7885 8625 7888
rect 9039 7885 9105 7888
rect 9423 7948 9489 7951
rect 28047 7948 28113 7951
rect 9423 7946 28113 7948
rect 9423 7890 9428 7946
rect 9484 7890 28052 7946
rect 28108 7890 28113 7946
rect 9423 7888 28113 7890
rect 9423 7885 9489 7888
rect 28047 7885 28113 7888
rect 38127 7948 38193 7951
rect 50031 7948 50097 7951
rect 38127 7946 50097 7948
rect 38127 7890 38132 7946
rect 38188 7890 50036 7946
rect 50092 7890 50097 7946
rect 38127 7888 50097 7890
rect 38127 7885 38193 7888
rect 50031 7885 50097 7888
rect 7599 7800 7665 7803
rect 8751 7800 8817 7803
rect 7599 7798 8817 7800
rect 7599 7742 7604 7798
rect 7660 7742 8756 7798
rect 8812 7742 8817 7798
rect 7599 7740 8817 7742
rect 7599 7737 7665 7740
rect 8751 7737 8817 7740
rect 10191 7800 10257 7803
rect 56367 7800 56433 7803
rect 10191 7798 56433 7800
rect 10191 7742 10196 7798
rect 10252 7742 56372 7798
rect 56428 7742 56433 7798
rect 10191 7740 56433 7742
rect 10191 7737 10257 7740
rect 56367 7737 56433 7740
rect 2511 7652 2577 7655
rect 38127 7652 38193 7655
rect 2511 7650 38193 7652
rect 2511 7594 2516 7650
rect 2572 7594 38132 7650
rect 38188 7594 38193 7650
rect 2511 7592 38193 7594
rect 2511 7589 2577 7592
rect 38127 7589 38193 7592
rect 8463 7504 8529 7507
rect 8751 7504 8817 7507
rect 9903 7506 9969 7507
rect 9850 7504 9856 7506
rect 8463 7502 8817 7504
rect 8463 7446 8468 7502
rect 8524 7446 8756 7502
rect 8812 7446 8817 7502
rect 8463 7444 8817 7446
rect 9812 7444 9856 7504
rect 9920 7502 9969 7506
rect 13935 7504 14001 7507
rect 52143 7504 52209 7507
rect 9964 7446 9969 7502
rect 8463 7441 8529 7444
rect 8751 7441 8817 7444
rect 9850 7442 9856 7444
rect 9920 7442 9969 7446
rect 9903 7441 9969 7442
rect 10050 7444 13758 7504
rect 6735 7356 6801 7359
rect 10050 7356 10110 7444
rect 6735 7354 10110 7356
rect 6735 7298 6740 7354
rect 6796 7298 10110 7354
rect 6735 7296 10110 7298
rect 12783 7356 12849 7359
rect 13263 7356 13329 7359
rect 12783 7354 13329 7356
rect 12783 7298 12788 7354
rect 12844 7298 13268 7354
rect 13324 7298 13329 7354
rect 12783 7296 13329 7298
rect 13698 7356 13758 7444
rect 13935 7502 52209 7504
rect 13935 7446 13940 7502
rect 13996 7446 52148 7502
rect 52204 7446 52209 7502
rect 13935 7444 52209 7446
rect 13935 7441 14001 7444
rect 52143 7441 52209 7444
rect 18927 7356 18993 7359
rect 13698 7354 18993 7356
rect 13698 7298 18932 7354
rect 18988 7298 18993 7354
rect 13698 7296 18993 7298
rect 6735 7293 6801 7296
rect 12783 7293 12849 7296
rect 13263 7293 13329 7296
rect 18927 7293 18993 7296
rect 19616 7358 19936 7359
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 7293 19936 7294
rect 20463 7356 20529 7359
rect 23151 7356 23217 7359
rect 20463 7354 23217 7356
rect 20463 7298 20468 7354
rect 20524 7298 23156 7354
rect 23212 7298 23217 7354
rect 20463 7296 23217 7298
rect 20463 7293 20529 7296
rect 23151 7293 23217 7296
rect 23823 7356 23889 7359
rect 27279 7356 27345 7359
rect 23823 7354 27345 7356
rect 23823 7298 23828 7354
rect 23884 7298 27284 7354
rect 27340 7298 27345 7354
rect 23823 7296 27345 7298
rect 23823 7293 23889 7296
rect 27279 7293 27345 7296
rect 28047 7356 28113 7359
rect 39375 7356 39441 7359
rect 28047 7354 39441 7356
rect 28047 7298 28052 7354
rect 28108 7298 39380 7354
rect 39436 7298 39441 7354
rect 28047 7296 39441 7298
rect 28047 7293 28113 7296
rect 39375 7293 39441 7296
rect 50336 7358 50656 7359
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 7293 50656 7294
rect 7311 7208 7377 7211
rect 7887 7208 7953 7211
rect 7311 7206 7953 7208
rect 7311 7150 7316 7206
rect 7372 7150 7892 7206
rect 7948 7150 7953 7206
rect 7311 7148 7953 7150
rect 7311 7145 7377 7148
rect 7887 7145 7953 7148
rect 12207 7208 12273 7211
rect 52719 7208 52785 7211
rect 12207 7206 52785 7208
rect 12207 7150 12212 7206
rect 12268 7150 52724 7206
rect 52780 7150 52785 7206
rect 12207 7148 52785 7150
rect 12207 7145 12273 7148
rect 52719 7145 52785 7148
rect 5391 7060 5457 7063
rect 46287 7060 46353 7063
rect 5391 7058 46353 7060
rect 5391 7002 5396 7058
rect 5452 7002 46292 7058
rect 46348 7002 46353 7058
rect 5391 7000 46353 7002
rect 5391 6997 5457 7000
rect 46287 6997 46353 7000
rect 4527 6912 4593 6915
rect 9999 6912 10065 6915
rect 4527 6910 10065 6912
rect 4527 6854 4532 6910
rect 4588 6854 10004 6910
rect 10060 6854 10065 6910
rect 4527 6852 10065 6854
rect 4527 6849 4593 6852
rect 9999 6849 10065 6852
rect 10575 6912 10641 6915
rect 53583 6912 53649 6915
rect 10575 6910 53649 6912
rect 10575 6854 10580 6910
rect 10636 6854 53588 6910
rect 53644 6854 53649 6910
rect 10575 6852 53649 6854
rect 10575 6849 10641 6852
rect 53583 6849 53649 6852
rect 10863 6764 10929 6767
rect 12975 6764 13041 6767
rect 10863 6762 13041 6764
rect 10863 6706 10868 6762
rect 10924 6706 12980 6762
rect 13036 6706 13041 6762
rect 10863 6704 13041 6706
rect 10863 6701 10929 6704
rect 12975 6701 13041 6704
rect 29050 6702 29056 6766
rect 29120 6764 29126 6766
rect 33039 6764 33105 6767
rect 29120 6762 33105 6764
rect 29120 6706 33044 6762
rect 33100 6706 33105 6762
rect 29120 6704 33105 6706
rect 29120 6702 29126 6704
rect 33039 6701 33105 6704
rect 33807 6764 33873 6767
rect 34575 6764 34641 6767
rect 33807 6762 34641 6764
rect 33807 6706 33812 6762
rect 33868 6706 34580 6762
rect 34636 6706 34641 6762
rect 33807 6704 34641 6706
rect 33807 6701 33873 6704
rect 34575 6701 34641 6704
rect 35439 6764 35505 6767
rect 39279 6764 39345 6767
rect 35439 6762 39345 6764
rect 35439 6706 35444 6762
rect 35500 6706 39284 6762
rect 39340 6706 39345 6762
rect 35439 6704 39345 6706
rect 35439 6701 35505 6704
rect 39279 6701 39345 6704
rect 42351 6764 42417 6767
rect 48495 6764 48561 6767
rect 42351 6762 48561 6764
rect 42351 6706 42356 6762
rect 42412 6706 48500 6762
rect 48556 6706 48561 6762
rect 42351 6704 48561 6706
rect 42351 6701 42417 6704
rect 48495 6701 48561 6704
rect 4256 6692 4576 6693
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 6627 4576 6628
rect 34976 6692 35296 6693
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 6627 35296 6628
rect 18351 6616 18417 6619
rect 23631 6616 23697 6619
rect 28282 6616 28288 6618
rect 18351 6614 23070 6616
rect 18351 6558 18356 6614
rect 18412 6558 23070 6614
rect 18351 6556 23070 6558
rect 18351 6553 18417 6556
rect 19599 6468 19665 6471
rect 22671 6468 22737 6471
rect 19599 6466 22737 6468
rect 19599 6410 19604 6466
rect 19660 6410 22676 6466
rect 22732 6410 22737 6466
rect 19599 6408 22737 6410
rect 23010 6468 23070 6556
rect 23631 6614 28288 6616
rect 23631 6558 23636 6614
rect 23692 6558 28288 6614
rect 23631 6556 28288 6558
rect 23631 6553 23697 6556
rect 28282 6554 28288 6556
rect 28352 6554 28358 6618
rect 28431 6616 28497 6619
rect 32847 6616 32913 6619
rect 28431 6614 32913 6616
rect 28431 6558 28436 6614
rect 28492 6558 32852 6614
rect 32908 6558 32913 6614
rect 28431 6556 32913 6558
rect 28431 6553 28497 6556
rect 32847 6553 32913 6556
rect 33135 6616 33201 6619
rect 33135 6614 34878 6616
rect 33135 6558 33140 6614
rect 33196 6558 34878 6614
rect 33135 6556 34878 6558
rect 33135 6553 33201 6556
rect 34671 6468 34737 6471
rect 23010 6466 34737 6468
rect 23010 6410 34676 6466
rect 34732 6410 34737 6466
rect 23010 6408 34737 6410
rect 34818 6468 34878 6556
rect 41871 6468 41937 6471
rect 34818 6466 41937 6468
rect 34818 6410 41876 6466
rect 41932 6410 41937 6466
rect 34818 6408 41937 6410
rect 19599 6405 19665 6408
rect 22671 6405 22737 6408
rect 34671 6405 34737 6408
rect 41871 6405 41937 6408
rect 24015 6320 24081 6323
rect 32751 6320 32817 6323
rect 24015 6318 32817 6320
rect 24015 6262 24020 6318
rect 24076 6262 32756 6318
rect 32812 6262 32817 6318
rect 24015 6260 32817 6262
rect 24015 6257 24081 6260
rect 32751 6257 32817 6260
rect 33039 6320 33105 6323
rect 43695 6320 43761 6323
rect 33039 6318 43761 6320
rect 33039 6262 33044 6318
rect 33100 6262 43700 6318
rect 43756 6262 43761 6318
rect 33039 6260 43761 6262
rect 33039 6257 33105 6260
rect 43695 6257 43761 6260
rect 17583 6172 17649 6175
rect 42351 6172 42417 6175
rect 17583 6170 42417 6172
rect 17583 6114 17588 6170
rect 17644 6114 42356 6170
rect 42412 6114 42417 6170
rect 17583 6112 42417 6114
rect 17583 6109 17649 6112
rect 42351 6109 42417 6112
rect 19616 6026 19936 6027
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 5961 19936 5962
rect 21327 6024 21393 6027
rect 46383 6024 46449 6027
rect 21327 6022 46449 6024
rect 21327 5966 21332 6022
rect 21388 5966 46388 6022
rect 46444 5966 46449 6022
rect 21327 5964 46449 5966
rect 21327 5961 21393 5964
rect 46383 5961 46449 5964
rect 50336 6026 50656 6027
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 5961 50656 5962
rect 17775 5876 17841 5879
rect 40719 5876 40785 5879
rect 17775 5874 40785 5876
rect 17775 5818 17780 5874
rect 17836 5818 40724 5874
rect 40780 5818 40785 5874
rect 17775 5816 40785 5818
rect 17775 5813 17841 5816
rect 40719 5813 40785 5816
rect 22671 5728 22737 5731
rect 30063 5728 30129 5731
rect 22671 5726 30129 5728
rect 22671 5670 22676 5726
rect 22732 5670 30068 5726
rect 30124 5670 30129 5726
rect 22671 5668 30129 5670
rect 22671 5665 22737 5668
rect 30063 5665 30129 5668
rect 4256 5360 4576 5361
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 5295 4576 5296
rect 34976 5360 35296 5361
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 5295 35296 5296
rect 56559 4988 56625 4991
rect 56514 4986 56625 4988
rect 56514 4930 56564 4986
rect 56620 4930 56625 4986
rect 56514 4925 56625 4930
rect 19616 4694 19936 4695
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 4629 19936 4630
rect 50336 4694 50656 4695
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 56514 4692 56574 4925
rect 56655 4692 56721 4695
rect 56514 4690 56721 4692
rect 56514 4634 56660 4690
rect 56716 4634 56721 4690
rect 56514 4632 56721 4634
rect 50336 4629 50656 4630
rect 56655 4629 56721 4632
rect 9711 4544 9777 4547
rect 8130 4542 9777 4544
rect 8130 4486 9716 4542
rect 9772 4486 9777 4542
rect 8130 4484 9777 4486
rect 8130 4399 8190 4484
rect 9711 4481 9777 4484
rect 8079 4394 8190 4399
rect 8079 4338 8084 4394
rect 8140 4338 8190 4394
rect 8079 4336 8190 4338
rect 8079 4333 8145 4336
rect 7983 4248 8049 4251
rect 19215 4248 19281 4251
rect 7983 4246 19281 4248
rect 7983 4190 7988 4246
rect 8044 4190 19220 4246
rect 19276 4190 19281 4246
rect 7983 4188 19281 4190
rect 7983 4185 8049 4188
rect 19215 4185 19281 4188
rect 4256 4028 4576 4029
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 3963 4576 3964
rect 34976 4028 35296 4029
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 3963 35296 3964
rect 9903 3954 9969 3955
rect 9850 3890 9856 3954
rect 9920 3952 9969 3954
rect 9920 3950 10012 3952
rect 9964 3894 10012 3950
rect 9920 3892 10012 3894
rect 9920 3890 9969 3892
rect 9903 3889 9969 3890
rect 8559 3804 8625 3807
rect 13743 3804 13809 3807
rect 34287 3804 34353 3807
rect 8559 3802 13809 3804
rect 8559 3746 8564 3802
rect 8620 3746 13748 3802
rect 13804 3746 13809 3802
rect 8559 3744 13809 3746
rect 8559 3741 8625 3744
rect 13743 3741 13809 3744
rect 34050 3802 34353 3804
rect 34050 3746 34292 3802
rect 34348 3746 34353 3802
rect 34050 3744 34353 3746
rect 10042 3594 10048 3658
rect 10112 3656 10118 3658
rect 10112 3596 12990 3656
rect 10112 3594 10118 3596
rect 12930 3508 12990 3596
rect 20847 3508 20913 3511
rect 12930 3506 20913 3508
rect 12930 3450 20852 3506
rect 20908 3450 20913 3506
rect 12930 3448 20913 3450
rect 20847 3445 20913 3448
rect 19616 3362 19936 3363
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 19616 3297 19936 3298
rect 33711 3360 33777 3363
rect 34050 3360 34110 3744
rect 34287 3741 34353 3744
rect 33711 3358 34110 3360
rect 33711 3302 33716 3358
rect 33772 3302 34110 3358
rect 33711 3300 34110 3302
rect 50336 3362 50656 3363
rect 33711 3297 33777 3300
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 50336 3297 50656 3298
rect 8314 3150 8320 3214
rect 8384 3212 8390 3214
rect 21135 3212 21201 3215
rect 8384 3210 21201 3212
rect 8384 3154 21140 3210
rect 21196 3154 21201 3210
rect 8384 3152 21201 3154
rect 8384 3150 8390 3152
rect 21135 3149 21201 3152
rect 7354 3002 7360 3066
rect 7424 3064 7430 3066
rect 56367 3064 56433 3067
rect 7424 3062 56433 3064
rect 7424 3006 56372 3062
rect 56428 3006 56433 3062
rect 7424 3004 56433 3006
rect 7424 3002 7430 3004
rect 56367 3001 56433 3004
rect 8122 2854 8128 2918
rect 8192 2916 8198 2918
rect 21135 2916 21201 2919
rect 8192 2914 21201 2916
rect 8192 2858 21140 2914
rect 21196 2858 21201 2914
rect 8192 2856 21201 2858
rect 8192 2854 8198 2856
rect 21135 2853 21201 2856
rect 4256 2696 4576 2697
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4256 2631 4576 2632
rect 34976 2696 35296 2697
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 34976 2631 35296 2632
<< via3 >>
rect 4264 57304 4328 57308
rect 4264 57248 4268 57304
rect 4268 57248 4324 57304
rect 4324 57248 4328 57304
rect 4264 57244 4328 57248
rect 4344 57304 4408 57308
rect 4344 57248 4348 57304
rect 4348 57248 4404 57304
rect 4404 57248 4408 57304
rect 4344 57244 4408 57248
rect 4424 57304 4488 57308
rect 4424 57248 4428 57304
rect 4428 57248 4484 57304
rect 4484 57248 4488 57304
rect 4424 57244 4488 57248
rect 4504 57304 4568 57308
rect 4504 57248 4508 57304
rect 4508 57248 4564 57304
rect 4564 57248 4568 57304
rect 4504 57244 4568 57248
rect 34984 57304 35048 57308
rect 34984 57248 34988 57304
rect 34988 57248 35044 57304
rect 35044 57248 35048 57304
rect 34984 57244 35048 57248
rect 35064 57304 35128 57308
rect 35064 57248 35068 57304
rect 35068 57248 35124 57304
rect 35124 57248 35128 57304
rect 35064 57244 35128 57248
rect 35144 57304 35208 57308
rect 35144 57248 35148 57304
rect 35148 57248 35204 57304
rect 35204 57248 35208 57304
rect 35144 57244 35208 57248
rect 35224 57304 35288 57308
rect 35224 57248 35228 57304
rect 35228 57248 35284 57304
rect 35284 57248 35288 57304
rect 35224 57244 35288 57248
rect 19624 56638 19688 56642
rect 19624 56582 19628 56638
rect 19628 56582 19684 56638
rect 19684 56582 19688 56638
rect 19624 56578 19688 56582
rect 19704 56638 19768 56642
rect 19704 56582 19708 56638
rect 19708 56582 19764 56638
rect 19764 56582 19768 56638
rect 19704 56578 19768 56582
rect 19784 56638 19848 56642
rect 19784 56582 19788 56638
rect 19788 56582 19844 56638
rect 19844 56582 19848 56638
rect 19784 56578 19848 56582
rect 19864 56638 19928 56642
rect 19864 56582 19868 56638
rect 19868 56582 19924 56638
rect 19924 56582 19928 56638
rect 19864 56578 19928 56582
rect 50344 56638 50408 56642
rect 50344 56582 50348 56638
rect 50348 56582 50404 56638
rect 50404 56582 50408 56638
rect 50344 56578 50408 56582
rect 50424 56638 50488 56642
rect 50424 56582 50428 56638
rect 50428 56582 50484 56638
rect 50484 56582 50488 56638
rect 50424 56578 50488 56582
rect 50504 56638 50568 56642
rect 50504 56582 50508 56638
rect 50508 56582 50564 56638
rect 50564 56582 50568 56638
rect 50504 56578 50568 56582
rect 50584 56638 50648 56642
rect 50584 56582 50588 56638
rect 50588 56582 50644 56638
rect 50644 56582 50648 56638
rect 50584 56578 50648 56582
rect 7360 56134 7424 56198
rect 4264 55972 4328 55976
rect 4264 55916 4268 55972
rect 4268 55916 4324 55972
rect 4324 55916 4328 55972
rect 4264 55912 4328 55916
rect 4344 55972 4408 55976
rect 4344 55916 4348 55972
rect 4348 55916 4404 55972
rect 4404 55916 4408 55972
rect 4344 55912 4408 55916
rect 4424 55972 4488 55976
rect 4424 55916 4428 55972
rect 4428 55916 4484 55972
rect 4484 55916 4488 55972
rect 4424 55912 4488 55916
rect 4504 55972 4568 55976
rect 4504 55916 4508 55972
rect 4508 55916 4564 55972
rect 4564 55916 4568 55972
rect 4504 55912 4568 55916
rect 34984 55972 35048 55976
rect 34984 55916 34988 55972
rect 34988 55916 35044 55972
rect 35044 55916 35048 55972
rect 34984 55912 35048 55916
rect 35064 55972 35128 55976
rect 35064 55916 35068 55972
rect 35068 55916 35124 55972
rect 35124 55916 35128 55972
rect 35064 55912 35128 55916
rect 35144 55972 35208 55976
rect 35144 55916 35148 55972
rect 35148 55916 35204 55972
rect 35204 55916 35208 55972
rect 35144 55912 35208 55916
rect 35224 55972 35288 55976
rect 35224 55916 35228 55972
rect 35228 55916 35284 55972
rect 35284 55916 35288 55972
rect 35224 55912 35288 55916
rect 19624 55306 19688 55310
rect 19624 55250 19628 55306
rect 19628 55250 19684 55306
rect 19684 55250 19688 55306
rect 19624 55246 19688 55250
rect 19704 55306 19768 55310
rect 19704 55250 19708 55306
rect 19708 55250 19764 55306
rect 19764 55250 19768 55306
rect 19704 55246 19768 55250
rect 19784 55306 19848 55310
rect 19784 55250 19788 55306
rect 19788 55250 19844 55306
rect 19844 55250 19848 55306
rect 19784 55246 19848 55250
rect 19864 55306 19928 55310
rect 19864 55250 19868 55306
rect 19868 55250 19924 55306
rect 19924 55250 19928 55306
rect 19864 55246 19928 55250
rect 50344 55306 50408 55310
rect 50344 55250 50348 55306
rect 50348 55250 50404 55306
rect 50404 55250 50408 55306
rect 50344 55246 50408 55250
rect 50424 55306 50488 55310
rect 50424 55250 50428 55306
rect 50428 55250 50484 55306
rect 50484 55250 50488 55306
rect 50424 55246 50488 55250
rect 50504 55306 50568 55310
rect 50504 55250 50508 55306
rect 50508 55250 50564 55306
rect 50564 55250 50568 55306
rect 50504 55246 50568 55250
rect 50584 55306 50648 55310
rect 50584 55250 50588 55306
rect 50588 55250 50644 55306
rect 50644 55250 50648 55306
rect 50584 55246 50648 55250
rect 4264 54640 4328 54644
rect 4264 54584 4268 54640
rect 4268 54584 4324 54640
rect 4324 54584 4328 54640
rect 4264 54580 4328 54584
rect 4344 54640 4408 54644
rect 4344 54584 4348 54640
rect 4348 54584 4404 54640
rect 4404 54584 4408 54640
rect 4344 54580 4408 54584
rect 4424 54640 4488 54644
rect 4424 54584 4428 54640
rect 4428 54584 4484 54640
rect 4484 54584 4488 54640
rect 4424 54580 4488 54584
rect 4504 54640 4568 54644
rect 4504 54584 4508 54640
rect 4508 54584 4564 54640
rect 4564 54584 4568 54640
rect 4504 54580 4568 54584
rect 34984 54640 35048 54644
rect 34984 54584 34988 54640
rect 34988 54584 35044 54640
rect 35044 54584 35048 54640
rect 34984 54580 35048 54584
rect 35064 54640 35128 54644
rect 35064 54584 35068 54640
rect 35068 54584 35124 54640
rect 35124 54584 35128 54640
rect 35064 54580 35128 54584
rect 35144 54640 35208 54644
rect 35144 54584 35148 54640
rect 35148 54584 35204 54640
rect 35204 54584 35208 54640
rect 35144 54580 35208 54584
rect 35224 54640 35288 54644
rect 35224 54584 35228 54640
rect 35228 54584 35284 54640
rect 35284 54584 35288 54640
rect 35224 54580 35288 54584
rect 19624 53974 19688 53978
rect 19624 53918 19628 53974
rect 19628 53918 19684 53974
rect 19684 53918 19688 53974
rect 19624 53914 19688 53918
rect 19704 53974 19768 53978
rect 19704 53918 19708 53974
rect 19708 53918 19764 53974
rect 19764 53918 19768 53974
rect 19704 53914 19768 53918
rect 19784 53974 19848 53978
rect 19784 53918 19788 53974
rect 19788 53918 19844 53974
rect 19844 53918 19848 53974
rect 19784 53914 19848 53918
rect 19864 53974 19928 53978
rect 19864 53918 19868 53974
rect 19868 53918 19924 53974
rect 19924 53918 19928 53974
rect 19864 53914 19928 53918
rect 50344 53974 50408 53978
rect 50344 53918 50348 53974
rect 50348 53918 50404 53974
rect 50404 53918 50408 53974
rect 50344 53914 50408 53918
rect 50424 53974 50488 53978
rect 50424 53918 50428 53974
rect 50428 53918 50484 53974
rect 50484 53918 50488 53974
rect 50424 53914 50488 53918
rect 50504 53974 50568 53978
rect 50504 53918 50508 53974
rect 50508 53918 50564 53974
rect 50564 53918 50568 53974
rect 50504 53914 50568 53918
rect 50584 53974 50648 53978
rect 50584 53918 50588 53974
rect 50588 53918 50644 53974
rect 50644 53918 50648 53974
rect 50584 53914 50648 53918
rect 4264 53308 4328 53312
rect 4264 53252 4268 53308
rect 4268 53252 4324 53308
rect 4324 53252 4328 53308
rect 4264 53248 4328 53252
rect 4344 53308 4408 53312
rect 4344 53252 4348 53308
rect 4348 53252 4404 53308
rect 4404 53252 4408 53308
rect 4344 53248 4408 53252
rect 4424 53308 4488 53312
rect 4424 53252 4428 53308
rect 4428 53252 4484 53308
rect 4484 53252 4488 53308
rect 4424 53248 4488 53252
rect 4504 53308 4568 53312
rect 4504 53252 4508 53308
rect 4508 53252 4564 53308
rect 4564 53252 4568 53308
rect 4504 53248 4568 53252
rect 34984 53308 35048 53312
rect 34984 53252 34988 53308
rect 34988 53252 35044 53308
rect 35044 53252 35048 53308
rect 34984 53248 35048 53252
rect 35064 53308 35128 53312
rect 35064 53252 35068 53308
rect 35068 53252 35124 53308
rect 35124 53252 35128 53308
rect 35064 53248 35128 53252
rect 35144 53308 35208 53312
rect 35144 53252 35148 53308
rect 35148 53252 35204 53308
rect 35204 53252 35208 53308
rect 35144 53248 35208 53252
rect 35224 53308 35288 53312
rect 35224 53252 35228 53308
rect 35228 53252 35284 53308
rect 35284 53252 35288 53308
rect 35224 53248 35288 53252
rect 19624 52642 19688 52646
rect 19624 52586 19628 52642
rect 19628 52586 19684 52642
rect 19684 52586 19688 52642
rect 19624 52582 19688 52586
rect 19704 52642 19768 52646
rect 19704 52586 19708 52642
rect 19708 52586 19764 52642
rect 19764 52586 19768 52642
rect 19704 52582 19768 52586
rect 19784 52642 19848 52646
rect 19784 52586 19788 52642
rect 19788 52586 19844 52642
rect 19844 52586 19848 52642
rect 19784 52582 19848 52586
rect 19864 52642 19928 52646
rect 19864 52586 19868 52642
rect 19868 52586 19924 52642
rect 19924 52586 19928 52642
rect 19864 52582 19928 52586
rect 50344 52642 50408 52646
rect 50344 52586 50348 52642
rect 50348 52586 50404 52642
rect 50404 52586 50408 52642
rect 50344 52582 50408 52586
rect 50424 52642 50488 52646
rect 50424 52586 50428 52642
rect 50428 52586 50484 52642
rect 50484 52586 50488 52642
rect 50424 52582 50488 52586
rect 50504 52642 50568 52646
rect 50504 52586 50508 52642
rect 50508 52586 50564 52642
rect 50564 52586 50568 52642
rect 50504 52582 50568 52586
rect 50584 52642 50648 52646
rect 50584 52586 50588 52642
rect 50588 52586 50644 52642
rect 50644 52586 50648 52642
rect 50584 52582 50648 52586
rect 4264 51976 4328 51980
rect 4264 51920 4268 51976
rect 4268 51920 4324 51976
rect 4324 51920 4328 51976
rect 4264 51916 4328 51920
rect 4344 51976 4408 51980
rect 4344 51920 4348 51976
rect 4348 51920 4404 51976
rect 4404 51920 4408 51976
rect 4344 51916 4408 51920
rect 4424 51976 4488 51980
rect 4424 51920 4428 51976
rect 4428 51920 4484 51976
rect 4484 51920 4488 51976
rect 4424 51916 4488 51920
rect 4504 51976 4568 51980
rect 4504 51920 4508 51976
rect 4508 51920 4564 51976
rect 4564 51920 4568 51976
rect 4504 51916 4568 51920
rect 34984 51976 35048 51980
rect 34984 51920 34988 51976
rect 34988 51920 35044 51976
rect 35044 51920 35048 51976
rect 34984 51916 35048 51920
rect 35064 51976 35128 51980
rect 35064 51920 35068 51976
rect 35068 51920 35124 51976
rect 35124 51920 35128 51976
rect 35064 51916 35128 51920
rect 35144 51976 35208 51980
rect 35144 51920 35148 51976
rect 35148 51920 35204 51976
rect 35204 51920 35208 51976
rect 35144 51916 35208 51920
rect 35224 51976 35288 51980
rect 35224 51920 35228 51976
rect 35228 51920 35284 51976
rect 35284 51920 35288 51976
rect 35224 51916 35288 51920
rect 19624 51310 19688 51314
rect 19624 51254 19628 51310
rect 19628 51254 19684 51310
rect 19684 51254 19688 51310
rect 19624 51250 19688 51254
rect 19704 51310 19768 51314
rect 19704 51254 19708 51310
rect 19708 51254 19764 51310
rect 19764 51254 19768 51310
rect 19704 51250 19768 51254
rect 19784 51310 19848 51314
rect 19784 51254 19788 51310
rect 19788 51254 19844 51310
rect 19844 51254 19848 51310
rect 19784 51250 19848 51254
rect 19864 51310 19928 51314
rect 19864 51254 19868 51310
rect 19868 51254 19924 51310
rect 19924 51254 19928 51310
rect 19864 51250 19928 51254
rect 50344 51310 50408 51314
rect 50344 51254 50348 51310
rect 50348 51254 50404 51310
rect 50404 51254 50408 51310
rect 50344 51250 50408 51254
rect 50424 51310 50488 51314
rect 50424 51254 50428 51310
rect 50428 51254 50484 51310
rect 50484 51254 50488 51310
rect 50424 51250 50488 51254
rect 50504 51310 50568 51314
rect 50504 51254 50508 51310
rect 50508 51254 50564 51310
rect 50564 51254 50568 51310
rect 50504 51250 50568 51254
rect 50584 51310 50648 51314
rect 50584 51254 50588 51310
rect 50588 51254 50644 51310
rect 50644 51254 50648 51310
rect 50584 51250 50648 51254
rect 4264 50644 4328 50648
rect 4264 50588 4268 50644
rect 4268 50588 4324 50644
rect 4324 50588 4328 50644
rect 4264 50584 4328 50588
rect 4344 50644 4408 50648
rect 4344 50588 4348 50644
rect 4348 50588 4404 50644
rect 4404 50588 4408 50644
rect 4344 50584 4408 50588
rect 4424 50644 4488 50648
rect 4424 50588 4428 50644
rect 4428 50588 4484 50644
rect 4484 50588 4488 50644
rect 4424 50584 4488 50588
rect 4504 50644 4568 50648
rect 4504 50588 4508 50644
rect 4508 50588 4564 50644
rect 4564 50588 4568 50644
rect 4504 50584 4568 50588
rect 34984 50644 35048 50648
rect 34984 50588 34988 50644
rect 34988 50588 35044 50644
rect 35044 50588 35048 50644
rect 34984 50584 35048 50588
rect 35064 50644 35128 50648
rect 35064 50588 35068 50644
rect 35068 50588 35124 50644
rect 35124 50588 35128 50644
rect 35064 50584 35128 50588
rect 35144 50644 35208 50648
rect 35144 50588 35148 50644
rect 35148 50588 35204 50644
rect 35204 50588 35208 50644
rect 35144 50584 35208 50588
rect 35224 50644 35288 50648
rect 35224 50588 35228 50644
rect 35228 50588 35284 50644
rect 35284 50588 35288 50644
rect 35224 50584 35288 50588
rect 19624 49978 19688 49982
rect 19624 49922 19628 49978
rect 19628 49922 19684 49978
rect 19684 49922 19688 49978
rect 19624 49918 19688 49922
rect 19704 49978 19768 49982
rect 19704 49922 19708 49978
rect 19708 49922 19764 49978
rect 19764 49922 19768 49978
rect 19704 49918 19768 49922
rect 19784 49978 19848 49982
rect 19784 49922 19788 49978
rect 19788 49922 19844 49978
rect 19844 49922 19848 49978
rect 19784 49918 19848 49922
rect 19864 49978 19928 49982
rect 19864 49922 19868 49978
rect 19868 49922 19924 49978
rect 19924 49922 19928 49978
rect 19864 49918 19928 49922
rect 50344 49978 50408 49982
rect 50344 49922 50348 49978
rect 50348 49922 50404 49978
rect 50404 49922 50408 49978
rect 50344 49918 50408 49922
rect 50424 49978 50488 49982
rect 50424 49922 50428 49978
rect 50428 49922 50484 49978
rect 50484 49922 50488 49978
rect 50424 49918 50488 49922
rect 50504 49978 50568 49982
rect 50504 49922 50508 49978
rect 50508 49922 50564 49978
rect 50564 49922 50568 49978
rect 50504 49918 50568 49922
rect 50584 49978 50648 49982
rect 50584 49922 50588 49978
rect 50588 49922 50644 49978
rect 50644 49922 50648 49978
rect 50584 49918 50648 49922
rect 4264 49312 4328 49316
rect 4264 49256 4268 49312
rect 4268 49256 4324 49312
rect 4324 49256 4328 49312
rect 4264 49252 4328 49256
rect 4344 49312 4408 49316
rect 4344 49256 4348 49312
rect 4348 49256 4404 49312
rect 4404 49256 4408 49312
rect 4344 49252 4408 49256
rect 4424 49312 4488 49316
rect 4424 49256 4428 49312
rect 4428 49256 4484 49312
rect 4484 49256 4488 49312
rect 4424 49252 4488 49256
rect 4504 49312 4568 49316
rect 4504 49256 4508 49312
rect 4508 49256 4564 49312
rect 4564 49256 4568 49312
rect 4504 49252 4568 49256
rect 34984 49312 35048 49316
rect 34984 49256 34988 49312
rect 34988 49256 35044 49312
rect 35044 49256 35048 49312
rect 34984 49252 35048 49256
rect 35064 49312 35128 49316
rect 35064 49256 35068 49312
rect 35068 49256 35124 49312
rect 35124 49256 35128 49312
rect 35064 49252 35128 49256
rect 35144 49312 35208 49316
rect 35144 49256 35148 49312
rect 35148 49256 35204 49312
rect 35204 49256 35208 49312
rect 35144 49252 35208 49256
rect 35224 49312 35288 49316
rect 35224 49256 35228 49312
rect 35228 49256 35284 49312
rect 35284 49256 35288 49312
rect 35224 49252 35288 49256
rect 19624 48646 19688 48650
rect 19624 48590 19628 48646
rect 19628 48590 19684 48646
rect 19684 48590 19688 48646
rect 19624 48586 19688 48590
rect 19704 48646 19768 48650
rect 19704 48590 19708 48646
rect 19708 48590 19764 48646
rect 19764 48590 19768 48646
rect 19704 48586 19768 48590
rect 19784 48646 19848 48650
rect 19784 48590 19788 48646
rect 19788 48590 19844 48646
rect 19844 48590 19848 48646
rect 19784 48586 19848 48590
rect 19864 48646 19928 48650
rect 19864 48590 19868 48646
rect 19868 48590 19924 48646
rect 19924 48590 19928 48646
rect 19864 48586 19928 48590
rect 50344 48646 50408 48650
rect 50344 48590 50348 48646
rect 50348 48590 50404 48646
rect 50404 48590 50408 48646
rect 50344 48586 50408 48590
rect 50424 48646 50488 48650
rect 50424 48590 50428 48646
rect 50428 48590 50484 48646
rect 50484 48590 50488 48646
rect 50424 48586 50488 48590
rect 50504 48646 50568 48650
rect 50504 48590 50508 48646
rect 50508 48590 50564 48646
rect 50564 48590 50568 48646
rect 50504 48586 50568 48590
rect 50584 48646 50648 48650
rect 50584 48590 50588 48646
rect 50588 48590 50644 48646
rect 50644 48590 50648 48646
rect 50584 48586 50648 48590
rect 4264 47980 4328 47984
rect 4264 47924 4268 47980
rect 4268 47924 4324 47980
rect 4324 47924 4328 47980
rect 4264 47920 4328 47924
rect 4344 47980 4408 47984
rect 4344 47924 4348 47980
rect 4348 47924 4404 47980
rect 4404 47924 4408 47980
rect 4344 47920 4408 47924
rect 4424 47980 4488 47984
rect 4424 47924 4428 47980
rect 4428 47924 4484 47980
rect 4484 47924 4488 47980
rect 4424 47920 4488 47924
rect 4504 47980 4568 47984
rect 4504 47924 4508 47980
rect 4508 47924 4564 47980
rect 4564 47924 4568 47980
rect 4504 47920 4568 47924
rect 34984 47980 35048 47984
rect 34984 47924 34988 47980
rect 34988 47924 35044 47980
rect 35044 47924 35048 47980
rect 34984 47920 35048 47924
rect 35064 47980 35128 47984
rect 35064 47924 35068 47980
rect 35068 47924 35124 47980
rect 35124 47924 35128 47980
rect 35064 47920 35128 47924
rect 35144 47980 35208 47984
rect 35144 47924 35148 47980
rect 35148 47924 35204 47980
rect 35204 47924 35208 47980
rect 35144 47920 35208 47924
rect 35224 47980 35288 47984
rect 35224 47924 35228 47980
rect 35228 47924 35284 47980
rect 35284 47924 35288 47980
rect 35224 47920 35288 47924
rect 19624 47314 19688 47318
rect 19624 47258 19628 47314
rect 19628 47258 19684 47314
rect 19684 47258 19688 47314
rect 19624 47254 19688 47258
rect 19704 47314 19768 47318
rect 19704 47258 19708 47314
rect 19708 47258 19764 47314
rect 19764 47258 19768 47314
rect 19704 47254 19768 47258
rect 19784 47314 19848 47318
rect 19784 47258 19788 47314
rect 19788 47258 19844 47314
rect 19844 47258 19848 47314
rect 19784 47254 19848 47258
rect 19864 47314 19928 47318
rect 19864 47258 19868 47314
rect 19868 47258 19924 47314
rect 19924 47258 19928 47314
rect 19864 47254 19928 47258
rect 50344 47314 50408 47318
rect 50344 47258 50348 47314
rect 50348 47258 50404 47314
rect 50404 47258 50408 47314
rect 50344 47254 50408 47258
rect 50424 47314 50488 47318
rect 50424 47258 50428 47314
rect 50428 47258 50484 47314
rect 50484 47258 50488 47314
rect 50424 47254 50488 47258
rect 50504 47314 50568 47318
rect 50504 47258 50508 47314
rect 50508 47258 50564 47314
rect 50564 47258 50568 47314
rect 50504 47254 50568 47258
rect 50584 47314 50648 47318
rect 50584 47258 50588 47314
rect 50588 47258 50644 47314
rect 50644 47258 50648 47314
rect 50584 47254 50648 47258
rect 4264 46648 4328 46652
rect 4264 46592 4268 46648
rect 4268 46592 4324 46648
rect 4324 46592 4328 46648
rect 4264 46588 4328 46592
rect 4344 46648 4408 46652
rect 4344 46592 4348 46648
rect 4348 46592 4404 46648
rect 4404 46592 4408 46648
rect 4344 46588 4408 46592
rect 4424 46648 4488 46652
rect 4424 46592 4428 46648
rect 4428 46592 4484 46648
rect 4484 46592 4488 46648
rect 4424 46588 4488 46592
rect 4504 46648 4568 46652
rect 4504 46592 4508 46648
rect 4508 46592 4564 46648
rect 4564 46592 4568 46648
rect 4504 46588 4568 46592
rect 34984 46648 35048 46652
rect 34984 46592 34988 46648
rect 34988 46592 35044 46648
rect 35044 46592 35048 46648
rect 34984 46588 35048 46592
rect 35064 46648 35128 46652
rect 35064 46592 35068 46648
rect 35068 46592 35124 46648
rect 35124 46592 35128 46648
rect 35064 46588 35128 46592
rect 35144 46648 35208 46652
rect 35144 46592 35148 46648
rect 35148 46592 35204 46648
rect 35204 46592 35208 46648
rect 35144 46588 35208 46592
rect 35224 46648 35288 46652
rect 35224 46592 35228 46648
rect 35228 46592 35284 46648
rect 35284 46592 35288 46648
rect 35224 46588 35288 46592
rect 19624 45982 19688 45986
rect 19624 45926 19628 45982
rect 19628 45926 19684 45982
rect 19684 45926 19688 45982
rect 19624 45922 19688 45926
rect 19704 45982 19768 45986
rect 19704 45926 19708 45982
rect 19708 45926 19764 45982
rect 19764 45926 19768 45982
rect 19704 45922 19768 45926
rect 19784 45982 19848 45986
rect 19784 45926 19788 45982
rect 19788 45926 19844 45982
rect 19844 45926 19848 45982
rect 19784 45922 19848 45926
rect 19864 45982 19928 45986
rect 19864 45926 19868 45982
rect 19868 45926 19924 45982
rect 19924 45926 19928 45982
rect 19864 45922 19928 45926
rect 50344 45982 50408 45986
rect 50344 45926 50348 45982
rect 50348 45926 50404 45982
rect 50404 45926 50408 45982
rect 50344 45922 50408 45926
rect 50424 45982 50488 45986
rect 50424 45926 50428 45982
rect 50428 45926 50484 45982
rect 50484 45926 50488 45982
rect 50424 45922 50488 45926
rect 50504 45982 50568 45986
rect 50504 45926 50508 45982
rect 50508 45926 50564 45982
rect 50564 45926 50568 45982
rect 50504 45922 50568 45926
rect 50584 45982 50648 45986
rect 50584 45926 50588 45982
rect 50588 45926 50644 45982
rect 50644 45926 50648 45982
rect 50584 45922 50648 45926
rect 4264 45316 4328 45320
rect 4264 45260 4268 45316
rect 4268 45260 4324 45316
rect 4324 45260 4328 45316
rect 4264 45256 4328 45260
rect 4344 45316 4408 45320
rect 4344 45260 4348 45316
rect 4348 45260 4404 45316
rect 4404 45260 4408 45316
rect 4344 45256 4408 45260
rect 4424 45316 4488 45320
rect 4424 45260 4428 45316
rect 4428 45260 4484 45316
rect 4484 45260 4488 45316
rect 4424 45256 4488 45260
rect 4504 45316 4568 45320
rect 4504 45260 4508 45316
rect 4508 45260 4564 45316
rect 4564 45260 4568 45316
rect 4504 45256 4568 45260
rect 34984 45316 35048 45320
rect 34984 45260 34988 45316
rect 34988 45260 35044 45316
rect 35044 45260 35048 45316
rect 34984 45256 35048 45260
rect 35064 45316 35128 45320
rect 35064 45260 35068 45316
rect 35068 45260 35124 45316
rect 35124 45260 35128 45316
rect 35064 45256 35128 45260
rect 35144 45316 35208 45320
rect 35144 45260 35148 45316
rect 35148 45260 35204 45316
rect 35204 45260 35208 45316
rect 35144 45256 35208 45260
rect 35224 45316 35288 45320
rect 35224 45260 35228 45316
rect 35228 45260 35284 45316
rect 35284 45260 35288 45316
rect 35224 45256 35288 45260
rect 19624 44650 19688 44654
rect 19624 44594 19628 44650
rect 19628 44594 19684 44650
rect 19684 44594 19688 44650
rect 19624 44590 19688 44594
rect 19704 44650 19768 44654
rect 19704 44594 19708 44650
rect 19708 44594 19764 44650
rect 19764 44594 19768 44650
rect 19704 44590 19768 44594
rect 19784 44650 19848 44654
rect 19784 44594 19788 44650
rect 19788 44594 19844 44650
rect 19844 44594 19848 44650
rect 19784 44590 19848 44594
rect 19864 44650 19928 44654
rect 19864 44594 19868 44650
rect 19868 44594 19924 44650
rect 19924 44594 19928 44650
rect 19864 44590 19928 44594
rect 50344 44650 50408 44654
rect 50344 44594 50348 44650
rect 50348 44594 50404 44650
rect 50404 44594 50408 44650
rect 50344 44590 50408 44594
rect 50424 44650 50488 44654
rect 50424 44594 50428 44650
rect 50428 44594 50484 44650
rect 50484 44594 50488 44650
rect 50424 44590 50488 44594
rect 50504 44650 50568 44654
rect 50504 44594 50508 44650
rect 50508 44594 50564 44650
rect 50564 44594 50568 44650
rect 50504 44590 50568 44594
rect 50584 44650 50648 44654
rect 50584 44594 50588 44650
rect 50588 44594 50644 44650
rect 50644 44594 50648 44650
rect 50584 44590 50648 44594
rect 4264 43984 4328 43988
rect 4264 43928 4268 43984
rect 4268 43928 4324 43984
rect 4324 43928 4328 43984
rect 4264 43924 4328 43928
rect 4344 43984 4408 43988
rect 4344 43928 4348 43984
rect 4348 43928 4404 43984
rect 4404 43928 4408 43984
rect 4344 43924 4408 43928
rect 4424 43984 4488 43988
rect 4424 43928 4428 43984
rect 4428 43928 4484 43984
rect 4484 43928 4488 43984
rect 4424 43924 4488 43928
rect 4504 43984 4568 43988
rect 4504 43928 4508 43984
rect 4508 43928 4564 43984
rect 4564 43928 4568 43984
rect 4504 43924 4568 43928
rect 34984 43984 35048 43988
rect 34984 43928 34988 43984
rect 34988 43928 35044 43984
rect 35044 43928 35048 43984
rect 34984 43924 35048 43928
rect 35064 43984 35128 43988
rect 35064 43928 35068 43984
rect 35068 43928 35124 43984
rect 35124 43928 35128 43984
rect 35064 43924 35128 43928
rect 35144 43984 35208 43988
rect 35144 43928 35148 43984
rect 35148 43928 35204 43984
rect 35204 43928 35208 43984
rect 35144 43924 35208 43928
rect 35224 43984 35288 43988
rect 35224 43928 35228 43984
rect 35228 43928 35284 43984
rect 35284 43928 35288 43984
rect 35224 43924 35288 43928
rect 19624 43318 19688 43322
rect 19624 43262 19628 43318
rect 19628 43262 19684 43318
rect 19684 43262 19688 43318
rect 19624 43258 19688 43262
rect 19704 43318 19768 43322
rect 19704 43262 19708 43318
rect 19708 43262 19764 43318
rect 19764 43262 19768 43318
rect 19704 43258 19768 43262
rect 19784 43318 19848 43322
rect 19784 43262 19788 43318
rect 19788 43262 19844 43318
rect 19844 43262 19848 43318
rect 19784 43258 19848 43262
rect 19864 43318 19928 43322
rect 19864 43262 19868 43318
rect 19868 43262 19924 43318
rect 19924 43262 19928 43318
rect 19864 43258 19928 43262
rect 50344 43318 50408 43322
rect 50344 43262 50348 43318
rect 50348 43262 50404 43318
rect 50404 43262 50408 43318
rect 50344 43258 50408 43262
rect 50424 43318 50488 43322
rect 50424 43262 50428 43318
rect 50428 43262 50484 43318
rect 50484 43262 50488 43318
rect 50424 43258 50488 43262
rect 50504 43318 50568 43322
rect 50504 43262 50508 43318
rect 50508 43262 50564 43318
rect 50564 43262 50568 43318
rect 50504 43258 50568 43262
rect 50584 43318 50648 43322
rect 50584 43262 50588 43318
rect 50588 43262 50644 43318
rect 50644 43262 50648 43318
rect 50584 43258 50648 43262
rect 4264 42652 4328 42656
rect 4264 42596 4268 42652
rect 4268 42596 4324 42652
rect 4324 42596 4328 42652
rect 4264 42592 4328 42596
rect 4344 42652 4408 42656
rect 4344 42596 4348 42652
rect 4348 42596 4404 42652
rect 4404 42596 4408 42652
rect 4344 42592 4408 42596
rect 4424 42652 4488 42656
rect 4424 42596 4428 42652
rect 4428 42596 4484 42652
rect 4484 42596 4488 42652
rect 4424 42592 4488 42596
rect 4504 42652 4568 42656
rect 4504 42596 4508 42652
rect 4508 42596 4564 42652
rect 4564 42596 4568 42652
rect 4504 42592 4568 42596
rect 34984 42652 35048 42656
rect 34984 42596 34988 42652
rect 34988 42596 35044 42652
rect 35044 42596 35048 42652
rect 34984 42592 35048 42596
rect 35064 42652 35128 42656
rect 35064 42596 35068 42652
rect 35068 42596 35124 42652
rect 35124 42596 35128 42652
rect 35064 42592 35128 42596
rect 35144 42652 35208 42656
rect 35144 42596 35148 42652
rect 35148 42596 35204 42652
rect 35204 42596 35208 42652
rect 35144 42592 35208 42596
rect 35224 42652 35288 42656
rect 35224 42596 35228 42652
rect 35228 42596 35284 42652
rect 35284 42596 35288 42652
rect 35224 42592 35288 42596
rect 19624 41986 19688 41990
rect 19624 41930 19628 41986
rect 19628 41930 19684 41986
rect 19684 41930 19688 41986
rect 19624 41926 19688 41930
rect 19704 41986 19768 41990
rect 19704 41930 19708 41986
rect 19708 41930 19764 41986
rect 19764 41930 19768 41986
rect 19704 41926 19768 41930
rect 19784 41986 19848 41990
rect 19784 41930 19788 41986
rect 19788 41930 19844 41986
rect 19844 41930 19848 41986
rect 19784 41926 19848 41930
rect 19864 41986 19928 41990
rect 19864 41930 19868 41986
rect 19868 41930 19924 41986
rect 19924 41930 19928 41986
rect 19864 41926 19928 41930
rect 50344 41986 50408 41990
rect 50344 41930 50348 41986
rect 50348 41930 50404 41986
rect 50404 41930 50408 41986
rect 50344 41926 50408 41930
rect 50424 41986 50488 41990
rect 50424 41930 50428 41986
rect 50428 41930 50484 41986
rect 50484 41930 50488 41986
rect 50424 41926 50488 41930
rect 50504 41986 50568 41990
rect 50504 41930 50508 41986
rect 50508 41930 50564 41986
rect 50564 41930 50568 41986
rect 50504 41926 50568 41930
rect 50584 41986 50648 41990
rect 50584 41930 50588 41986
rect 50588 41930 50644 41986
rect 50644 41930 50648 41986
rect 50584 41926 50648 41930
rect 4264 41320 4328 41324
rect 4264 41264 4268 41320
rect 4268 41264 4324 41320
rect 4324 41264 4328 41320
rect 4264 41260 4328 41264
rect 4344 41320 4408 41324
rect 4344 41264 4348 41320
rect 4348 41264 4404 41320
rect 4404 41264 4408 41320
rect 4344 41260 4408 41264
rect 4424 41320 4488 41324
rect 4424 41264 4428 41320
rect 4428 41264 4484 41320
rect 4484 41264 4488 41320
rect 4424 41260 4488 41264
rect 4504 41320 4568 41324
rect 4504 41264 4508 41320
rect 4508 41264 4564 41320
rect 4564 41264 4568 41320
rect 4504 41260 4568 41264
rect 34984 41320 35048 41324
rect 34984 41264 34988 41320
rect 34988 41264 35044 41320
rect 35044 41264 35048 41320
rect 34984 41260 35048 41264
rect 35064 41320 35128 41324
rect 35064 41264 35068 41320
rect 35068 41264 35124 41320
rect 35124 41264 35128 41320
rect 35064 41260 35128 41264
rect 35144 41320 35208 41324
rect 35144 41264 35148 41320
rect 35148 41264 35204 41320
rect 35204 41264 35208 41320
rect 35144 41260 35208 41264
rect 35224 41320 35288 41324
rect 35224 41264 35228 41320
rect 35228 41264 35284 41320
rect 35284 41264 35288 41320
rect 35224 41260 35288 41264
rect 19624 40654 19688 40658
rect 19624 40598 19628 40654
rect 19628 40598 19684 40654
rect 19684 40598 19688 40654
rect 19624 40594 19688 40598
rect 19704 40654 19768 40658
rect 19704 40598 19708 40654
rect 19708 40598 19764 40654
rect 19764 40598 19768 40654
rect 19704 40594 19768 40598
rect 19784 40654 19848 40658
rect 19784 40598 19788 40654
rect 19788 40598 19844 40654
rect 19844 40598 19848 40654
rect 19784 40594 19848 40598
rect 19864 40654 19928 40658
rect 19864 40598 19868 40654
rect 19868 40598 19924 40654
rect 19924 40598 19928 40654
rect 19864 40594 19928 40598
rect 50344 40654 50408 40658
rect 50344 40598 50348 40654
rect 50348 40598 50404 40654
rect 50404 40598 50408 40654
rect 50344 40594 50408 40598
rect 50424 40654 50488 40658
rect 50424 40598 50428 40654
rect 50428 40598 50484 40654
rect 50484 40598 50488 40654
rect 50424 40594 50488 40598
rect 50504 40654 50568 40658
rect 50504 40598 50508 40654
rect 50508 40598 50564 40654
rect 50564 40598 50568 40654
rect 50504 40594 50568 40598
rect 50584 40654 50648 40658
rect 50584 40598 50588 40654
rect 50588 40598 50644 40654
rect 50644 40598 50648 40654
rect 50584 40594 50648 40598
rect 4264 39988 4328 39992
rect 4264 39932 4268 39988
rect 4268 39932 4324 39988
rect 4324 39932 4328 39988
rect 4264 39928 4328 39932
rect 4344 39988 4408 39992
rect 4344 39932 4348 39988
rect 4348 39932 4404 39988
rect 4404 39932 4408 39988
rect 4344 39928 4408 39932
rect 4424 39988 4488 39992
rect 4424 39932 4428 39988
rect 4428 39932 4484 39988
rect 4484 39932 4488 39988
rect 4424 39928 4488 39932
rect 4504 39988 4568 39992
rect 4504 39932 4508 39988
rect 4508 39932 4564 39988
rect 4564 39932 4568 39988
rect 4504 39928 4568 39932
rect 34984 39988 35048 39992
rect 34984 39932 34988 39988
rect 34988 39932 35044 39988
rect 35044 39932 35048 39988
rect 34984 39928 35048 39932
rect 35064 39988 35128 39992
rect 35064 39932 35068 39988
rect 35068 39932 35124 39988
rect 35124 39932 35128 39988
rect 35064 39928 35128 39932
rect 35144 39988 35208 39992
rect 35144 39932 35148 39988
rect 35148 39932 35204 39988
rect 35204 39932 35208 39988
rect 35144 39928 35208 39932
rect 35224 39988 35288 39992
rect 35224 39932 35228 39988
rect 35228 39932 35284 39988
rect 35284 39932 35288 39988
rect 35224 39928 35288 39932
rect 19624 39322 19688 39326
rect 19624 39266 19628 39322
rect 19628 39266 19684 39322
rect 19684 39266 19688 39322
rect 19624 39262 19688 39266
rect 19704 39322 19768 39326
rect 19704 39266 19708 39322
rect 19708 39266 19764 39322
rect 19764 39266 19768 39322
rect 19704 39262 19768 39266
rect 19784 39322 19848 39326
rect 19784 39266 19788 39322
rect 19788 39266 19844 39322
rect 19844 39266 19848 39322
rect 19784 39262 19848 39266
rect 19864 39322 19928 39326
rect 19864 39266 19868 39322
rect 19868 39266 19924 39322
rect 19924 39266 19928 39322
rect 19864 39262 19928 39266
rect 50344 39322 50408 39326
rect 50344 39266 50348 39322
rect 50348 39266 50404 39322
rect 50404 39266 50408 39322
rect 50344 39262 50408 39266
rect 50424 39322 50488 39326
rect 50424 39266 50428 39322
rect 50428 39266 50484 39322
rect 50484 39266 50488 39322
rect 50424 39262 50488 39266
rect 50504 39322 50568 39326
rect 50504 39266 50508 39322
rect 50508 39266 50564 39322
rect 50564 39266 50568 39322
rect 50504 39262 50568 39266
rect 50584 39322 50648 39326
rect 50584 39266 50588 39322
rect 50588 39266 50644 39322
rect 50644 39266 50648 39322
rect 50584 39262 50648 39266
rect 4264 38656 4328 38660
rect 4264 38600 4268 38656
rect 4268 38600 4324 38656
rect 4324 38600 4328 38656
rect 4264 38596 4328 38600
rect 4344 38656 4408 38660
rect 4344 38600 4348 38656
rect 4348 38600 4404 38656
rect 4404 38600 4408 38656
rect 4344 38596 4408 38600
rect 4424 38656 4488 38660
rect 4424 38600 4428 38656
rect 4428 38600 4484 38656
rect 4484 38600 4488 38656
rect 4424 38596 4488 38600
rect 4504 38656 4568 38660
rect 4504 38600 4508 38656
rect 4508 38600 4564 38656
rect 4564 38600 4568 38656
rect 4504 38596 4568 38600
rect 34984 38656 35048 38660
rect 34984 38600 34988 38656
rect 34988 38600 35044 38656
rect 35044 38600 35048 38656
rect 34984 38596 35048 38600
rect 35064 38656 35128 38660
rect 35064 38600 35068 38656
rect 35068 38600 35124 38656
rect 35124 38600 35128 38656
rect 35064 38596 35128 38600
rect 35144 38656 35208 38660
rect 35144 38600 35148 38656
rect 35148 38600 35204 38656
rect 35204 38600 35208 38656
rect 35144 38596 35208 38600
rect 35224 38656 35288 38660
rect 35224 38600 35228 38656
rect 35228 38600 35284 38656
rect 35284 38600 35288 38656
rect 35224 38596 35288 38600
rect 19624 37990 19688 37994
rect 19624 37934 19628 37990
rect 19628 37934 19684 37990
rect 19684 37934 19688 37990
rect 19624 37930 19688 37934
rect 19704 37990 19768 37994
rect 19704 37934 19708 37990
rect 19708 37934 19764 37990
rect 19764 37934 19768 37990
rect 19704 37930 19768 37934
rect 19784 37990 19848 37994
rect 19784 37934 19788 37990
rect 19788 37934 19844 37990
rect 19844 37934 19848 37990
rect 19784 37930 19848 37934
rect 19864 37990 19928 37994
rect 19864 37934 19868 37990
rect 19868 37934 19924 37990
rect 19924 37934 19928 37990
rect 19864 37930 19928 37934
rect 50344 37990 50408 37994
rect 50344 37934 50348 37990
rect 50348 37934 50404 37990
rect 50404 37934 50408 37990
rect 50344 37930 50408 37934
rect 50424 37990 50488 37994
rect 50424 37934 50428 37990
rect 50428 37934 50484 37990
rect 50484 37934 50488 37990
rect 50424 37930 50488 37934
rect 50504 37990 50568 37994
rect 50504 37934 50508 37990
rect 50508 37934 50564 37990
rect 50564 37934 50568 37990
rect 50504 37930 50568 37934
rect 50584 37990 50648 37994
rect 50584 37934 50588 37990
rect 50588 37934 50644 37990
rect 50644 37934 50648 37990
rect 50584 37930 50648 37934
rect 4264 37324 4328 37328
rect 4264 37268 4268 37324
rect 4268 37268 4324 37324
rect 4324 37268 4328 37324
rect 4264 37264 4328 37268
rect 4344 37324 4408 37328
rect 4344 37268 4348 37324
rect 4348 37268 4404 37324
rect 4404 37268 4408 37324
rect 4344 37264 4408 37268
rect 4424 37324 4488 37328
rect 4424 37268 4428 37324
rect 4428 37268 4484 37324
rect 4484 37268 4488 37324
rect 4424 37264 4488 37268
rect 4504 37324 4568 37328
rect 4504 37268 4508 37324
rect 4508 37268 4564 37324
rect 4564 37268 4568 37324
rect 4504 37264 4568 37268
rect 34984 37324 35048 37328
rect 34984 37268 34988 37324
rect 34988 37268 35044 37324
rect 35044 37268 35048 37324
rect 34984 37264 35048 37268
rect 35064 37324 35128 37328
rect 35064 37268 35068 37324
rect 35068 37268 35124 37324
rect 35124 37268 35128 37324
rect 35064 37264 35128 37268
rect 35144 37324 35208 37328
rect 35144 37268 35148 37324
rect 35148 37268 35204 37324
rect 35204 37268 35208 37324
rect 35144 37264 35208 37268
rect 35224 37324 35288 37328
rect 35224 37268 35228 37324
rect 35228 37268 35284 37324
rect 35284 37268 35288 37324
rect 35224 37264 35288 37268
rect 19624 36658 19688 36662
rect 19624 36602 19628 36658
rect 19628 36602 19684 36658
rect 19684 36602 19688 36658
rect 19624 36598 19688 36602
rect 19704 36658 19768 36662
rect 19704 36602 19708 36658
rect 19708 36602 19764 36658
rect 19764 36602 19768 36658
rect 19704 36598 19768 36602
rect 19784 36658 19848 36662
rect 19784 36602 19788 36658
rect 19788 36602 19844 36658
rect 19844 36602 19848 36658
rect 19784 36598 19848 36602
rect 19864 36658 19928 36662
rect 19864 36602 19868 36658
rect 19868 36602 19924 36658
rect 19924 36602 19928 36658
rect 19864 36598 19928 36602
rect 50344 36658 50408 36662
rect 50344 36602 50348 36658
rect 50348 36602 50404 36658
rect 50404 36602 50408 36658
rect 50344 36598 50408 36602
rect 50424 36658 50488 36662
rect 50424 36602 50428 36658
rect 50428 36602 50484 36658
rect 50484 36602 50488 36658
rect 50424 36598 50488 36602
rect 50504 36658 50568 36662
rect 50504 36602 50508 36658
rect 50508 36602 50564 36658
rect 50564 36602 50568 36658
rect 50504 36598 50568 36602
rect 50584 36658 50648 36662
rect 50584 36602 50588 36658
rect 50588 36602 50644 36658
rect 50644 36602 50648 36658
rect 50584 36598 50648 36602
rect 4264 35992 4328 35996
rect 4264 35936 4268 35992
rect 4268 35936 4324 35992
rect 4324 35936 4328 35992
rect 4264 35932 4328 35936
rect 4344 35992 4408 35996
rect 4344 35936 4348 35992
rect 4348 35936 4404 35992
rect 4404 35936 4408 35992
rect 4344 35932 4408 35936
rect 4424 35992 4488 35996
rect 4424 35936 4428 35992
rect 4428 35936 4484 35992
rect 4484 35936 4488 35992
rect 4424 35932 4488 35936
rect 4504 35992 4568 35996
rect 4504 35936 4508 35992
rect 4508 35936 4564 35992
rect 4564 35936 4568 35992
rect 4504 35932 4568 35936
rect 34984 35992 35048 35996
rect 34984 35936 34988 35992
rect 34988 35936 35044 35992
rect 35044 35936 35048 35992
rect 34984 35932 35048 35936
rect 35064 35992 35128 35996
rect 35064 35936 35068 35992
rect 35068 35936 35124 35992
rect 35124 35936 35128 35992
rect 35064 35932 35128 35936
rect 35144 35992 35208 35996
rect 35144 35936 35148 35992
rect 35148 35936 35204 35992
rect 35204 35936 35208 35992
rect 35144 35932 35208 35936
rect 35224 35992 35288 35996
rect 35224 35936 35228 35992
rect 35228 35936 35284 35992
rect 35284 35936 35288 35992
rect 35224 35932 35288 35936
rect 19624 35326 19688 35330
rect 19624 35270 19628 35326
rect 19628 35270 19684 35326
rect 19684 35270 19688 35326
rect 19624 35266 19688 35270
rect 19704 35326 19768 35330
rect 19704 35270 19708 35326
rect 19708 35270 19764 35326
rect 19764 35270 19768 35326
rect 19704 35266 19768 35270
rect 19784 35326 19848 35330
rect 19784 35270 19788 35326
rect 19788 35270 19844 35326
rect 19844 35270 19848 35326
rect 19784 35266 19848 35270
rect 19864 35326 19928 35330
rect 19864 35270 19868 35326
rect 19868 35270 19924 35326
rect 19924 35270 19928 35326
rect 19864 35266 19928 35270
rect 50344 35326 50408 35330
rect 50344 35270 50348 35326
rect 50348 35270 50404 35326
rect 50404 35270 50408 35326
rect 50344 35266 50408 35270
rect 50424 35326 50488 35330
rect 50424 35270 50428 35326
rect 50428 35270 50484 35326
rect 50484 35270 50488 35326
rect 50424 35266 50488 35270
rect 50504 35326 50568 35330
rect 50504 35270 50508 35326
rect 50508 35270 50564 35326
rect 50564 35270 50568 35326
rect 50504 35266 50568 35270
rect 50584 35326 50648 35330
rect 50584 35270 50588 35326
rect 50588 35270 50644 35326
rect 50644 35270 50648 35326
rect 50584 35266 50648 35270
rect 4264 34660 4328 34664
rect 4264 34604 4268 34660
rect 4268 34604 4324 34660
rect 4324 34604 4328 34660
rect 4264 34600 4328 34604
rect 4344 34660 4408 34664
rect 4344 34604 4348 34660
rect 4348 34604 4404 34660
rect 4404 34604 4408 34660
rect 4344 34600 4408 34604
rect 4424 34660 4488 34664
rect 4424 34604 4428 34660
rect 4428 34604 4484 34660
rect 4484 34604 4488 34660
rect 4424 34600 4488 34604
rect 4504 34660 4568 34664
rect 4504 34604 4508 34660
rect 4508 34604 4564 34660
rect 4564 34604 4568 34660
rect 4504 34600 4568 34604
rect 34984 34660 35048 34664
rect 34984 34604 34988 34660
rect 34988 34604 35044 34660
rect 35044 34604 35048 34660
rect 34984 34600 35048 34604
rect 35064 34660 35128 34664
rect 35064 34604 35068 34660
rect 35068 34604 35124 34660
rect 35124 34604 35128 34660
rect 35064 34600 35128 34604
rect 35144 34660 35208 34664
rect 35144 34604 35148 34660
rect 35148 34604 35204 34660
rect 35204 34604 35208 34660
rect 35144 34600 35208 34604
rect 35224 34660 35288 34664
rect 35224 34604 35228 34660
rect 35228 34604 35284 34660
rect 35284 34604 35288 34660
rect 35224 34600 35288 34604
rect 19624 33994 19688 33998
rect 19624 33938 19628 33994
rect 19628 33938 19684 33994
rect 19684 33938 19688 33994
rect 19624 33934 19688 33938
rect 19704 33994 19768 33998
rect 19704 33938 19708 33994
rect 19708 33938 19764 33994
rect 19764 33938 19768 33994
rect 19704 33934 19768 33938
rect 19784 33994 19848 33998
rect 19784 33938 19788 33994
rect 19788 33938 19844 33994
rect 19844 33938 19848 33994
rect 19784 33934 19848 33938
rect 19864 33994 19928 33998
rect 19864 33938 19868 33994
rect 19868 33938 19924 33994
rect 19924 33938 19928 33994
rect 19864 33934 19928 33938
rect 50344 33994 50408 33998
rect 50344 33938 50348 33994
rect 50348 33938 50404 33994
rect 50404 33938 50408 33994
rect 50344 33934 50408 33938
rect 50424 33994 50488 33998
rect 50424 33938 50428 33994
rect 50428 33938 50484 33994
rect 50484 33938 50488 33994
rect 50424 33934 50488 33938
rect 50504 33994 50568 33998
rect 50504 33938 50508 33994
rect 50508 33938 50564 33994
rect 50564 33938 50568 33994
rect 50504 33934 50568 33938
rect 50584 33994 50648 33998
rect 50584 33938 50588 33994
rect 50588 33938 50644 33994
rect 50644 33938 50648 33994
rect 50584 33934 50648 33938
rect 4264 33328 4328 33332
rect 4264 33272 4268 33328
rect 4268 33272 4324 33328
rect 4324 33272 4328 33328
rect 4264 33268 4328 33272
rect 4344 33328 4408 33332
rect 4344 33272 4348 33328
rect 4348 33272 4404 33328
rect 4404 33272 4408 33328
rect 4344 33268 4408 33272
rect 4424 33328 4488 33332
rect 4424 33272 4428 33328
rect 4428 33272 4484 33328
rect 4484 33272 4488 33328
rect 4424 33268 4488 33272
rect 4504 33328 4568 33332
rect 4504 33272 4508 33328
rect 4508 33272 4564 33328
rect 4564 33272 4568 33328
rect 4504 33268 4568 33272
rect 34984 33328 35048 33332
rect 34984 33272 34988 33328
rect 34988 33272 35044 33328
rect 35044 33272 35048 33328
rect 34984 33268 35048 33272
rect 35064 33328 35128 33332
rect 35064 33272 35068 33328
rect 35068 33272 35124 33328
rect 35124 33272 35128 33328
rect 35064 33268 35128 33272
rect 35144 33328 35208 33332
rect 35144 33272 35148 33328
rect 35148 33272 35204 33328
rect 35204 33272 35208 33328
rect 35144 33268 35208 33272
rect 35224 33328 35288 33332
rect 35224 33272 35228 33328
rect 35228 33272 35284 33328
rect 35284 33272 35288 33328
rect 35224 33268 35288 33272
rect 19624 32662 19688 32666
rect 19624 32606 19628 32662
rect 19628 32606 19684 32662
rect 19684 32606 19688 32662
rect 19624 32602 19688 32606
rect 19704 32662 19768 32666
rect 19704 32606 19708 32662
rect 19708 32606 19764 32662
rect 19764 32606 19768 32662
rect 19704 32602 19768 32606
rect 19784 32662 19848 32666
rect 19784 32606 19788 32662
rect 19788 32606 19844 32662
rect 19844 32606 19848 32662
rect 19784 32602 19848 32606
rect 19864 32662 19928 32666
rect 19864 32606 19868 32662
rect 19868 32606 19924 32662
rect 19924 32606 19928 32662
rect 19864 32602 19928 32606
rect 50344 32662 50408 32666
rect 50344 32606 50348 32662
rect 50348 32606 50404 32662
rect 50404 32606 50408 32662
rect 50344 32602 50408 32606
rect 50424 32662 50488 32666
rect 50424 32606 50428 32662
rect 50428 32606 50484 32662
rect 50484 32606 50488 32662
rect 50424 32602 50488 32606
rect 50504 32662 50568 32666
rect 50504 32606 50508 32662
rect 50508 32606 50564 32662
rect 50564 32606 50568 32662
rect 50504 32602 50568 32606
rect 50584 32662 50648 32666
rect 50584 32606 50588 32662
rect 50588 32606 50644 32662
rect 50644 32606 50648 32662
rect 50584 32602 50648 32606
rect 4264 31996 4328 32000
rect 4264 31940 4268 31996
rect 4268 31940 4324 31996
rect 4324 31940 4328 31996
rect 4264 31936 4328 31940
rect 4344 31996 4408 32000
rect 4344 31940 4348 31996
rect 4348 31940 4404 31996
rect 4404 31940 4408 31996
rect 4344 31936 4408 31940
rect 4424 31996 4488 32000
rect 4424 31940 4428 31996
rect 4428 31940 4484 31996
rect 4484 31940 4488 31996
rect 4424 31936 4488 31940
rect 4504 31996 4568 32000
rect 4504 31940 4508 31996
rect 4508 31940 4564 31996
rect 4564 31940 4568 31996
rect 4504 31936 4568 31940
rect 34984 31996 35048 32000
rect 34984 31940 34988 31996
rect 34988 31940 35044 31996
rect 35044 31940 35048 31996
rect 34984 31936 35048 31940
rect 35064 31996 35128 32000
rect 35064 31940 35068 31996
rect 35068 31940 35124 31996
rect 35124 31940 35128 31996
rect 35064 31936 35128 31940
rect 35144 31996 35208 32000
rect 35144 31940 35148 31996
rect 35148 31940 35204 31996
rect 35204 31940 35208 31996
rect 35144 31936 35208 31940
rect 35224 31996 35288 32000
rect 35224 31940 35228 31996
rect 35228 31940 35284 31996
rect 35284 31940 35288 31996
rect 35224 31936 35288 31940
rect 19624 31330 19688 31334
rect 19624 31274 19628 31330
rect 19628 31274 19684 31330
rect 19684 31274 19688 31330
rect 19624 31270 19688 31274
rect 19704 31330 19768 31334
rect 19704 31274 19708 31330
rect 19708 31274 19764 31330
rect 19764 31274 19768 31330
rect 19704 31270 19768 31274
rect 19784 31330 19848 31334
rect 19784 31274 19788 31330
rect 19788 31274 19844 31330
rect 19844 31274 19848 31330
rect 19784 31270 19848 31274
rect 19864 31330 19928 31334
rect 19864 31274 19868 31330
rect 19868 31274 19924 31330
rect 19924 31274 19928 31330
rect 19864 31270 19928 31274
rect 50344 31330 50408 31334
rect 50344 31274 50348 31330
rect 50348 31274 50404 31330
rect 50404 31274 50408 31330
rect 50344 31270 50408 31274
rect 50424 31330 50488 31334
rect 50424 31274 50428 31330
rect 50428 31274 50484 31330
rect 50484 31274 50488 31330
rect 50424 31270 50488 31274
rect 50504 31330 50568 31334
rect 50504 31274 50508 31330
rect 50508 31274 50564 31330
rect 50564 31274 50568 31330
rect 50504 31270 50568 31274
rect 50584 31330 50648 31334
rect 50584 31274 50588 31330
rect 50588 31274 50644 31330
rect 50644 31274 50648 31330
rect 50584 31270 50648 31274
rect 4264 30664 4328 30668
rect 4264 30608 4268 30664
rect 4268 30608 4324 30664
rect 4324 30608 4328 30664
rect 4264 30604 4328 30608
rect 4344 30664 4408 30668
rect 4344 30608 4348 30664
rect 4348 30608 4404 30664
rect 4404 30608 4408 30664
rect 4344 30604 4408 30608
rect 4424 30664 4488 30668
rect 4424 30608 4428 30664
rect 4428 30608 4484 30664
rect 4484 30608 4488 30664
rect 4424 30604 4488 30608
rect 4504 30664 4568 30668
rect 4504 30608 4508 30664
rect 4508 30608 4564 30664
rect 4564 30608 4568 30664
rect 4504 30604 4568 30608
rect 34984 30664 35048 30668
rect 34984 30608 34988 30664
rect 34988 30608 35044 30664
rect 35044 30608 35048 30664
rect 34984 30604 35048 30608
rect 35064 30664 35128 30668
rect 35064 30608 35068 30664
rect 35068 30608 35124 30664
rect 35124 30608 35128 30664
rect 35064 30604 35128 30608
rect 35144 30664 35208 30668
rect 35144 30608 35148 30664
rect 35148 30608 35204 30664
rect 35204 30608 35208 30664
rect 35144 30604 35208 30608
rect 35224 30664 35288 30668
rect 35224 30608 35228 30664
rect 35228 30608 35284 30664
rect 35284 30608 35288 30664
rect 35224 30604 35288 30608
rect 19624 29998 19688 30002
rect 19624 29942 19628 29998
rect 19628 29942 19684 29998
rect 19684 29942 19688 29998
rect 19624 29938 19688 29942
rect 19704 29998 19768 30002
rect 19704 29942 19708 29998
rect 19708 29942 19764 29998
rect 19764 29942 19768 29998
rect 19704 29938 19768 29942
rect 19784 29998 19848 30002
rect 19784 29942 19788 29998
rect 19788 29942 19844 29998
rect 19844 29942 19848 29998
rect 19784 29938 19848 29942
rect 19864 29998 19928 30002
rect 19864 29942 19868 29998
rect 19868 29942 19924 29998
rect 19924 29942 19928 29998
rect 19864 29938 19928 29942
rect 50344 29998 50408 30002
rect 50344 29942 50348 29998
rect 50348 29942 50404 29998
rect 50404 29942 50408 29998
rect 50344 29938 50408 29942
rect 50424 29998 50488 30002
rect 50424 29942 50428 29998
rect 50428 29942 50484 29998
rect 50484 29942 50488 29998
rect 50424 29938 50488 29942
rect 50504 29998 50568 30002
rect 50504 29942 50508 29998
rect 50508 29942 50564 29998
rect 50564 29942 50568 29998
rect 50504 29938 50568 29942
rect 50584 29998 50648 30002
rect 50584 29942 50588 29998
rect 50588 29942 50644 29998
rect 50644 29942 50648 29998
rect 50584 29938 50648 29942
rect 4264 29332 4328 29336
rect 4264 29276 4268 29332
rect 4268 29276 4324 29332
rect 4324 29276 4328 29332
rect 4264 29272 4328 29276
rect 4344 29332 4408 29336
rect 4344 29276 4348 29332
rect 4348 29276 4404 29332
rect 4404 29276 4408 29332
rect 4344 29272 4408 29276
rect 4424 29332 4488 29336
rect 4424 29276 4428 29332
rect 4428 29276 4484 29332
rect 4484 29276 4488 29332
rect 4424 29272 4488 29276
rect 4504 29332 4568 29336
rect 4504 29276 4508 29332
rect 4508 29276 4564 29332
rect 4564 29276 4568 29332
rect 4504 29272 4568 29276
rect 34984 29332 35048 29336
rect 34984 29276 34988 29332
rect 34988 29276 35044 29332
rect 35044 29276 35048 29332
rect 34984 29272 35048 29276
rect 35064 29332 35128 29336
rect 35064 29276 35068 29332
rect 35068 29276 35124 29332
rect 35124 29276 35128 29332
rect 35064 29272 35128 29276
rect 35144 29332 35208 29336
rect 35144 29276 35148 29332
rect 35148 29276 35204 29332
rect 35204 29276 35208 29332
rect 35144 29272 35208 29276
rect 35224 29332 35288 29336
rect 35224 29276 35228 29332
rect 35228 29276 35284 29332
rect 35284 29276 35288 29332
rect 35224 29272 35288 29276
rect 8128 28902 8192 28966
rect 19624 28666 19688 28670
rect 19624 28610 19628 28666
rect 19628 28610 19684 28666
rect 19684 28610 19688 28666
rect 19624 28606 19688 28610
rect 19704 28666 19768 28670
rect 19704 28610 19708 28666
rect 19708 28610 19764 28666
rect 19764 28610 19768 28666
rect 19704 28606 19768 28610
rect 19784 28666 19848 28670
rect 19784 28610 19788 28666
rect 19788 28610 19844 28666
rect 19844 28610 19848 28666
rect 19784 28606 19848 28610
rect 19864 28666 19928 28670
rect 19864 28610 19868 28666
rect 19868 28610 19924 28666
rect 19924 28610 19928 28666
rect 19864 28606 19928 28610
rect 50344 28666 50408 28670
rect 50344 28610 50348 28666
rect 50348 28610 50404 28666
rect 50404 28610 50408 28666
rect 50344 28606 50408 28610
rect 50424 28666 50488 28670
rect 50424 28610 50428 28666
rect 50428 28610 50484 28666
rect 50484 28610 50488 28666
rect 50424 28606 50488 28610
rect 50504 28666 50568 28670
rect 50504 28610 50508 28666
rect 50508 28610 50564 28666
rect 50564 28610 50568 28666
rect 50504 28606 50568 28610
rect 50584 28666 50648 28670
rect 50584 28610 50588 28666
rect 50588 28610 50644 28666
rect 50644 28610 50648 28666
rect 50584 28606 50648 28610
rect 4264 28000 4328 28004
rect 4264 27944 4268 28000
rect 4268 27944 4324 28000
rect 4324 27944 4328 28000
rect 4264 27940 4328 27944
rect 4344 28000 4408 28004
rect 4344 27944 4348 28000
rect 4348 27944 4404 28000
rect 4404 27944 4408 28000
rect 4344 27940 4408 27944
rect 4424 28000 4488 28004
rect 4424 27944 4428 28000
rect 4428 27944 4484 28000
rect 4484 27944 4488 28000
rect 4424 27940 4488 27944
rect 4504 28000 4568 28004
rect 4504 27944 4508 28000
rect 4508 27944 4564 28000
rect 4564 27944 4568 28000
rect 4504 27940 4568 27944
rect 34984 28000 35048 28004
rect 34984 27944 34988 28000
rect 34988 27944 35044 28000
rect 35044 27944 35048 28000
rect 34984 27940 35048 27944
rect 35064 28000 35128 28004
rect 35064 27944 35068 28000
rect 35068 27944 35124 28000
rect 35124 27944 35128 28000
rect 35064 27940 35128 27944
rect 35144 28000 35208 28004
rect 35144 27944 35148 28000
rect 35148 27944 35204 28000
rect 35204 27944 35208 28000
rect 35144 27940 35208 27944
rect 35224 28000 35288 28004
rect 35224 27944 35228 28000
rect 35228 27944 35284 28000
rect 35284 27944 35288 28000
rect 35224 27940 35288 27944
rect 19624 27334 19688 27338
rect 19624 27278 19628 27334
rect 19628 27278 19684 27334
rect 19684 27278 19688 27334
rect 19624 27274 19688 27278
rect 19704 27334 19768 27338
rect 19704 27278 19708 27334
rect 19708 27278 19764 27334
rect 19764 27278 19768 27334
rect 19704 27274 19768 27278
rect 19784 27334 19848 27338
rect 19784 27278 19788 27334
rect 19788 27278 19844 27334
rect 19844 27278 19848 27334
rect 19784 27274 19848 27278
rect 19864 27334 19928 27338
rect 19864 27278 19868 27334
rect 19868 27278 19924 27334
rect 19924 27278 19928 27334
rect 19864 27274 19928 27278
rect 50344 27334 50408 27338
rect 50344 27278 50348 27334
rect 50348 27278 50404 27334
rect 50404 27278 50408 27334
rect 50344 27274 50408 27278
rect 50424 27334 50488 27338
rect 50424 27278 50428 27334
rect 50428 27278 50484 27334
rect 50484 27278 50488 27334
rect 50424 27274 50488 27278
rect 50504 27334 50568 27338
rect 50504 27278 50508 27334
rect 50508 27278 50564 27334
rect 50564 27278 50568 27334
rect 50504 27274 50568 27278
rect 50584 27334 50648 27338
rect 50584 27278 50588 27334
rect 50588 27278 50644 27334
rect 50644 27278 50648 27334
rect 50584 27274 50648 27278
rect 4264 26668 4328 26672
rect 4264 26612 4268 26668
rect 4268 26612 4324 26668
rect 4324 26612 4328 26668
rect 4264 26608 4328 26612
rect 4344 26668 4408 26672
rect 4344 26612 4348 26668
rect 4348 26612 4404 26668
rect 4404 26612 4408 26668
rect 4344 26608 4408 26612
rect 4424 26668 4488 26672
rect 4424 26612 4428 26668
rect 4428 26612 4484 26668
rect 4484 26612 4488 26668
rect 4424 26608 4488 26612
rect 4504 26668 4568 26672
rect 4504 26612 4508 26668
rect 4508 26612 4564 26668
rect 4564 26612 4568 26668
rect 4504 26608 4568 26612
rect 34984 26668 35048 26672
rect 34984 26612 34988 26668
rect 34988 26612 35044 26668
rect 35044 26612 35048 26668
rect 34984 26608 35048 26612
rect 35064 26668 35128 26672
rect 35064 26612 35068 26668
rect 35068 26612 35124 26668
rect 35124 26612 35128 26668
rect 35064 26608 35128 26612
rect 35144 26668 35208 26672
rect 35144 26612 35148 26668
rect 35148 26612 35204 26668
rect 35204 26612 35208 26668
rect 35144 26608 35208 26612
rect 35224 26668 35288 26672
rect 35224 26612 35228 26668
rect 35228 26612 35284 26668
rect 35284 26612 35288 26668
rect 35224 26608 35288 26612
rect 8320 26150 8384 26154
rect 8320 26094 8372 26150
rect 8372 26094 8384 26150
rect 8320 26090 8384 26094
rect 19624 26002 19688 26006
rect 19624 25946 19628 26002
rect 19628 25946 19684 26002
rect 19684 25946 19688 26002
rect 19624 25942 19688 25946
rect 19704 26002 19768 26006
rect 19704 25946 19708 26002
rect 19708 25946 19764 26002
rect 19764 25946 19768 26002
rect 19704 25942 19768 25946
rect 19784 26002 19848 26006
rect 19784 25946 19788 26002
rect 19788 25946 19844 26002
rect 19844 25946 19848 26002
rect 19784 25942 19848 25946
rect 19864 26002 19928 26006
rect 19864 25946 19868 26002
rect 19868 25946 19924 26002
rect 19924 25946 19928 26002
rect 19864 25942 19928 25946
rect 50344 26002 50408 26006
rect 50344 25946 50348 26002
rect 50348 25946 50404 26002
rect 50404 25946 50408 26002
rect 50344 25942 50408 25946
rect 50424 26002 50488 26006
rect 50424 25946 50428 26002
rect 50428 25946 50484 26002
rect 50484 25946 50488 26002
rect 50424 25942 50488 25946
rect 50504 26002 50568 26006
rect 50504 25946 50508 26002
rect 50508 25946 50564 26002
rect 50564 25946 50568 26002
rect 50504 25942 50568 25946
rect 50584 26002 50648 26006
rect 50584 25946 50588 26002
rect 50588 25946 50644 26002
rect 50644 25946 50648 26002
rect 50584 25942 50648 25946
rect 4264 25336 4328 25340
rect 4264 25280 4268 25336
rect 4268 25280 4324 25336
rect 4324 25280 4328 25336
rect 4264 25276 4328 25280
rect 4344 25336 4408 25340
rect 4344 25280 4348 25336
rect 4348 25280 4404 25336
rect 4404 25280 4408 25336
rect 4344 25276 4408 25280
rect 4424 25336 4488 25340
rect 4424 25280 4428 25336
rect 4428 25280 4484 25336
rect 4484 25280 4488 25336
rect 4424 25276 4488 25280
rect 4504 25336 4568 25340
rect 4504 25280 4508 25336
rect 4508 25280 4564 25336
rect 4564 25280 4568 25336
rect 4504 25276 4568 25280
rect 34984 25336 35048 25340
rect 34984 25280 34988 25336
rect 34988 25280 35044 25336
rect 35044 25280 35048 25336
rect 34984 25276 35048 25280
rect 35064 25336 35128 25340
rect 35064 25280 35068 25336
rect 35068 25280 35124 25336
rect 35124 25280 35128 25336
rect 35064 25276 35128 25280
rect 35144 25336 35208 25340
rect 35144 25280 35148 25336
rect 35148 25280 35204 25336
rect 35204 25280 35208 25336
rect 35144 25276 35208 25280
rect 35224 25336 35288 25340
rect 35224 25280 35228 25336
rect 35228 25280 35284 25336
rect 35284 25280 35288 25336
rect 35224 25276 35288 25280
rect 19624 24670 19688 24674
rect 19624 24614 19628 24670
rect 19628 24614 19684 24670
rect 19684 24614 19688 24670
rect 19624 24610 19688 24614
rect 19704 24670 19768 24674
rect 19704 24614 19708 24670
rect 19708 24614 19764 24670
rect 19764 24614 19768 24670
rect 19704 24610 19768 24614
rect 19784 24670 19848 24674
rect 19784 24614 19788 24670
rect 19788 24614 19844 24670
rect 19844 24614 19848 24670
rect 19784 24610 19848 24614
rect 19864 24670 19928 24674
rect 19864 24614 19868 24670
rect 19868 24614 19924 24670
rect 19924 24614 19928 24670
rect 19864 24610 19928 24614
rect 50344 24670 50408 24674
rect 50344 24614 50348 24670
rect 50348 24614 50404 24670
rect 50404 24614 50408 24670
rect 50344 24610 50408 24614
rect 50424 24670 50488 24674
rect 50424 24614 50428 24670
rect 50428 24614 50484 24670
rect 50484 24614 50488 24670
rect 50424 24610 50488 24614
rect 50504 24670 50568 24674
rect 50504 24614 50508 24670
rect 50508 24614 50564 24670
rect 50564 24614 50568 24670
rect 50504 24610 50568 24614
rect 50584 24670 50648 24674
rect 50584 24614 50588 24670
rect 50588 24614 50644 24670
rect 50644 24614 50648 24670
rect 50584 24610 50648 24614
rect 4264 24004 4328 24008
rect 4264 23948 4268 24004
rect 4268 23948 4324 24004
rect 4324 23948 4328 24004
rect 4264 23944 4328 23948
rect 4344 24004 4408 24008
rect 4344 23948 4348 24004
rect 4348 23948 4404 24004
rect 4404 23948 4408 24004
rect 4344 23944 4408 23948
rect 4424 24004 4488 24008
rect 4424 23948 4428 24004
rect 4428 23948 4484 24004
rect 4484 23948 4488 24004
rect 4424 23944 4488 23948
rect 4504 24004 4568 24008
rect 4504 23948 4508 24004
rect 4508 23948 4564 24004
rect 4564 23948 4568 24004
rect 4504 23944 4568 23948
rect 34984 24004 35048 24008
rect 34984 23948 34988 24004
rect 34988 23948 35044 24004
rect 35044 23948 35048 24004
rect 34984 23944 35048 23948
rect 35064 24004 35128 24008
rect 35064 23948 35068 24004
rect 35068 23948 35124 24004
rect 35124 23948 35128 24004
rect 35064 23944 35128 23948
rect 35144 24004 35208 24008
rect 35144 23948 35148 24004
rect 35148 23948 35204 24004
rect 35204 23948 35208 24004
rect 35144 23944 35208 23948
rect 35224 24004 35288 24008
rect 35224 23948 35228 24004
rect 35228 23948 35284 24004
rect 35284 23948 35288 24004
rect 35224 23944 35288 23948
rect 19624 23338 19688 23342
rect 19624 23282 19628 23338
rect 19628 23282 19684 23338
rect 19684 23282 19688 23338
rect 19624 23278 19688 23282
rect 19704 23338 19768 23342
rect 19704 23282 19708 23338
rect 19708 23282 19764 23338
rect 19764 23282 19768 23338
rect 19704 23278 19768 23282
rect 19784 23338 19848 23342
rect 19784 23282 19788 23338
rect 19788 23282 19844 23338
rect 19844 23282 19848 23338
rect 19784 23278 19848 23282
rect 19864 23338 19928 23342
rect 19864 23282 19868 23338
rect 19868 23282 19924 23338
rect 19924 23282 19928 23338
rect 19864 23278 19928 23282
rect 50344 23338 50408 23342
rect 50344 23282 50348 23338
rect 50348 23282 50404 23338
rect 50404 23282 50408 23338
rect 50344 23278 50408 23282
rect 50424 23338 50488 23342
rect 50424 23282 50428 23338
rect 50428 23282 50484 23338
rect 50484 23282 50488 23338
rect 50424 23278 50488 23282
rect 50504 23338 50568 23342
rect 50504 23282 50508 23338
rect 50508 23282 50564 23338
rect 50564 23282 50568 23338
rect 50504 23278 50568 23282
rect 50584 23338 50648 23342
rect 50584 23282 50588 23338
rect 50588 23282 50644 23338
rect 50644 23282 50648 23338
rect 50584 23278 50648 23282
rect 4264 22672 4328 22676
rect 4264 22616 4268 22672
rect 4268 22616 4324 22672
rect 4324 22616 4328 22672
rect 4264 22612 4328 22616
rect 4344 22672 4408 22676
rect 4344 22616 4348 22672
rect 4348 22616 4404 22672
rect 4404 22616 4408 22672
rect 4344 22612 4408 22616
rect 4424 22672 4488 22676
rect 4424 22616 4428 22672
rect 4428 22616 4484 22672
rect 4484 22616 4488 22672
rect 4424 22612 4488 22616
rect 4504 22672 4568 22676
rect 4504 22616 4508 22672
rect 4508 22616 4564 22672
rect 4564 22616 4568 22672
rect 4504 22612 4568 22616
rect 34984 22672 35048 22676
rect 34984 22616 34988 22672
rect 34988 22616 35044 22672
rect 35044 22616 35048 22672
rect 34984 22612 35048 22616
rect 35064 22672 35128 22676
rect 35064 22616 35068 22672
rect 35068 22616 35124 22672
rect 35124 22616 35128 22672
rect 35064 22612 35128 22616
rect 35144 22672 35208 22676
rect 35144 22616 35148 22672
rect 35148 22616 35204 22672
rect 35204 22616 35208 22672
rect 35144 22612 35208 22616
rect 35224 22672 35288 22676
rect 35224 22616 35228 22672
rect 35228 22616 35284 22672
rect 35284 22616 35288 22672
rect 35224 22612 35288 22616
rect 19624 22006 19688 22010
rect 19624 21950 19628 22006
rect 19628 21950 19684 22006
rect 19684 21950 19688 22006
rect 19624 21946 19688 21950
rect 19704 22006 19768 22010
rect 19704 21950 19708 22006
rect 19708 21950 19764 22006
rect 19764 21950 19768 22006
rect 19704 21946 19768 21950
rect 19784 22006 19848 22010
rect 19784 21950 19788 22006
rect 19788 21950 19844 22006
rect 19844 21950 19848 22006
rect 19784 21946 19848 21950
rect 19864 22006 19928 22010
rect 19864 21950 19868 22006
rect 19868 21950 19924 22006
rect 19924 21950 19928 22006
rect 19864 21946 19928 21950
rect 50344 22006 50408 22010
rect 50344 21950 50348 22006
rect 50348 21950 50404 22006
rect 50404 21950 50408 22006
rect 50344 21946 50408 21950
rect 50424 22006 50488 22010
rect 50424 21950 50428 22006
rect 50428 21950 50484 22006
rect 50484 21950 50488 22006
rect 50424 21946 50488 21950
rect 50504 22006 50568 22010
rect 50504 21950 50508 22006
rect 50508 21950 50564 22006
rect 50564 21950 50568 22006
rect 50504 21946 50568 21950
rect 50584 22006 50648 22010
rect 50584 21950 50588 22006
rect 50588 21950 50644 22006
rect 50644 21950 50648 22006
rect 50584 21946 50648 21950
rect 4264 21340 4328 21344
rect 4264 21284 4268 21340
rect 4268 21284 4324 21340
rect 4324 21284 4328 21340
rect 4264 21280 4328 21284
rect 4344 21340 4408 21344
rect 4344 21284 4348 21340
rect 4348 21284 4404 21340
rect 4404 21284 4408 21340
rect 4344 21280 4408 21284
rect 4424 21340 4488 21344
rect 4424 21284 4428 21340
rect 4428 21284 4484 21340
rect 4484 21284 4488 21340
rect 4424 21280 4488 21284
rect 4504 21340 4568 21344
rect 4504 21284 4508 21340
rect 4508 21284 4564 21340
rect 4564 21284 4568 21340
rect 4504 21280 4568 21284
rect 34984 21340 35048 21344
rect 34984 21284 34988 21340
rect 34988 21284 35044 21340
rect 35044 21284 35048 21340
rect 34984 21280 35048 21284
rect 35064 21340 35128 21344
rect 35064 21284 35068 21340
rect 35068 21284 35124 21340
rect 35124 21284 35128 21340
rect 35064 21280 35128 21284
rect 35144 21340 35208 21344
rect 35144 21284 35148 21340
rect 35148 21284 35204 21340
rect 35204 21284 35208 21340
rect 35144 21280 35208 21284
rect 35224 21340 35288 21344
rect 35224 21284 35228 21340
rect 35228 21284 35284 21340
rect 35284 21284 35288 21340
rect 35224 21280 35288 21284
rect 19624 20674 19688 20678
rect 19624 20618 19628 20674
rect 19628 20618 19684 20674
rect 19684 20618 19688 20674
rect 19624 20614 19688 20618
rect 19704 20674 19768 20678
rect 19704 20618 19708 20674
rect 19708 20618 19764 20674
rect 19764 20618 19768 20674
rect 19704 20614 19768 20618
rect 19784 20674 19848 20678
rect 19784 20618 19788 20674
rect 19788 20618 19844 20674
rect 19844 20618 19848 20674
rect 19784 20614 19848 20618
rect 19864 20674 19928 20678
rect 19864 20618 19868 20674
rect 19868 20618 19924 20674
rect 19924 20618 19928 20674
rect 19864 20614 19928 20618
rect 50344 20674 50408 20678
rect 50344 20618 50348 20674
rect 50348 20618 50404 20674
rect 50404 20618 50408 20674
rect 50344 20614 50408 20618
rect 50424 20674 50488 20678
rect 50424 20618 50428 20674
rect 50428 20618 50484 20674
rect 50484 20618 50488 20674
rect 50424 20614 50488 20618
rect 50504 20674 50568 20678
rect 50504 20618 50508 20674
rect 50508 20618 50564 20674
rect 50564 20618 50568 20674
rect 50504 20614 50568 20618
rect 50584 20674 50648 20678
rect 50584 20618 50588 20674
rect 50588 20618 50644 20674
rect 50644 20618 50648 20674
rect 50584 20614 50648 20618
rect 4264 20008 4328 20012
rect 4264 19952 4268 20008
rect 4268 19952 4324 20008
rect 4324 19952 4328 20008
rect 4264 19948 4328 19952
rect 4344 20008 4408 20012
rect 4344 19952 4348 20008
rect 4348 19952 4404 20008
rect 4404 19952 4408 20008
rect 4344 19948 4408 19952
rect 4424 20008 4488 20012
rect 4424 19952 4428 20008
rect 4428 19952 4484 20008
rect 4484 19952 4488 20008
rect 4424 19948 4488 19952
rect 4504 20008 4568 20012
rect 4504 19952 4508 20008
rect 4508 19952 4564 20008
rect 4564 19952 4568 20008
rect 4504 19948 4568 19952
rect 34984 20008 35048 20012
rect 34984 19952 34988 20008
rect 34988 19952 35044 20008
rect 35044 19952 35048 20008
rect 34984 19948 35048 19952
rect 35064 20008 35128 20012
rect 35064 19952 35068 20008
rect 35068 19952 35124 20008
rect 35124 19952 35128 20008
rect 35064 19948 35128 19952
rect 35144 20008 35208 20012
rect 35144 19952 35148 20008
rect 35148 19952 35204 20008
rect 35204 19952 35208 20008
rect 35144 19948 35208 19952
rect 35224 20008 35288 20012
rect 35224 19952 35228 20008
rect 35228 19952 35284 20008
rect 35284 19952 35288 20008
rect 35224 19948 35288 19952
rect 19624 19342 19688 19346
rect 19624 19286 19628 19342
rect 19628 19286 19684 19342
rect 19684 19286 19688 19342
rect 19624 19282 19688 19286
rect 19704 19342 19768 19346
rect 19704 19286 19708 19342
rect 19708 19286 19764 19342
rect 19764 19286 19768 19342
rect 19704 19282 19768 19286
rect 19784 19342 19848 19346
rect 19784 19286 19788 19342
rect 19788 19286 19844 19342
rect 19844 19286 19848 19342
rect 19784 19282 19848 19286
rect 19864 19342 19928 19346
rect 19864 19286 19868 19342
rect 19868 19286 19924 19342
rect 19924 19286 19928 19342
rect 19864 19282 19928 19286
rect 50344 19342 50408 19346
rect 50344 19286 50348 19342
rect 50348 19286 50404 19342
rect 50404 19286 50408 19342
rect 50344 19282 50408 19286
rect 50424 19342 50488 19346
rect 50424 19286 50428 19342
rect 50428 19286 50484 19342
rect 50484 19286 50488 19342
rect 50424 19282 50488 19286
rect 50504 19342 50568 19346
rect 50504 19286 50508 19342
rect 50508 19286 50564 19342
rect 50564 19286 50568 19342
rect 50504 19282 50568 19286
rect 50584 19342 50648 19346
rect 50584 19286 50588 19342
rect 50588 19286 50644 19342
rect 50644 19286 50648 19342
rect 50584 19282 50648 19286
rect 4264 18676 4328 18680
rect 4264 18620 4268 18676
rect 4268 18620 4324 18676
rect 4324 18620 4328 18676
rect 4264 18616 4328 18620
rect 4344 18676 4408 18680
rect 4344 18620 4348 18676
rect 4348 18620 4404 18676
rect 4404 18620 4408 18676
rect 4344 18616 4408 18620
rect 4424 18676 4488 18680
rect 4424 18620 4428 18676
rect 4428 18620 4484 18676
rect 4484 18620 4488 18676
rect 4424 18616 4488 18620
rect 4504 18676 4568 18680
rect 4504 18620 4508 18676
rect 4508 18620 4564 18676
rect 4564 18620 4568 18676
rect 4504 18616 4568 18620
rect 34984 18676 35048 18680
rect 34984 18620 34988 18676
rect 34988 18620 35044 18676
rect 35044 18620 35048 18676
rect 34984 18616 35048 18620
rect 35064 18676 35128 18680
rect 35064 18620 35068 18676
rect 35068 18620 35124 18676
rect 35124 18620 35128 18676
rect 35064 18616 35128 18620
rect 35144 18676 35208 18680
rect 35144 18620 35148 18676
rect 35148 18620 35204 18676
rect 35204 18620 35208 18676
rect 35144 18616 35208 18620
rect 35224 18676 35288 18680
rect 35224 18620 35228 18676
rect 35228 18620 35284 18676
rect 35284 18620 35288 18676
rect 35224 18616 35288 18620
rect 19624 18010 19688 18014
rect 19624 17954 19628 18010
rect 19628 17954 19684 18010
rect 19684 17954 19688 18010
rect 19624 17950 19688 17954
rect 19704 18010 19768 18014
rect 19704 17954 19708 18010
rect 19708 17954 19764 18010
rect 19764 17954 19768 18010
rect 19704 17950 19768 17954
rect 19784 18010 19848 18014
rect 19784 17954 19788 18010
rect 19788 17954 19844 18010
rect 19844 17954 19848 18010
rect 19784 17950 19848 17954
rect 19864 18010 19928 18014
rect 19864 17954 19868 18010
rect 19868 17954 19924 18010
rect 19924 17954 19928 18010
rect 19864 17950 19928 17954
rect 50344 18010 50408 18014
rect 50344 17954 50348 18010
rect 50348 17954 50404 18010
rect 50404 17954 50408 18010
rect 50344 17950 50408 17954
rect 50424 18010 50488 18014
rect 50424 17954 50428 18010
rect 50428 17954 50484 18010
rect 50484 17954 50488 18010
rect 50424 17950 50488 17954
rect 50504 18010 50568 18014
rect 50504 17954 50508 18010
rect 50508 17954 50564 18010
rect 50564 17954 50568 18010
rect 50504 17950 50568 17954
rect 50584 18010 50648 18014
rect 50584 17954 50588 18010
rect 50588 17954 50644 18010
rect 50644 17954 50648 18010
rect 50584 17950 50648 17954
rect 4264 17344 4328 17348
rect 4264 17288 4268 17344
rect 4268 17288 4324 17344
rect 4324 17288 4328 17344
rect 4264 17284 4328 17288
rect 4344 17344 4408 17348
rect 4344 17288 4348 17344
rect 4348 17288 4404 17344
rect 4404 17288 4408 17344
rect 4344 17284 4408 17288
rect 4424 17344 4488 17348
rect 4424 17288 4428 17344
rect 4428 17288 4484 17344
rect 4484 17288 4488 17344
rect 4424 17284 4488 17288
rect 4504 17344 4568 17348
rect 4504 17288 4508 17344
rect 4508 17288 4564 17344
rect 4564 17288 4568 17344
rect 4504 17284 4568 17288
rect 34984 17344 35048 17348
rect 34984 17288 34988 17344
rect 34988 17288 35044 17344
rect 35044 17288 35048 17344
rect 34984 17284 35048 17288
rect 35064 17344 35128 17348
rect 35064 17288 35068 17344
rect 35068 17288 35124 17344
rect 35124 17288 35128 17344
rect 35064 17284 35128 17288
rect 35144 17344 35208 17348
rect 35144 17288 35148 17344
rect 35148 17288 35204 17344
rect 35204 17288 35208 17344
rect 35144 17284 35208 17288
rect 35224 17344 35288 17348
rect 35224 17288 35228 17344
rect 35228 17288 35284 17344
rect 35284 17288 35288 17344
rect 35224 17284 35288 17288
rect 19624 16678 19688 16682
rect 19624 16622 19628 16678
rect 19628 16622 19684 16678
rect 19684 16622 19688 16678
rect 19624 16618 19688 16622
rect 19704 16678 19768 16682
rect 19704 16622 19708 16678
rect 19708 16622 19764 16678
rect 19764 16622 19768 16678
rect 19704 16618 19768 16622
rect 19784 16678 19848 16682
rect 19784 16622 19788 16678
rect 19788 16622 19844 16678
rect 19844 16622 19848 16678
rect 19784 16618 19848 16622
rect 19864 16678 19928 16682
rect 19864 16622 19868 16678
rect 19868 16622 19924 16678
rect 19924 16622 19928 16678
rect 19864 16618 19928 16622
rect 50344 16678 50408 16682
rect 50344 16622 50348 16678
rect 50348 16622 50404 16678
rect 50404 16622 50408 16678
rect 50344 16618 50408 16622
rect 50424 16678 50488 16682
rect 50424 16622 50428 16678
rect 50428 16622 50484 16678
rect 50484 16622 50488 16678
rect 50424 16618 50488 16622
rect 50504 16678 50568 16682
rect 50504 16622 50508 16678
rect 50508 16622 50564 16678
rect 50564 16622 50568 16678
rect 50504 16618 50568 16622
rect 50584 16678 50648 16682
rect 50584 16622 50588 16678
rect 50588 16622 50644 16678
rect 50644 16622 50648 16678
rect 50584 16618 50648 16622
rect 4264 16012 4328 16016
rect 4264 15956 4268 16012
rect 4268 15956 4324 16012
rect 4324 15956 4328 16012
rect 4264 15952 4328 15956
rect 4344 16012 4408 16016
rect 4344 15956 4348 16012
rect 4348 15956 4404 16012
rect 4404 15956 4408 16012
rect 4344 15952 4408 15956
rect 4424 16012 4488 16016
rect 4424 15956 4428 16012
rect 4428 15956 4484 16012
rect 4484 15956 4488 16012
rect 4424 15952 4488 15956
rect 4504 16012 4568 16016
rect 4504 15956 4508 16012
rect 4508 15956 4564 16012
rect 4564 15956 4568 16012
rect 4504 15952 4568 15956
rect 34984 16012 35048 16016
rect 34984 15956 34988 16012
rect 34988 15956 35044 16012
rect 35044 15956 35048 16012
rect 34984 15952 35048 15956
rect 35064 16012 35128 16016
rect 35064 15956 35068 16012
rect 35068 15956 35124 16012
rect 35124 15956 35128 16012
rect 35064 15952 35128 15956
rect 35144 16012 35208 16016
rect 35144 15956 35148 16012
rect 35148 15956 35204 16012
rect 35204 15956 35208 16012
rect 35144 15952 35208 15956
rect 35224 16012 35288 16016
rect 35224 15956 35228 16012
rect 35228 15956 35284 16012
rect 35284 15956 35288 16012
rect 35224 15952 35288 15956
rect 19624 15346 19688 15350
rect 19624 15290 19628 15346
rect 19628 15290 19684 15346
rect 19684 15290 19688 15346
rect 19624 15286 19688 15290
rect 19704 15346 19768 15350
rect 19704 15290 19708 15346
rect 19708 15290 19764 15346
rect 19764 15290 19768 15346
rect 19704 15286 19768 15290
rect 19784 15346 19848 15350
rect 19784 15290 19788 15346
rect 19788 15290 19844 15346
rect 19844 15290 19848 15346
rect 19784 15286 19848 15290
rect 19864 15346 19928 15350
rect 19864 15290 19868 15346
rect 19868 15290 19924 15346
rect 19924 15290 19928 15346
rect 19864 15286 19928 15290
rect 50344 15346 50408 15350
rect 50344 15290 50348 15346
rect 50348 15290 50404 15346
rect 50404 15290 50408 15346
rect 50344 15286 50408 15290
rect 50424 15346 50488 15350
rect 50424 15290 50428 15346
rect 50428 15290 50484 15346
rect 50484 15290 50488 15346
rect 50424 15286 50488 15290
rect 50504 15346 50568 15350
rect 50504 15290 50508 15346
rect 50508 15290 50564 15346
rect 50564 15290 50568 15346
rect 50504 15286 50568 15290
rect 50584 15346 50648 15350
rect 50584 15290 50588 15346
rect 50588 15290 50644 15346
rect 50644 15290 50648 15346
rect 50584 15286 50648 15290
rect 4264 14680 4328 14684
rect 4264 14624 4268 14680
rect 4268 14624 4324 14680
rect 4324 14624 4328 14680
rect 4264 14620 4328 14624
rect 4344 14680 4408 14684
rect 4344 14624 4348 14680
rect 4348 14624 4404 14680
rect 4404 14624 4408 14680
rect 4344 14620 4408 14624
rect 4424 14680 4488 14684
rect 4424 14624 4428 14680
rect 4428 14624 4484 14680
rect 4484 14624 4488 14680
rect 4424 14620 4488 14624
rect 4504 14680 4568 14684
rect 4504 14624 4508 14680
rect 4508 14624 4564 14680
rect 4564 14624 4568 14680
rect 4504 14620 4568 14624
rect 34984 14680 35048 14684
rect 34984 14624 34988 14680
rect 34988 14624 35044 14680
rect 35044 14624 35048 14680
rect 34984 14620 35048 14624
rect 35064 14680 35128 14684
rect 35064 14624 35068 14680
rect 35068 14624 35124 14680
rect 35124 14624 35128 14680
rect 35064 14620 35128 14624
rect 35144 14680 35208 14684
rect 35144 14624 35148 14680
rect 35148 14624 35204 14680
rect 35204 14624 35208 14680
rect 35144 14620 35208 14624
rect 35224 14680 35288 14684
rect 35224 14624 35228 14680
rect 35228 14624 35284 14680
rect 35284 14624 35288 14680
rect 35224 14620 35288 14624
rect 19624 14014 19688 14018
rect 19624 13958 19628 14014
rect 19628 13958 19684 14014
rect 19684 13958 19688 14014
rect 19624 13954 19688 13958
rect 19704 14014 19768 14018
rect 19704 13958 19708 14014
rect 19708 13958 19764 14014
rect 19764 13958 19768 14014
rect 19704 13954 19768 13958
rect 19784 14014 19848 14018
rect 19784 13958 19788 14014
rect 19788 13958 19844 14014
rect 19844 13958 19848 14014
rect 19784 13954 19848 13958
rect 19864 14014 19928 14018
rect 19864 13958 19868 14014
rect 19868 13958 19924 14014
rect 19924 13958 19928 14014
rect 19864 13954 19928 13958
rect 50344 14014 50408 14018
rect 50344 13958 50348 14014
rect 50348 13958 50404 14014
rect 50404 13958 50408 14014
rect 50344 13954 50408 13958
rect 50424 14014 50488 14018
rect 50424 13958 50428 14014
rect 50428 13958 50484 14014
rect 50484 13958 50488 14014
rect 50424 13954 50488 13958
rect 50504 14014 50568 14018
rect 50504 13958 50508 14014
rect 50508 13958 50564 14014
rect 50564 13958 50568 14014
rect 50504 13954 50568 13958
rect 50584 14014 50648 14018
rect 50584 13958 50588 14014
rect 50588 13958 50644 14014
rect 50644 13958 50648 14014
rect 50584 13954 50648 13958
rect 4264 13348 4328 13352
rect 4264 13292 4268 13348
rect 4268 13292 4324 13348
rect 4324 13292 4328 13348
rect 4264 13288 4328 13292
rect 4344 13348 4408 13352
rect 4344 13292 4348 13348
rect 4348 13292 4404 13348
rect 4404 13292 4408 13348
rect 4344 13288 4408 13292
rect 4424 13348 4488 13352
rect 4424 13292 4428 13348
rect 4428 13292 4484 13348
rect 4484 13292 4488 13348
rect 4424 13288 4488 13292
rect 4504 13348 4568 13352
rect 4504 13292 4508 13348
rect 4508 13292 4564 13348
rect 4564 13292 4568 13348
rect 4504 13288 4568 13292
rect 34984 13348 35048 13352
rect 34984 13292 34988 13348
rect 34988 13292 35044 13348
rect 35044 13292 35048 13348
rect 34984 13288 35048 13292
rect 35064 13348 35128 13352
rect 35064 13292 35068 13348
rect 35068 13292 35124 13348
rect 35124 13292 35128 13348
rect 35064 13288 35128 13292
rect 35144 13348 35208 13352
rect 35144 13292 35148 13348
rect 35148 13292 35204 13348
rect 35204 13292 35208 13348
rect 35144 13288 35208 13292
rect 35224 13348 35288 13352
rect 35224 13292 35228 13348
rect 35228 13292 35284 13348
rect 35284 13292 35288 13348
rect 35224 13288 35288 13292
rect 19624 12682 19688 12686
rect 19624 12626 19628 12682
rect 19628 12626 19684 12682
rect 19684 12626 19688 12682
rect 19624 12622 19688 12626
rect 19704 12682 19768 12686
rect 19704 12626 19708 12682
rect 19708 12626 19764 12682
rect 19764 12626 19768 12682
rect 19704 12622 19768 12626
rect 19784 12682 19848 12686
rect 19784 12626 19788 12682
rect 19788 12626 19844 12682
rect 19844 12626 19848 12682
rect 19784 12622 19848 12626
rect 19864 12682 19928 12686
rect 19864 12626 19868 12682
rect 19868 12626 19924 12682
rect 19924 12626 19928 12682
rect 19864 12622 19928 12626
rect 50344 12682 50408 12686
rect 50344 12626 50348 12682
rect 50348 12626 50404 12682
rect 50404 12626 50408 12682
rect 50344 12622 50408 12626
rect 50424 12682 50488 12686
rect 50424 12626 50428 12682
rect 50428 12626 50484 12682
rect 50484 12626 50488 12682
rect 50424 12622 50488 12626
rect 50504 12682 50568 12686
rect 50504 12626 50508 12682
rect 50508 12626 50564 12682
rect 50564 12626 50568 12682
rect 50504 12622 50568 12626
rect 50584 12682 50648 12686
rect 50584 12626 50588 12682
rect 50588 12626 50644 12682
rect 50644 12626 50648 12682
rect 50584 12622 50648 12626
rect 4264 12016 4328 12020
rect 4264 11960 4268 12016
rect 4268 11960 4324 12016
rect 4324 11960 4328 12016
rect 4264 11956 4328 11960
rect 4344 12016 4408 12020
rect 4344 11960 4348 12016
rect 4348 11960 4404 12016
rect 4404 11960 4408 12016
rect 4344 11956 4408 11960
rect 4424 12016 4488 12020
rect 4424 11960 4428 12016
rect 4428 11960 4484 12016
rect 4484 11960 4488 12016
rect 4424 11956 4488 11960
rect 4504 12016 4568 12020
rect 4504 11960 4508 12016
rect 4508 11960 4564 12016
rect 4564 11960 4568 12016
rect 4504 11956 4568 11960
rect 34984 12016 35048 12020
rect 34984 11960 34988 12016
rect 34988 11960 35044 12016
rect 35044 11960 35048 12016
rect 34984 11956 35048 11960
rect 35064 12016 35128 12020
rect 35064 11960 35068 12016
rect 35068 11960 35124 12016
rect 35124 11960 35128 12016
rect 35064 11956 35128 11960
rect 35144 12016 35208 12020
rect 35144 11960 35148 12016
rect 35148 11960 35204 12016
rect 35204 11960 35208 12016
rect 35144 11956 35208 11960
rect 35224 12016 35288 12020
rect 35224 11960 35228 12016
rect 35228 11960 35284 12016
rect 35284 11960 35288 12016
rect 35224 11956 35288 11960
rect 19624 11350 19688 11354
rect 19624 11294 19628 11350
rect 19628 11294 19684 11350
rect 19684 11294 19688 11350
rect 19624 11290 19688 11294
rect 19704 11350 19768 11354
rect 19704 11294 19708 11350
rect 19708 11294 19764 11350
rect 19764 11294 19768 11350
rect 19704 11290 19768 11294
rect 19784 11350 19848 11354
rect 19784 11294 19788 11350
rect 19788 11294 19844 11350
rect 19844 11294 19848 11350
rect 19784 11290 19848 11294
rect 19864 11350 19928 11354
rect 19864 11294 19868 11350
rect 19868 11294 19924 11350
rect 19924 11294 19928 11350
rect 19864 11290 19928 11294
rect 50344 11350 50408 11354
rect 50344 11294 50348 11350
rect 50348 11294 50404 11350
rect 50404 11294 50408 11350
rect 50344 11290 50408 11294
rect 50424 11350 50488 11354
rect 50424 11294 50428 11350
rect 50428 11294 50484 11350
rect 50484 11294 50488 11350
rect 50424 11290 50488 11294
rect 50504 11350 50568 11354
rect 50504 11294 50508 11350
rect 50508 11294 50564 11350
rect 50564 11294 50568 11350
rect 50504 11290 50568 11294
rect 50584 11350 50648 11354
rect 50584 11294 50588 11350
rect 50588 11294 50644 11350
rect 50644 11294 50648 11350
rect 50584 11290 50648 11294
rect 4264 10684 4328 10688
rect 4264 10628 4268 10684
rect 4268 10628 4324 10684
rect 4324 10628 4328 10684
rect 4264 10624 4328 10628
rect 4344 10684 4408 10688
rect 4344 10628 4348 10684
rect 4348 10628 4404 10684
rect 4404 10628 4408 10684
rect 4344 10624 4408 10628
rect 4424 10684 4488 10688
rect 4424 10628 4428 10684
rect 4428 10628 4484 10684
rect 4484 10628 4488 10684
rect 4424 10624 4488 10628
rect 4504 10684 4568 10688
rect 4504 10628 4508 10684
rect 4508 10628 4564 10684
rect 4564 10628 4568 10684
rect 4504 10624 4568 10628
rect 34984 10684 35048 10688
rect 34984 10628 34988 10684
rect 34988 10628 35044 10684
rect 35044 10628 35048 10684
rect 34984 10624 35048 10628
rect 35064 10684 35128 10688
rect 35064 10628 35068 10684
rect 35068 10628 35124 10684
rect 35124 10628 35128 10684
rect 35064 10624 35128 10628
rect 35144 10684 35208 10688
rect 35144 10628 35148 10684
rect 35148 10628 35204 10684
rect 35204 10628 35208 10684
rect 35144 10624 35208 10628
rect 35224 10684 35288 10688
rect 35224 10628 35228 10684
rect 35228 10628 35284 10684
rect 35284 10628 35288 10684
rect 35224 10624 35288 10628
rect 19624 10018 19688 10022
rect 19624 9962 19628 10018
rect 19628 9962 19684 10018
rect 19684 9962 19688 10018
rect 19624 9958 19688 9962
rect 19704 10018 19768 10022
rect 19704 9962 19708 10018
rect 19708 9962 19764 10018
rect 19764 9962 19768 10018
rect 19704 9958 19768 9962
rect 19784 10018 19848 10022
rect 19784 9962 19788 10018
rect 19788 9962 19844 10018
rect 19844 9962 19848 10018
rect 19784 9958 19848 9962
rect 19864 10018 19928 10022
rect 19864 9962 19868 10018
rect 19868 9962 19924 10018
rect 19924 9962 19928 10018
rect 19864 9958 19928 9962
rect 50344 10018 50408 10022
rect 50344 9962 50348 10018
rect 50348 9962 50404 10018
rect 50404 9962 50408 10018
rect 50344 9958 50408 9962
rect 50424 10018 50488 10022
rect 50424 9962 50428 10018
rect 50428 9962 50484 10018
rect 50484 9962 50488 10018
rect 50424 9958 50488 9962
rect 50504 10018 50568 10022
rect 50504 9962 50508 10018
rect 50508 9962 50564 10018
rect 50564 9962 50568 10018
rect 50504 9958 50568 9962
rect 50584 10018 50648 10022
rect 50584 9962 50588 10018
rect 50588 9962 50644 10018
rect 50644 9962 50648 10018
rect 50584 9958 50648 9962
rect 4264 9352 4328 9356
rect 4264 9296 4268 9352
rect 4268 9296 4324 9352
rect 4324 9296 4328 9352
rect 4264 9292 4328 9296
rect 4344 9352 4408 9356
rect 4344 9296 4348 9352
rect 4348 9296 4404 9352
rect 4404 9296 4408 9352
rect 4344 9292 4408 9296
rect 4424 9352 4488 9356
rect 4424 9296 4428 9352
rect 4428 9296 4484 9352
rect 4484 9296 4488 9352
rect 4424 9292 4488 9296
rect 4504 9352 4568 9356
rect 4504 9296 4508 9352
rect 4508 9296 4564 9352
rect 4564 9296 4568 9352
rect 4504 9292 4568 9296
rect 34984 9352 35048 9356
rect 34984 9296 34988 9352
rect 34988 9296 35044 9352
rect 35044 9296 35048 9352
rect 34984 9292 35048 9296
rect 35064 9352 35128 9356
rect 35064 9296 35068 9352
rect 35068 9296 35124 9352
rect 35124 9296 35128 9352
rect 35064 9292 35128 9296
rect 35144 9352 35208 9356
rect 35144 9296 35148 9352
rect 35148 9296 35204 9352
rect 35204 9296 35208 9352
rect 35144 9292 35208 9296
rect 35224 9352 35288 9356
rect 35224 9296 35228 9352
rect 35228 9296 35284 9352
rect 35284 9296 35288 9352
rect 35224 9292 35288 9296
rect 10048 9070 10112 9134
rect 19624 8686 19688 8690
rect 19624 8630 19628 8686
rect 19628 8630 19684 8686
rect 19684 8630 19688 8686
rect 19624 8626 19688 8630
rect 19704 8686 19768 8690
rect 19704 8630 19708 8686
rect 19708 8630 19764 8686
rect 19764 8630 19768 8686
rect 19704 8626 19768 8630
rect 19784 8686 19848 8690
rect 19784 8630 19788 8686
rect 19788 8630 19844 8686
rect 19844 8630 19848 8686
rect 19784 8626 19848 8630
rect 19864 8686 19928 8690
rect 19864 8630 19868 8686
rect 19868 8630 19924 8686
rect 19924 8630 19928 8686
rect 19864 8626 19928 8630
rect 50344 8686 50408 8690
rect 50344 8630 50348 8686
rect 50348 8630 50404 8686
rect 50404 8630 50408 8686
rect 50344 8626 50408 8630
rect 50424 8686 50488 8690
rect 50424 8630 50428 8686
rect 50428 8630 50484 8686
rect 50484 8630 50488 8686
rect 50424 8626 50488 8630
rect 50504 8686 50568 8690
rect 50504 8630 50508 8686
rect 50508 8630 50564 8686
rect 50564 8630 50568 8686
rect 50504 8626 50568 8630
rect 50584 8686 50648 8690
rect 50584 8630 50588 8686
rect 50588 8630 50644 8686
rect 50644 8630 50648 8686
rect 50584 8626 50648 8630
rect 4264 8020 4328 8024
rect 4264 7964 4268 8020
rect 4268 7964 4324 8020
rect 4324 7964 4328 8020
rect 4264 7960 4328 7964
rect 4344 8020 4408 8024
rect 4344 7964 4348 8020
rect 4348 7964 4404 8020
rect 4404 7964 4408 8020
rect 4344 7960 4408 7964
rect 4424 8020 4488 8024
rect 4424 7964 4428 8020
rect 4428 7964 4484 8020
rect 4484 7964 4488 8020
rect 4424 7960 4488 7964
rect 4504 8020 4568 8024
rect 4504 7964 4508 8020
rect 4508 7964 4564 8020
rect 4564 7964 4568 8020
rect 4504 7960 4568 7964
rect 34984 8020 35048 8024
rect 34984 7964 34988 8020
rect 34988 7964 35044 8020
rect 35044 7964 35048 8020
rect 34984 7960 35048 7964
rect 35064 8020 35128 8024
rect 35064 7964 35068 8020
rect 35068 7964 35124 8020
rect 35124 7964 35128 8020
rect 35064 7960 35128 7964
rect 35144 8020 35208 8024
rect 35144 7964 35148 8020
rect 35148 7964 35204 8020
rect 35204 7964 35208 8020
rect 35144 7960 35208 7964
rect 35224 8020 35288 8024
rect 35224 7964 35228 8020
rect 35228 7964 35284 8020
rect 35284 7964 35288 8020
rect 35224 7960 35288 7964
rect 9856 7502 9920 7506
rect 9856 7446 9908 7502
rect 9908 7446 9920 7502
rect 9856 7442 9920 7446
rect 19624 7354 19688 7358
rect 19624 7298 19628 7354
rect 19628 7298 19684 7354
rect 19684 7298 19688 7354
rect 19624 7294 19688 7298
rect 19704 7354 19768 7358
rect 19704 7298 19708 7354
rect 19708 7298 19764 7354
rect 19764 7298 19768 7354
rect 19704 7294 19768 7298
rect 19784 7354 19848 7358
rect 19784 7298 19788 7354
rect 19788 7298 19844 7354
rect 19844 7298 19848 7354
rect 19784 7294 19848 7298
rect 19864 7354 19928 7358
rect 19864 7298 19868 7354
rect 19868 7298 19924 7354
rect 19924 7298 19928 7354
rect 19864 7294 19928 7298
rect 50344 7354 50408 7358
rect 50344 7298 50348 7354
rect 50348 7298 50404 7354
rect 50404 7298 50408 7354
rect 50344 7294 50408 7298
rect 50424 7354 50488 7358
rect 50424 7298 50428 7354
rect 50428 7298 50484 7354
rect 50484 7298 50488 7354
rect 50424 7294 50488 7298
rect 50504 7354 50568 7358
rect 50504 7298 50508 7354
rect 50508 7298 50564 7354
rect 50564 7298 50568 7354
rect 50504 7294 50568 7298
rect 50584 7354 50648 7358
rect 50584 7298 50588 7354
rect 50588 7298 50644 7354
rect 50644 7298 50648 7354
rect 50584 7294 50648 7298
rect 29056 6702 29120 6766
rect 4264 6688 4328 6692
rect 4264 6632 4268 6688
rect 4268 6632 4324 6688
rect 4324 6632 4328 6688
rect 4264 6628 4328 6632
rect 4344 6688 4408 6692
rect 4344 6632 4348 6688
rect 4348 6632 4404 6688
rect 4404 6632 4408 6688
rect 4344 6628 4408 6632
rect 4424 6688 4488 6692
rect 4424 6632 4428 6688
rect 4428 6632 4484 6688
rect 4484 6632 4488 6688
rect 4424 6628 4488 6632
rect 4504 6688 4568 6692
rect 4504 6632 4508 6688
rect 4508 6632 4564 6688
rect 4564 6632 4568 6688
rect 4504 6628 4568 6632
rect 34984 6688 35048 6692
rect 34984 6632 34988 6688
rect 34988 6632 35044 6688
rect 35044 6632 35048 6688
rect 34984 6628 35048 6632
rect 35064 6688 35128 6692
rect 35064 6632 35068 6688
rect 35068 6632 35124 6688
rect 35124 6632 35128 6688
rect 35064 6628 35128 6632
rect 35144 6688 35208 6692
rect 35144 6632 35148 6688
rect 35148 6632 35204 6688
rect 35204 6632 35208 6688
rect 35144 6628 35208 6632
rect 35224 6688 35288 6692
rect 35224 6632 35228 6688
rect 35228 6632 35284 6688
rect 35284 6632 35288 6688
rect 35224 6628 35288 6632
rect 28288 6554 28352 6618
rect 19624 6022 19688 6026
rect 19624 5966 19628 6022
rect 19628 5966 19684 6022
rect 19684 5966 19688 6022
rect 19624 5962 19688 5966
rect 19704 6022 19768 6026
rect 19704 5966 19708 6022
rect 19708 5966 19764 6022
rect 19764 5966 19768 6022
rect 19704 5962 19768 5966
rect 19784 6022 19848 6026
rect 19784 5966 19788 6022
rect 19788 5966 19844 6022
rect 19844 5966 19848 6022
rect 19784 5962 19848 5966
rect 19864 6022 19928 6026
rect 19864 5966 19868 6022
rect 19868 5966 19924 6022
rect 19924 5966 19928 6022
rect 19864 5962 19928 5966
rect 50344 6022 50408 6026
rect 50344 5966 50348 6022
rect 50348 5966 50404 6022
rect 50404 5966 50408 6022
rect 50344 5962 50408 5966
rect 50424 6022 50488 6026
rect 50424 5966 50428 6022
rect 50428 5966 50484 6022
rect 50484 5966 50488 6022
rect 50424 5962 50488 5966
rect 50504 6022 50568 6026
rect 50504 5966 50508 6022
rect 50508 5966 50564 6022
rect 50564 5966 50568 6022
rect 50504 5962 50568 5966
rect 50584 6022 50648 6026
rect 50584 5966 50588 6022
rect 50588 5966 50644 6022
rect 50644 5966 50648 6022
rect 50584 5962 50648 5966
rect 4264 5356 4328 5360
rect 4264 5300 4268 5356
rect 4268 5300 4324 5356
rect 4324 5300 4328 5356
rect 4264 5296 4328 5300
rect 4344 5356 4408 5360
rect 4344 5300 4348 5356
rect 4348 5300 4404 5356
rect 4404 5300 4408 5356
rect 4344 5296 4408 5300
rect 4424 5356 4488 5360
rect 4424 5300 4428 5356
rect 4428 5300 4484 5356
rect 4484 5300 4488 5356
rect 4424 5296 4488 5300
rect 4504 5356 4568 5360
rect 4504 5300 4508 5356
rect 4508 5300 4564 5356
rect 4564 5300 4568 5356
rect 4504 5296 4568 5300
rect 34984 5356 35048 5360
rect 34984 5300 34988 5356
rect 34988 5300 35044 5356
rect 35044 5300 35048 5356
rect 34984 5296 35048 5300
rect 35064 5356 35128 5360
rect 35064 5300 35068 5356
rect 35068 5300 35124 5356
rect 35124 5300 35128 5356
rect 35064 5296 35128 5300
rect 35144 5356 35208 5360
rect 35144 5300 35148 5356
rect 35148 5300 35204 5356
rect 35204 5300 35208 5356
rect 35144 5296 35208 5300
rect 35224 5356 35288 5360
rect 35224 5300 35228 5356
rect 35228 5300 35284 5356
rect 35284 5300 35288 5356
rect 35224 5296 35288 5300
rect 19624 4690 19688 4694
rect 19624 4634 19628 4690
rect 19628 4634 19684 4690
rect 19684 4634 19688 4690
rect 19624 4630 19688 4634
rect 19704 4690 19768 4694
rect 19704 4634 19708 4690
rect 19708 4634 19764 4690
rect 19764 4634 19768 4690
rect 19704 4630 19768 4634
rect 19784 4690 19848 4694
rect 19784 4634 19788 4690
rect 19788 4634 19844 4690
rect 19844 4634 19848 4690
rect 19784 4630 19848 4634
rect 19864 4690 19928 4694
rect 19864 4634 19868 4690
rect 19868 4634 19924 4690
rect 19924 4634 19928 4690
rect 19864 4630 19928 4634
rect 50344 4690 50408 4694
rect 50344 4634 50348 4690
rect 50348 4634 50404 4690
rect 50404 4634 50408 4690
rect 50344 4630 50408 4634
rect 50424 4690 50488 4694
rect 50424 4634 50428 4690
rect 50428 4634 50484 4690
rect 50484 4634 50488 4690
rect 50424 4630 50488 4634
rect 50504 4690 50568 4694
rect 50504 4634 50508 4690
rect 50508 4634 50564 4690
rect 50564 4634 50568 4690
rect 50504 4630 50568 4634
rect 50584 4690 50648 4694
rect 50584 4634 50588 4690
rect 50588 4634 50644 4690
rect 50644 4634 50648 4690
rect 50584 4630 50648 4634
rect 4264 4024 4328 4028
rect 4264 3968 4268 4024
rect 4268 3968 4324 4024
rect 4324 3968 4328 4024
rect 4264 3964 4328 3968
rect 4344 4024 4408 4028
rect 4344 3968 4348 4024
rect 4348 3968 4404 4024
rect 4404 3968 4408 4024
rect 4344 3964 4408 3968
rect 4424 4024 4488 4028
rect 4424 3968 4428 4024
rect 4428 3968 4484 4024
rect 4484 3968 4488 4024
rect 4424 3964 4488 3968
rect 4504 4024 4568 4028
rect 4504 3968 4508 4024
rect 4508 3968 4564 4024
rect 4564 3968 4568 4024
rect 4504 3964 4568 3968
rect 34984 4024 35048 4028
rect 34984 3968 34988 4024
rect 34988 3968 35044 4024
rect 35044 3968 35048 4024
rect 34984 3964 35048 3968
rect 35064 4024 35128 4028
rect 35064 3968 35068 4024
rect 35068 3968 35124 4024
rect 35124 3968 35128 4024
rect 35064 3964 35128 3968
rect 35144 4024 35208 4028
rect 35144 3968 35148 4024
rect 35148 3968 35204 4024
rect 35204 3968 35208 4024
rect 35144 3964 35208 3968
rect 35224 4024 35288 4028
rect 35224 3968 35228 4024
rect 35228 3968 35284 4024
rect 35284 3968 35288 4024
rect 35224 3964 35288 3968
rect 9856 3950 9920 3954
rect 9856 3894 9908 3950
rect 9908 3894 9920 3950
rect 9856 3890 9920 3894
rect 10048 3594 10112 3658
rect 19624 3358 19688 3362
rect 19624 3302 19628 3358
rect 19628 3302 19684 3358
rect 19684 3302 19688 3358
rect 19624 3298 19688 3302
rect 19704 3358 19768 3362
rect 19704 3302 19708 3358
rect 19708 3302 19764 3358
rect 19764 3302 19768 3358
rect 19704 3298 19768 3302
rect 19784 3358 19848 3362
rect 19784 3302 19788 3358
rect 19788 3302 19844 3358
rect 19844 3302 19848 3358
rect 19784 3298 19848 3302
rect 19864 3358 19928 3362
rect 19864 3302 19868 3358
rect 19868 3302 19924 3358
rect 19924 3302 19928 3358
rect 19864 3298 19928 3302
rect 50344 3358 50408 3362
rect 50344 3302 50348 3358
rect 50348 3302 50404 3358
rect 50404 3302 50408 3358
rect 50344 3298 50408 3302
rect 50424 3358 50488 3362
rect 50424 3302 50428 3358
rect 50428 3302 50484 3358
rect 50484 3302 50488 3358
rect 50424 3298 50488 3302
rect 50504 3358 50568 3362
rect 50504 3302 50508 3358
rect 50508 3302 50564 3358
rect 50564 3302 50568 3358
rect 50504 3298 50568 3302
rect 50584 3358 50648 3362
rect 50584 3302 50588 3358
rect 50588 3302 50644 3358
rect 50644 3302 50648 3358
rect 50584 3298 50648 3302
rect 8320 3150 8384 3214
rect 7360 3002 7424 3066
rect 8128 2854 8192 2918
rect 4264 2692 4328 2696
rect 4264 2636 4268 2692
rect 4268 2636 4324 2692
rect 4324 2636 4328 2692
rect 4264 2632 4328 2636
rect 4344 2692 4408 2696
rect 4344 2636 4348 2692
rect 4348 2636 4404 2692
rect 4404 2636 4408 2692
rect 4344 2632 4408 2636
rect 4424 2692 4488 2696
rect 4424 2636 4428 2692
rect 4428 2636 4484 2692
rect 4484 2636 4488 2692
rect 4424 2632 4488 2636
rect 4504 2692 4568 2696
rect 4504 2636 4508 2692
rect 4508 2636 4564 2692
rect 4564 2636 4568 2692
rect 4504 2632 4568 2636
rect 34984 2692 35048 2696
rect 34984 2636 34988 2692
rect 34988 2636 35044 2692
rect 35044 2636 35048 2692
rect 34984 2632 35048 2636
rect 35064 2692 35128 2696
rect 35064 2636 35068 2692
rect 35068 2636 35124 2692
rect 35124 2636 35128 2692
rect 35064 2632 35128 2636
rect 35144 2692 35208 2696
rect 35144 2636 35148 2692
rect 35148 2636 35204 2692
rect 35204 2636 35208 2692
rect 35144 2632 35208 2636
rect 35224 2692 35288 2696
rect 35224 2636 35228 2692
rect 35228 2636 35284 2692
rect 35284 2636 35288 2692
rect 35224 2632 35288 2636
<< metal4 >>
rect 4256 57308 4576 57324
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 55976 4576 57244
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 54644 4576 55912
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 53312 4576 54580
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 51980 4576 53248
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 50648 4576 51916
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 49316 4576 50584
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 47984 4576 49252
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 46652 4576 47920
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 45320 4576 46588
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 43988 4576 45256
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 42656 4576 43924
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 41324 4576 42592
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 39992 4576 41260
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 38660 4576 39928
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 37328 4576 38596
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 35996 4576 37264
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 34664 4576 35932
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 33332 4576 34600
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 32000 4576 33268
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 30668 4576 31936
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 29336 4576 30604
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 28004 4576 29272
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 26672 4576 27940
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 25340 4576 26608
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 24008 4576 25276
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 22676 4576 23944
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 21344 4576 22612
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 20012 4576 21280
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 18680 4576 19948
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 17348 4576 18616
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 16016 4576 17284
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 14684 4576 15952
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 13352 4576 14620
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 12020 4576 13288
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 10688 4576 11956
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 9356 4576 10624
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 8024 4576 9292
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 6692 4576 7960
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 5360 4576 6628
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 4028 4576 5296
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 2696 4576 3964
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4916 2664 5236 57276
rect 5576 2664 5896 57276
rect 6236 2664 6556 57276
rect 19616 56642 19936 57324
rect 34976 57308 35296 57324
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 7359 56198 7425 56199
rect 7359 56134 7360 56198
rect 7424 56134 7425 56198
rect 7359 56133 7425 56134
rect 7362 3067 7422 56133
rect 19616 55310 19936 56578
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 53978 19936 55246
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 52646 19936 53914
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 51314 19936 52582
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 49982 19936 51250
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 48650 19936 49918
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 47318 19936 48586
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 45986 19936 47254
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 44654 19936 45922
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 43322 19936 44590
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 41990 19936 43258
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 40658 19936 41926
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 39326 19936 40594
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 37994 19936 39262
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 36662 19936 37930
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 35330 19936 36598
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 33998 19936 35266
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 32666 19936 33934
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 31334 19936 32602
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 30002 19936 31270
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 8127 28966 8193 28967
rect 8127 28902 8128 28966
rect 8192 28902 8193 28966
rect 8127 28901 8193 28902
rect 7359 3066 7425 3067
rect 7359 3002 7360 3066
rect 7424 3002 7425 3066
rect 7359 3001 7425 3002
rect 8130 2919 8190 28901
rect 19616 28670 19936 29938
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 27338 19936 28606
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 8319 26154 8385 26155
rect 8319 26090 8320 26154
rect 8384 26090 8385 26154
rect 8319 26089 8385 26090
rect 8322 3215 8382 26089
rect 19616 26006 19936 27274
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 24674 19936 25942
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 23342 19936 24610
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 22010 19936 23278
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 20678 19936 21946
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 19346 19936 20614
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 18014 19936 19282
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 16682 19936 17950
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 15350 19936 16618
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 14018 19936 15286
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 12686 19936 13954
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 11354 19936 12622
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 10022 19936 11290
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 10047 9134 10113 9135
rect 10047 9070 10048 9134
rect 10112 9070 10113 9134
rect 10047 9069 10113 9070
rect 9855 7506 9921 7507
rect 9855 7442 9856 7506
rect 9920 7442 9921 7506
rect 9855 7441 9921 7442
rect 9858 3955 9918 7441
rect 9855 3954 9921 3955
rect 9855 3890 9856 3954
rect 9920 3890 9921 3954
rect 9855 3889 9921 3890
rect 10050 3659 10110 9069
rect 19616 8690 19936 9958
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 7358 19936 8626
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 6026 19936 7294
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 4694 19936 5962
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 10047 3658 10113 3659
rect 10047 3594 10048 3658
rect 10112 3594 10113 3658
rect 10047 3593 10113 3594
rect 19616 3362 19936 4630
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 8319 3214 8385 3215
rect 8319 3150 8320 3214
rect 8384 3150 8385 3214
rect 8319 3149 8385 3150
rect 8127 2918 8193 2919
rect 8127 2854 8128 2918
rect 8192 2854 8193 2918
rect 8127 2853 8193 2854
rect 4256 2616 4576 2632
rect 19616 2616 19936 3298
rect 20276 2664 20596 57276
rect 20936 2664 21256 57276
rect 21596 2664 21916 57276
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 55976 35296 57244
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 54644 35296 55912
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 53312 35296 54580
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 51980 35296 53248
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 50648 35296 51916
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 49316 35296 50584
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 47984 35296 49252
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 46652 35296 47920
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 45320 35296 46588
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 43988 35296 45256
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 42656 35296 43924
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 41324 35296 42592
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 39992 35296 41260
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 38660 35296 39928
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 37328 35296 38596
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 35996 35296 37264
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 34664 35296 35932
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 33332 35296 34600
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 32000 35296 33268
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 30668 35296 31936
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 29336 35296 30604
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 28004 35296 29272
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 26672 35296 27940
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 25340 35296 26608
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 24008 35296 25276
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 22676 35296 23944
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 21344 35296 22612
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 20012 35296 21280
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 18680 35296 19948
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 17348 35296 18616
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 16016 35296 17284
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 14684 35296 15952
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 13352 35296 14620
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 12020 35296 13288
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 10688 35296 11956
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 9356 35296 10624
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 8024 35296 9292
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 28290 6963 29118 7023
rect 28290 6619 28350 6963
rect 29058 6767 29118 6963
rect 29055 6766 29121 6767
rect 29055 6702 29056 6766
rect 29120 6702 29121 6766
rect 29055 6701 29121 6702
rect 34976 6692 35296 7960
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 28287 6618 28353 6619
rect 28287 6554 28288 6618
rect 28352 6554 28353 6618
rect 28287 6553 28353 6554
rect 34976 5360 35296 6628
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 4028 35296 5296
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 2696 35296 3964
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 35636 2664 35956 57276
rect 36296 2664 36616 57276
rect 36956 2664 37276 57276
rect 50336 56642 50656 57324
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 55310 50656 56578
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 53978 50656 55246
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 52646 50656 53914
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 51314 50656 52582
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 49982 50656 51250
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 48650 50656 49918
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 47318 50656 48586
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 45986 50656 47254
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 44654 50656 45922
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 43322 50656 44590
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 41990 50656 43258
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 40658 50656 41926
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 39326 50656 40594
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 37994 50656 39262
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 36662 50656 37930
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 35330 50656 36598
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 33998 50656 35266
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 32666 50656 33934
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 31334 50656 32602
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 30002 50656 31270
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 28670 50656 29938
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 27338 50656 28606
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 26006 50656 27274
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 24674 50656 25942
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 23342 50656 24610
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 22010 50656 23278
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 20678 50656 21946
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 19346 50656 20614
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 18014 50656 19282
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 16682 50656 17950
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 15350 50656 16618
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 14018 50656 15286
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 12686 50656 13954
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 11354 50656 12622
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 10022 50656 11290
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 8690 50656 9958
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 7358 50656 8626
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 6026 50656 7294
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 4694 50656 5962
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 3362 50656 4630
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 34976 2616 35296 2632
rect 50336 2616 50656 3298
rect 50996 2664 51316 57276
rect 51656 2664 51976 57276
rect 52316 2664 52636 57276
use sky130_fd_sc_ls__clkbuf_1  input296 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input295
timestamp 1621261055
transform 1 0 1536 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_0
timestamp 1621261055
transform 1 0 1152 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_8
timestamp 1621261055
transform 1 0 1920 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_8
timestamp 1621261055
transform 1 0 1920 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input319
timestamp 1621261055
transform 1 0 2304 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input297
timestamp 1621261055
transform 1 0 2304 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_16
timestamp 1621261055
transform 1 0 2688 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_16
timestamp 1621261055
transform 1 0 2688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input323
timestamp 1621261055
transform 1 0 3072 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input322
timestamp 1621261055
transform 1 0 3072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_24
timestamp 1621261055
transform 1 0 3456 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3936 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_24
timestamp 1621261055
transform 1 0 3456 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input324
timestamp 1621261055
transform 1 0 3840 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_164 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3840 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_32
timestamp 1621261055
transform 1 0 4224 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 4704 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input325
timestamp 1621261055
transform 1 0 4608 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_40
timestamp 1621261055
transform 1 0 4992 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input298
timestamp 1621261055
transform 1 0 4896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_44
timestamp 1621261055
transform 1 0 5376 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_43
timestamp 1621261055
transform 1 0 5280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input300
timestamp 1621261055
transform 1 0 5568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_50
timestamp 1621261055
transform 1 0 5952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_51
timestamp 1621261055
transform 1 0 6048 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input299
timestamp 1621261055
transform 1 0 5664 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_56
timestamp 1621261055
transform 1 0 6528 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_54 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 6336 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_0_55
timestamp 1621261055
transform 1 0 6432 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_185
timestamp 1621261055
transform 1 0 6432 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_165
timestamp 1621261055
transform 1 0 6528 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_57
timestamp 1621261055
transform 1 0 6624 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input302
timestamp 1621261055
transform 1 0 6912 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input301
timestamp 1621261055
transform 1 0 7008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_64
timestamp 1621261055
transform 1 0 7296 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_65
timestamp 1621261055
transform 1 0 7392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input304
timestamp 1621261055
transform 1 0 7680 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input303
timestamp 1621261055
transform 1 0 7776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_80
timestamp 1621261055
transform 1 0 8832 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_72
timestamp 1621261055
transform 1 0 8064 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_73
timestamp 1621261055
transform 1 0 8160 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input306
timestamp 1621261055
transform 1 0 8448 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_83
timestamp 1621261055
transform 1 0 9120 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_81
timestamp 1621261055
transform 1 0 8928 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input309
timestamp 1621261055
transform 1 0 9216 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_166
timestamp 1621261055
transform 1 0 9216 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_88
timestamp 1621261055
transform 1 0 9600 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_85
timestamp 1621261055
transform 1 0 9312 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input311
timestamp 1621261055
transform 1 0 9984 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input307
timestamp 1621261055
transform 1 0 9696 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_96
timestamp 1621261055
transform 1 0 10368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_101
timestamp 1621261055
transform 1 0 10848 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_93
timestamp 1621261055
transform 1 0 10080 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input313
timestamp 1621261055
transform 1 0 10752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input310
timestamp 1621261055
transform 1 0 10464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_104
timestamp 1621261055
transform 1 0 11136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_111
timestamp 1621261055
transform 1 0 11808 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_108
timestamp 1621261055
transform 1 0 11520 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_113
timestamp 1621261055
transform 1 0 12000 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_0_111
timestamp 1621261055
transform 1 0 11808 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_109
timestamp 1621261055
transform 1 0 11616 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_186
timestamp 1621261055
transform 1 0 11712 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_167
timestamp 1621261055
transform 1 0 11904 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_118
timestamp 1621261055
transform 1 0 12480 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_121
timestamp 1621261055
transform 1 0 12768 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input167
timestamp 1621261055
transform 1 0 12864 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _114_ $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 12192 0 1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_126
timestamp 1621261055
transform 1 0 13248 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input39
timestamp 1621261055
transform 1 0 12960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_127
timestamp 1621261055
transform 1 0 13344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input89
timestamp 1621261055
transform 1 0 13632 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_134
timestamp 1621261055
transform 1 0 14016 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_135
timestamp 1621261055
transform 1 0 14112 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input78
timestamp 1621261055
transform 1 0 13728 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_139
timestamp 1621261055
transform 1 0 14496 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input100
timestamp 1621261055
transform 1 0 14400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_168
timestamp 1621261055
transform 1 0 14592 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_142
timestamp 1621261055
transform 1 0 14784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_141
timestamp 1621261055
transform 1 0 14688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input111 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 15072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input122
timestamp 1621261055
transform 1 0 15168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_150
timestamp 1621261055
transform 1 0 15552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_149
timestamp 1621261055
transform 1 0 15456 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input133
timestamp 1621261055
transform 1 0 15936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_164
timestamp 1621261055
transform 1 0 16896 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_162
timestamp 1621261055
transform 1 0 16704 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_158
timestamp 1621261055
transform 1 0 16320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_164
timestamp 1621261055
transform 1 0 16896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_159
timestamp 1621261055
transform 1 0 16416 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_157
timestamp 1621261055
transform 1 0 16224 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input50
timestamp 1621261055
transform 1 0 16512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_166
timestamp 1621261055
transform 1 0 17088 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_187
timestamp 1621261055
transform 1 0 16992 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_169
timestamp 1621261055
transform 1 0 17280 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_169
timestamp 1621261055
transform 1 0 17376 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input70
timestamp 1621261055
transform 1 0 17472 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_174
timestamp 1621261055
transform 1 0 17856 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_177
timestamp 1621261055
transform 1 0 18144 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input61
timestamp 1621261055
transform 1 0 17760 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_182
timestamp 1621261055
transform 1 0 18624 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input72
timestamp 1621261055
transform 1 0 18240 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input71
timestamp 1621261055
transform 1 0 18528 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_185
timestamp 1621261055
transform 1 0 18912 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_33 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 19104 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input73
timestamp 1621261055
transform 1 0 19008 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _020_
timestamp 1621261055
transform 1 0 19296 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_190
timestamp 1621261055
transform 1 0 19392 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_192
timestamp 1621261055
transform 1 0 19584 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_198
timestamp 1621261055
transform 1 0 20160 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_197
timestamp 1621261055
transform 1 0 20064 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input75
timestamp 1621261055
transform 1 0 19776 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_170
timestamp 1621261055
transform 1 0 19968 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__buf_1  input77
timestamp 1621261055
transform 1 0 20544 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input74
timestamp 1621261055
transform 1 0 20448 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_206
timestamp 1621261055
transform 1 0 20928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_205
timestamp 1621261055
transform 1 0 20832 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input80
timestamp 1621261055
transform 1 0 21312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input76
timestamp 1621261055
transform 1 0 21216 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_214
timestamp 1621261055
transform 1 0 21696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_213
timestamp 1621261055
transform 1 0 21600 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_218
timestamp 1621261055
transform 1 0 22080 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _082_
timestamp 1621261055
transform 1 0 21984 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_221
timestamp 1621261055
transform 1 0 22368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_220
timestamp 1621261055
transform 1 0 22272 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_188
timestamp 1621261055
transform 1 0 22272 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_171
timestamp 1621261055
transform 1 0 22656 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_229
timestamp 1621261055
transform 1 0 23136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_225
timestamp 1621261055
transform 1 0 22752 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input84
timestamp 1621261055
transform 1 0 22752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input82
timestamp 1621261055
transform 1 0 23136 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_237
timestamp 1621261055
transform 1 0 23904 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_233
timestamp 1621261055
transform 1 0 23520 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input86
timestamp 1621261055
transform 1 0 23520 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input85
timestamp 1621261055
transform 1 0 23904 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_245
timestamp 1621261055
transform 1 0 24672 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_241
timestamp 1621261055
transform 1 0 24288 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input88
timestamp 1621261055
transform 1 0 24288 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_251
timestamp 1621261055
transform 1 0 25248 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_249
timestamp 1621261055
transform 1 0 25056 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input91
timestamp 1621261055
transform 1 0 25056 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_172
timestamp 1621261055
transform 1 0 25344 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_253
timestamp 1621261055
transform 1 0 25440 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_253
timestamp 1621261055
transform 1 0 25440 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input92
timestamp 1621261055
transform 1 0 25824 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input90
timestamp 1621261055
transform 1 0 25824 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_269
timestamp 1621261055
transform 1 0 26976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_261
timestamp 1621261055
transform 1 0 26208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_269
timestamp 1621261055
transform 1 0 26976 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_261
timestamp 1621261055
transform 1 0 26208 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input95
timestamp 1621261055
transform 1 0 26592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input93
timestamp 1621261055
transform 1 0 26592 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_273
timestamp 1621261055
transform 1 0 27360 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_276
timestamp 1621261055
transform 1 0 27648 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_277
timestamp 1621261055
transform 1 0 27744 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_189
timestamp 1621261055
transform 1 0 27552 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_281
timestamp 1621261055
transform 1 0 28128 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_279
timestamp 1621261055
transform 1 0 27936 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input99
timestamp 1621261055
transform 1 0 28032 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_173
timestamp 1621261055
transform 1 0 28032 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_284
timestamp 1621261055
transform 1 0 28416 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input98
timestamp 1621261055
transform 1 0 28512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_292
timestamp 1621261055
transform 1 0 29184 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_289
timestamp 1621261055
transform 1 0 28896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input102
timestamp 1621261055
transform 1 0 28800 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input101
timestamp 1621261055
transform 1 0 29280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_300
timestamp 1621261055
transform 1 0 29952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_297
timestamp 1621261055
transform 1 0 29664 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input104
timestamp 1621261055
transform 1 0 29568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_308
timestamp 1621261055
transform 1 0 30720 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_309
timestamp 1621261055
transform 1 0 30816 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_307
timestamp 1621261055
transform 1 0 30624 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_305
timestamp 1621261055
transform 1 0 30432 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input106
timestamp 1621261055
transform 1 0 30336 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_174
timestamp 1621261055
transform 1 0 30720 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input108
timestamp 1621261055
transform 1 0 31104 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input107
timestamp 1621261055
transform 1 0 31200 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_316
timestamp 1621261055
transform 1 0 31488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_317
timestamp 1621261055
transform 1 0 31584 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input112
timestamp 1621261055
transform 1 0 31872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input109
timestamp 1621261055
transform 1 0 31968 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_331
timestamp 1621261055
transform 1 0 32928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_328
timestamp 1621261055
transform 1 0 32640 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_324
timestamp 1621261055
transform 1 0 32256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_325
timestamp 1621261055
transform 1 0 32352 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_190
timestamp 1621261055
transform 1 0 32832 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_0_335
timestamp 1621261055
transform 1 0 33312 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_333
timestamp 1621261055
transform 1 0 33120 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input115
timestamp 1621261055
transform 1 0 33312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_175
timestamp 1621261055
transform 1 0 33408 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_339
timestamp 1621261055
transform 1 0 33696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_337
timestamp 1621261055
transform 1 0 33504 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_345
timestamp 1621261055
transform 1 0 34272 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input118
timestamp 1621261055
transform 1 0 34080 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input114
timestamp 1621261055
transform 1 0 33888 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_347
timestamp 1621261055
transform 1 0 34464 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input117
timestamp 1621261055
transform 1 0 34656 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_355
timestamp 1621261055
transform 1 0 35232 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_353
timestamp 1621261055
transform 1 0 35040 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_12
timestamp 1621261055
transform -1 0 35424 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input120
timestamp 1621261055
transform 1 0 34848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _006_
timestamp 1621261055
transform -1 0 35712 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_360
timestamp 1621261055
transform 1 0 35712 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input123
timestamp 1621261055
transform 1 0 35616 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_363
timestamp 1621261055
transform 1 0 36000 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_365
timestamp 1621261055
transform 1 0 36192 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_176
timestamp 1621261055
transform 1 0 36096 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_371
timestamp 1621261055
transform 1 0 36768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input125
timestamp 1621261055
transform 1 0 36384 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input124
timestamp 1621261055
transform 1 0 36576 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_373
timestamp 1621261055
transform 1 0 36960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input127
timestamp 1621261055
transform 1 0 37152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input126
timestamp 1621261055
transform 1 0 37344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_386
timestamp 1621261055
transform 1 0 38208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_383
timestamp 1621261055
transform 1 0 37920 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_379
timestamp 1621261055
transform 1 0 37536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_381
timestamp 1621261055
transform 1 0 37728 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_191
timestamp 1621261055
transform 1 0 38112 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_394
timestamp 1621261055
transform 1 0 38976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_393
timestamp 1621261055
transform 1 0 38880 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_391
timestamp 1621261055
transform 1 0 38688 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_389
timestamp 1621261055
transform 1 0 38496 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input131
timestamp 1621261055
transform 1 0 38592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_177
timestamp 1621261055
transform 1 0 38784 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input134
timestamp 1621261055
transform 1 0 39360 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input130
timestamp 1621261055
transform 1 0 39264 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_402
timestamp 1621261055
transform 1 0 39744 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_401
timestamp 1621261055
transform 1 0 39648 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input136
timestamp 1621261055
transform 1 0 40128 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input132
timestamp 1621261055
transform 1 0 40032 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_410
timestamp 1621261055
transform 1 0 40512 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_409
timestamp 1621261055
transform 1 0 40416 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input138
timestamp 1621261055
transform 1 0 40896 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_418
timestamp 1621261055
transform 1 0 41280 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_419
timestamp 1621261055
transform 1 0 41376 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_417
timestamp 1621261055
transform 1 0 41184 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_178
timestamp 1621261055
transform 1 0 41472 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_421
timestamp 1621261055
transform 1 0 41568 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input140
timestamp 1621261055
transform 1 0 41664 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input139
timestamp 1621261055
transform 1 0 41952 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_426
timestamp 1621261055
transform 1 0 42048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_429
timestamp 1621261055
transform 1 0 42336 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_434
timestamp 1621261055
transform 1 0 42816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input142
timestamp 1621261055
transform 1 0 42432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input141
timestamp 1621261055
transform 1 0 42720 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_438
timestamp 1621261055
transform 1 0 43200 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_437
timestamp 1621261055
transform 1 0 43104 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_441
timestamp 1621261055
transform 1 0 43488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_192
timestamp 1621261055
transform 1 0 43392 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _139_
timestamp 1621261055
transform 1 0 43488 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_444
timestamp 1621261055
transform 1 0 43776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input146
timestamp 1621261055
transform 1 0 43872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_449
timestamp 1621261055
transform 1 0 44256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_449
timestamp 1621261055
transform 1 0 44256 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_179
timestamp 1621261055
transform 1 0 44160 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input149
timestamp 1621261055
transform 1 0 44640 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input147
timestamp 1621261055
transform 1 0 44640 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_457
timestamp 1621261055
transform 1 0 45024 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_457
timestamp 1621261055
transform 1 0 45024 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input151
timestamp 1621261055
transform 1 0 45408 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input150
timestamp 1621261055
transform 1 0 45408 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_465
timestamp 1621261055
transform 1 0 45792 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_465
timestamp 1621261055
transform 1 0 45792 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input153
timestamp 1621261055
transform 1 0 46176 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _195_
timestamp 1621261055
transform 1 0 46176 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_473
timestamp 1621261055
transform 1 0 46560 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_472
timestamp 1621261055
transform 1 0 46464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_180
timestamp 1621261055
transform 1 0 46848 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_481
timestamp 1621261055
transform 1 0 47328 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_477
timestamp 1621261055
transform 1 0 46944 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input156
timestamp 1621261055
transform 1 0 46944 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input154
timestamp 1621261055
transform 1 0 47328 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_489
timestamp 1621261055
transform 1 0 48096 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_485
timestamp 1621261055
transform 1 0 47712 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input159
timestamp 1621261055
transform 1 0 47712 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input157
timestamp 1621261055
transform 1 0 48096 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_496
timestamp 1621261055
transform 1 0 48768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_493
timestamp 1621261055
transform 1 0 48480 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_493
timestamp 1621261055
transform 1 0 48480 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input162
timestamp 1621261055
transform 1 0 49152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_193
timestamp 1621261055
transform 1 0 48672 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_504
timestamp 1621261055
transform 1 0 49536 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_0_503
timestamp 1621261055
transform 1 0 49440 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_501
timestamp 1621261055
transform 1 0 49248 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_181
timestamp 1621261055
transform 1 0 49536 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_505
timestamp 1621261055
transform 1 0 49632 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input40
timestamp 1621261055
transform 1 0 50016 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_512
timestamp 1621261055
transform 1 0 50304 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_513
timestamp 1621261055
transform 1 0 50400 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input42
timestamp 1621261055
transform 1 0 50400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_517
timestamp 1621261055
transform 1 0 50784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input41
timestamp 1621261055
transform 1 0 50784 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_521
timestamp 1621261055
transform 1 0 51168 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input43
timestamp 1621261055
transform 1 0 51168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_525
timestamp 1621261055
transform 1 0 51552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _130_
timestamp 1621261055
transform 1 0 51552 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_533
timestamp 1621261055
transform 1 0 52320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_533
timestamp 1621261055
transform 1 0 52320 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_528
timestamp 1621261055
transform 1 0 51840 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input44
timestamp 1621261055
transform 1 0 51936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_182
timestamp 1621261055
transform 1 0 52224 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_541
timestamp 1621261055
transform 1 0 53088 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_541
timestamp 1621261055
transform 1 0 53088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input46
timestamp 1621261055
transform 1 0 52704 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input45
timestamp 1621261055
transform 1 0 52704 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input47
timestamp 1621261055
transform 1 0 53472 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_551
timestamp 1621261055
transform 1 0 54048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_549
timestamp 1621261055
transform 1 0 53856 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_549
timestamp 1621261055
transform 1 0 53856 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_194
timestamp 1621261055
transform 1 0 53952 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input51
timestamp 1621261055
transform 1 0 54432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _120_
timestamp 1621261055
transform 1 0 54240 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_559
timestamp 1621261055
transform 1 0 54816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_556
timestamp 1621261055
transform 1 0 54528 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_183
timestamp 1621261055
transform 1 0 54912 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_561
timestamp 1621261055
transform 1 0 55008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input54
timestamp 1621261055
transform 1 0 55200 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input52
timestamp 1621261055
transform 1 0 55392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_567
timestamp 1621261055
transform 1 0 55584 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_569
timestamp 1621261055
transform 1 0 55776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input56
timestamp 1621261055
transform 1 0 55968 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_575
timestamp 1621261055
transform 1 0 56352 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input55
timestamp 1621261055
transform 1 0 56160 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_577
timestamp 1621261055
transform 1 0 56544 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_31
timestamp 1621261055
transform 1 0 56736 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input58
timestamp 1621261055
transform 1 0 56736 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _019_
timestamp 1621261055
transform 1 0 56928 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_583
timestamp 1621261055
transform 1 0 57120 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_584
timestamp 1621261055
transform 1 0 57216 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input59
timestamp 1621261055
transform 1 0 57504 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_184
timestamp 1621261055
transform 1 0 57600 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_1
timestamp 1621261055
transform -1 0 58848 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_3
timestamp 1621261055
transform -1 0 58848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_589
timestamp 1621261055
transform 1 0 57696 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_1_591
timestamp 1621261055
transform 1 0 57888 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_595
timestamp 1621261055
transform 1 0 58272 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_4
timestamp 1621261055
transform 1 0 1152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input308
timestamp 1621261055
transform 1 0 1536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input330
timestamp 1621261055
transform 1 0 2304 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input341
timestamp 1621261055
transform 1 0 3072 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_8
timestamp 1621261055
transform 1 0 1920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_16
timestamp 1621261055
transform 1 0 2688 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_195
timestamp 1621261055
transform 1 0 3840 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input326
timestamp 1621261055
transform 1 0 4320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input328
timestamp 1621261055
transform 1 0 5088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_24
timestamp 1621261055
transform 1 0 3456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_29
timestamp 1621261055
transform 1 0 3936 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_37
timestamp 1621261055
transform 1 0 4704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input331
timestamp 1621261055
transform 1 0 5856 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input333
timestamp 1621261055
transform 1 0 6624 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_45
timestamp 1621261055
transform 1 0 5472 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_53
timestamp 1621261055
transform 1 0 6240 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_61
timestamp 1621261055
transform 1 0 7008 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_196
timestamp 1621261055
transform 1 0 9120 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input305
timestamp 1621261055
transform 1 0 7392 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input335
timestamp 1621261055
transform 1 0 8160 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_69
timestamp 1621261055
transform 1 0 7776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_77
timestamp 1621261055
transform 1 0 8544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_81
timestamp 1621261055
transform 1 0 8928 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_84
timestamp 1621261055
transform 1 0 9216 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input312
timestamp 1621261055
transform 1 0 9600 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input314
timestamp 1621261055
transform 1 0 10368 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input315
timestamp 1621261055
transform 1 0 11136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_92
timestamp 1621261055
transform 1 0 9984 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_100
timestamp 1621261055
transform 1 0 10752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input316
timestamp 1621261055
transform 1 0 11904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input317
timestamp 1621261055
transform 1 0 12672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_108
timestamp 1621261055
transform 1 0 11520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_116
timestamp 1621261055
transform 1 0 12288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_124
timestamp 1621261055
transform 1 0 13056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_197
timestamp 1621261055
transform 1 0 14400 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input206
timestamp 1621261055
transform 1 0 13536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_128
timestamp 1621261055
transform 1 0 13440 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_133
timestamp 1621261055
transform 1 0 13920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_137
timestamp 1621261055
transform 1 0 14304 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_139
timestamp 1621261055
transform 1 0 14496 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_147
timestamp 1621261055
transform 1 0 15264 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input144
timestamp 1621261055
transform 1 0 15456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input155
timestamp 1621261055
transform 1 0 16224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input166
timestamp 1621261055
transform 1 0 16992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_153
timestamp 1621261055
transform 1 0 15840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_161
timestamp 1621261055
transform 1 0 16608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input178
timestamp 1621261055
transform 1 0 17760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input198
timestamp 1621261055
transform 1 0 18528 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_169
timestamp 1621261055
transform 1 0 17376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_177
timestamp 1621261055
transform 1 0 18144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_185
timestamp 1621261055
transform 1 0 18912 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_198
timestamp 1621261055
transform 1 0 19680 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input79
timestamp 1621261055
transform 1 0 20256 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input81
timestamp 1621261055
transform 1 0 21024 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_194
timestamp 1621261055
transform 1 0 19776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_198
timestamp 1621261055
transform 1 0 20160 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_203
timestamp 1621261055
transform 1 0 20640 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _074_
timestamp 1621261055
transform 1 0 22560 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input83
timestamp 1621261055
transform 1 0 21792 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input87
timestamp 1621261055
transform 1 0 23232 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_211
timestamp 1621261055
transform 1 0 21408 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_219
timestamp 1621261055
transform 1 0 22176 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_226
timestamp 1621261055
transform 1 0 22848 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_199
timestamp 1621261055
transform 1 0 24960 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input211
timestamp 1621261055
transform 1 0 24000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_234
timestamp 1621261055
transform 1 0 23616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_242
timestamp 1621261055
transform 1 0 24384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_246
timestamp 1621261055
transform 1 0 24768 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_249
timestamp 1621261055
transform 1 0 25056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input94
timestamp 1621261055
transform 1 0 25440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input96
timestamp 1621261055
transform 1 0 26208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input97
timestamp 1621261055
transform 1 0 26976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_257
timestamp 1621261055
transform 1 0 25824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_265
timestamp 1621261055
transform 1 0 26592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_273
timestamp 1621261055
transform 1 0 27360 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input103
timestamp 1621261055
transform 1 0 28320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input105
timestamp 1621261055
transform 1 0 29088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_281
timestamp 1621261055
transform 1 0 28128 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_287
timestamp 1621261055
transform 1 0 28704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_200
timestamp 1621261055
transform 1 0 30240 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input110
timestamp 1621261055
transform 1 0 30912 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_295
timestamp 1621261055
transform 1 0 29472 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_304
timestamp 1621261055
transform 1 0 30336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_308
timestamp 1621261055
transform 1 0 30720 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_314
timestamp 1621261055
transform 1 0 31296 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input113
timestamp 1621261055
transform 1 0 31680 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input116
timestamp 1621261055
transform 1 0 32736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_322
timestamp 1621261055
transform 1 0 32064 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_326
timestamp 1621261055
transform 1 0 32448 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_328
timestamp 1621261055
transform 1 0 32640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_333
timestamp 1621261055
transform 1 0 33120 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input119
timestamp 1621261055
transform 1 0 33888 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input121
timestamp 1621261055
transform 1 0 34656 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_345
timestamp 1621261055
transform 1 0 34272 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_353
timestamp 1621261055
transform 1 0 35040 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_357
timestamp 1621261055
transform 1 0 35424 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_201
timestamp 1621261055
transform 1 0 35520 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input128
timestamp 1621261055
transform 1 0 36768 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input247
timestamp 1621261055
transform 1 0 36000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_359
timestamp 1621261055
transform 1 0 35616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_367
timestamp 1621261055
transform 1 0 36384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_375
timestamp 1621261055
transform 1 0 37152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input129
timestamp 1621261055
transform 1 0 37536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input135
timestamp 1621261055
transform 1 0 38976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_383
timestamp 1621261055
transform 1 0 37920 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_391
timestamp 1621261055
transform 1 0 38688 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_393
timestamp 1621261055
transform 1 0 38880 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_398
timestamp 1621261055
transform 1 0 39360 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_202
timestamp 1621261055
transform 1 0 40800 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input137
timestamp 1621261055
transform 1 0 39744 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_406
timestamp 1621261055
transform 1 0 40128 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_410
timestamp 1621261055
transform 1 0 40512 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_412
timestamp 1621261055
transform 1 0 40704 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_414
timestamp 1621261055
transform 1 0 40896 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input143
timestamp 1621261055
transform 1 0 41952 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input145
timestamp 1621261055
transform 1 0 42720 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input148
timestamp 1621261055
transform 1 0 43488 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_422
timestamp 1621261055
transform 1 0 41664 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_424
timestamp 1621261055
transform 1 0 41856 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_429
timestamp 1621261055
transform 1 0 42336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_437
timestamp 1621261055
transform 1 0 43104 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _048_
timestamp 1621261055
transform -1 0 44544 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input152
timestamp 1621261055
transform 1 0 44928 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_53
timestamp 1621261055
transform -1 0 44256 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_445
timestamp 1621261055
transform 1 0 43872 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_452
timestamp 1621261055
transform 1 0 44544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_460
timestamp 1621261055
transform 1 0 45312 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_203
timestamp 1621261055
transform 1 0 46080 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input158
timestamp 1621261055
transform 1 0 46752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input160
timestamp 1621261055
transform 1 0 47520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_469
timestamp 1621261055
transform 1 0 46176 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_473
timestamp 1621261055
transform 1 0 46560 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_479
timestamp 1621261055
transform 1 0 47136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input161
timestamp 1621261055
transform 1 0 48288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input163
timestamp 1621261055
transform 1 0 49056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_487
timestamp 1621261055
transform 1 0 47904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_495
timestamp 1621261055
transform 1 0 48672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_503
timestamp 1621261055
transform 1 0 49440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_204
timestamp 1621261055
transform 1 0 51360 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input164
timestamp 1621261055
transform 1 0 49824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input168
timestamp 1621261055
transform 1 0 50592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_511
timestamp 1621261055
transform 1 0 50208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_519
timestamp 1621261055
transform 1 0 50976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_524
timestamp 1621261055
transform 1 0 51456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input48
timestamp 1621261055
transform 1 0 52608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input49
timestamp 1621261055
transform 1 0 53376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input171
timestamp 1621261055
transform 1 0 51840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_532
timestamp 1621261055
transform 1 0 52224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_540
timestamp 1621261055
transform 1 0 52992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _079_
timestamp 1621261055
transform 1 0 54912 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input53
timestamp 1621261055
transform 1 0 54144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input57
timestamp 1621261055
transform 1 0 55584 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_548
timestamp 1621261055
transform 1 0 53760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_556
timestamp 1621261055
transform 1 0 54528 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_563
timestamp 1621261055
transform 1 0 55200 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_205
timestamp 1621261055
transform 1 0 56640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input60
timestamp 1621261055
transform 1 0 57120 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_571
timestamp 1621261055
transform 1 0 55968 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_575
timestamp 1621261055
transform 1 0 56352 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_577
timestamp 1621261055
transform 1 0 56544 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_579
timestamp 1621261055
transform 1 0 56736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_587
timestamp 1621261055
transform 1 0 57504 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_5
timestamp 1621261055
transform -1 0 58848 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_595
timestamp 1621261055
transform 1 0 58272 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_6
timestamp 1621261055
transform 1 0 1152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input329
timestamp 1621261055
transform 1 0 1536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input352
timestamp 1621261055
transform 1 0 2304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input355
timestamp 1621261055
transform 1 0 3072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_8
timestamp 1621261055
transform 1 0 1920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_16
timestamp 1621261055
transform 1 0 2688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input327
timestamp 1621261055
transform 1 0 4128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_24
timestamp 1621261055
transform 1 0 3456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_28
timestamp 1621261055
transform 1 0 3840 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_30
timestamp 1621261055
transform 1 0 4032 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_3_35
timestamp 1621261055
transform 1 0 4512 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_206
timestamp 1621261055
transform 1 0 6432 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input332
timestamp 1621261055
transform 1 0 5376 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input334
timestamp 1621261055
transform 1 0 6912 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_43
timestamp 1621261055
transform 1 0 5280 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_3_48
timestamp 1621261055
transform 1 0 5760 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_52
timestamp 1621261055
transform 1 0 6144 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_54
timestamp 1621261055
transform 1 0 6336 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_3_56
timestamp 1621261055
transform 1 0 6528 0 1 4662
box -38 -49 422 715
use AND2X1  AND2X1
timestamp 1624074425
transform 1 0 7680 0 1 4662
box 0 -48 1152 714
use sky130_fd_sc_ls__clkbuf_1  input339
timestamp 1621261055
transform 1 0 9216 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_71
timestamp 1621261055
transform 1 0 7488 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_64
timestamp 1621261055
transform 1 0 7296 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_80
timestamp 1621261055
transform 1 0 8832 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input340
timestamp 1621261055
transform 1 0 9984 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input343
timestamp 1621261055
transform 1 0 10752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_88
timestamp 1621261055
transform 1 0 9600 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_96
timestamp 1621261055
transform 1 0 10368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_104
timestamp 1621261055
transform 1 0 11136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_207
timestamp 1621261055
transform 1 0 11712 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input318
timestamp 1621261055
transform 1 0 12192 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input320
timestamp 1621261055
transform 1 0 12960 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_108
timestamp 1621261055
transform 1 0 11520 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_111
timestamp 1621261055
transform 1 0 11808 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_119
timestamp 1621261055
transform 1 0 12576 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input217
timestamp 1621261055
transform 1 0 13920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input228
timestamp 1621261055
transform 1 0 14688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_127
timestamp 1621261055
transform 1 0 13344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_131
timestamp 1621261055
transform 1 0 13728 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_137
timestamp 1621261055
transform 1 0 14304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_145
timestamp 1621261055
transform 1 0 15072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_208
timestamp 1621261055
transform 1 0 16992 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input239
timestamp 1621261055
transform 1 0 15456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input261
timestamp 1621261055
transform 1 0 16224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_153
timestamp 1621261055
transform 1 0 15840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_161
timestamp 1621261055
transform 1 0 16608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_166
timestamp 1621261055
transform 1 0 17088 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input189
timestamp 1621261055
transform 1 0 17472 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input199
timestamp 1621261055
transform 1 0 18240 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input200
timestamp 1621261055
transform 1 0 19008 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_174
timestamp 1621261055
transform 1 0 17856 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_182
timestamp 1621261055
transform 1 0 18624 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input202
timestamp 1621261055
transform 1 0 19776 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input203
timestamp 1621261055
transform 1 0 20544 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input205
timestamp 1621261055
transform 1 0 21312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_190
timestamp 1621261055
transform 1 0 19392 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_198
timestamp 1621261055
transform 1 0 20160 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_206
timestamp 1621261055
transform 1 0 20928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_209
timestamp 1621261055
transform 1 0 22272 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input209
timestamp 1621261055
transform 1 0 22752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_214
timestamp 1621261055
transform 1 0 21696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_218
timestamp 1621261055
transform 1 0 22080 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_221
timestamp 1621261055
transform 1 0 22368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_229
timestamp 1621261055
transform 1 0 23136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input212
timestamp 1621261055
transform 1 0 23520 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input214
timestamp 1621261055
transform 1 0 24288 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input216
timestamp 1621261055
transform 1 0 25056 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_237
timestamp 1621261055
transform 1 0 23904 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_245
timestamp 1621261055
transform 1 0 24672 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input218
timestamp 1621261055
transform 1 0 25824 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input220
timestamp 1621261055
transform 1 0 26592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_253
timestamp 1621261055
transform 1 0 25440 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_261
timestamp 1621261055
transform 1 0 26208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_269
timestamp 1621261055
transform 1 0 26976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_273
timestamp 1621261055
transform 1 0 27360 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_210
timestamp 1621261055
transform 1 0 27552 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input224
timestamp 1621261055
transform 1 0 28032 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input227
timestamp 1621261055
transform 1 0 28800 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_276
timestamp 1621261055
transform 1 0 27648 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_284
timestamp 1621261055
transform 1 0 28416 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_292
timestamp 1621261055
transform 1 0 29184 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input230
timestamp 1621261055
transform 1 0 29568 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input232
timestamp 1621261055
transform 1 0 30336 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input233
timestamp 1621261055
transform 1 0 31104 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_300
timestamp 1621261055
transform 1 0 29952 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_308
timestamp 1621261055
transform 1 0 30720 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_211
timestamp 1621261055
transform 1 0 32832 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input236
timestamp 1621261055
transform 1 0 31872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input241
timestamp 1621261055
transform 1 0 33312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_316
timestamp 1621261055
transform 1 0 31488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_324
timestamp 1621261055
transform 1 0 32256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_328
timestamp 1621261055
transform 1 0 32640 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_331
timestamp 1621261055
transform 1 0 32928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input243
timestamp 1621261055
transform 1 0 34080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input245
timestamp 1621261055
transform 1 0 34848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_339
timestamp 1621261055
transform 1 0 33696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_347
timestamp 1621261055
transform 1 0 34464 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_355
timestamp 1621261055
transform 1 0 35232 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input248
timestamp 1621261055
transform 1 0 35616 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input249
timestamp 1621261055
transform 1 0 36384 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input252
timestamp 1621261055
transform 1 0 37152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_363
timestamp 1621261055
transform 1 0 36000 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_371
timestamp 1621261055
transform 1 0 36768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_212
timestamp 1621261055
transform 1 0 38112 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input256
timestamp 1621261055
transform 1 0 38592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input258
timestamp 1621261055
transform 1 0 39360 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_379
timestamp 1621261055
transform 1 0 37536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_383
timestamp 1621261055
transform 1 0 37920 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_386
timestamp 1621261055
transform 1 0 38208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_394
timestamp 1621261055
transform 1 0 38976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input260
timestamp 1621261055
transform 1 0 40128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input264
timestamp 1621261055
transform 1 0 40896 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_402
timestamp 1621261055
transform 1 0 39744 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_410
timestamp 1621261055
transform 1 0 40512 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_418
timestamp 1621261055
transform 1 0 41280 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_213
timestamp 1621261055
transform 1 0 43392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input265
timestamp 1621261055
transform 1 0 41664 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input268
timestamp 1621261055
transform 1 0 42432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_426
timestamp 1621261055
transform 1 0 42048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_434
timestamp 1621261055
transform 1 0 42816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_438
timestamp 1621261055
transform 1 0 43200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_441
timestamp 1621261055
transform 1 0 43488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input273
timestamp 1621261055
transform 1 0 43872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input275
timestamp 1621261055
transform 1 0 44640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input277
timestamp 1621261055
transform 1 0 45408 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_449
timestamp 1621261055
transform 1 0 44256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_457
timestamp 1621261055
transform 1 0 45024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input279
timestamp 1621261055
transform 1 0 46176 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input280
timestamp 1621261055
transform 1 0 46944 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_465
timestamp 1621261055
transform 1 0 45792 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_473
timestamp 1621261055
transform 1 0 46560 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_481
timestamp 1621261055
transform 1 0 47328 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_214
timestamp 1621261055
transform 1 0 48672 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input165
timestamp 1621261055
transform 1 0 49344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input284
timestamp 1621261055
transform 1 0 47712 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_489
timestamp 1621261055
transform 1 0 48096 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_493
timestamp 1621261055
transform 1 0 48480 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_496
timestamp 1621261055
transform 1 0 48768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_500
timestamp 1621261055
transform 1 0 49152 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input169
timestamp 1621261055
transform 1 0 50304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input170
timestamp 1621261055
transform 1 0 51072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_506
timestamp 1621261055
transform 1 0 49728 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_510
timestamp 1621261055
transform 1 0 50112 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_516
timestamp 1621261055
transform 1 0 50688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_524
timestamp 1621261055
transform 1 0 51456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input172
timestamp 1621261055
transform 1 0 51840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input173
timestamp 1621261055
transform 1 0 52608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_532
timestamp 1621261055
transform 1 0 52224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_540
timestamp 1621261055
transform 1 0 52992 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_215
timestamp 1621261055
transform 1 0 53952 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input68
timestamp 1621261055
transform 1 0 55488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input177
timestamp 1621261055
transform 1 0 54432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_548
timestamp 1621261055
transform 1 0 53760 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_551
timestamp 1621261055
transform 1 0 54048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_559
timestamp 1621261055
transform 1 0 54816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_563
timestamp 1621261055
transform 1 0 55200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_565
timestamp 1621261055
transform 1 0 55392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input62
timestamp 1621261055
transform 1 0 57024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input64
timestamp 1621261055
transform 1 0 56256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_14
timestamp 1621261055
transform 1 0 57600 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_570
timestamp 1621261055
transform 1 0 55872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_578
timestamp 1621261055
transform 1 0 56640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_586
timestamp 1621261055
transform 1 0 57408 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _007_
timestamp 1621261055
transform 1 0 57792 0 1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_7
timestamp 1621261055
transform -1 0 58848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_593
timestamp 1621261055
transform 1 0 58080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_8
timestamp 1621261055
transform 1 0 1152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input356
timestamp 1621261055
transform 1 0 2784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input362
timestamp 1621261055
transform 1 0 1536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_8
timestamp 1621261055
transform 1 0 1920 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_4_16
timestamp 1621261055
transform 1 0 2688 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_21
timestamp 1621261055
transform 1 0 3168 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_216
timestamp 1621261055
transform 1 0 3840 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input358
timestamp 1621261055
transform 1 0 4320 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input360
timestamp 1621261055
transform 1 0 5088 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_25
timestamp 1621261055
transform 1 0 3552 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_27
timestamp 1621261055
transform 1 0 3744 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_29
timestamp 1621261055
transform 1 0 3936 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_37
timestamp 1621261055
transform 1 0 4704 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input336
timestamp 1621261055
transform 1 0 6816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output574 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 5856 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_211
timestamp 1621261055
transform 1 0 5664 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_45
timestamp 1621261055
transform 1 0 5472 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_53
timestamp 1621261055
transform 1 0 6240 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_57
timestamp 1621261055
transform 1 0 6624 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_63
timestamp 1621261055
transform 1 0 7200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_217
timestamp 1621261055
transform 1 0 9120 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input337
timestamp 1621261055
transform 1 0 7584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input338
timestamp 1621261055
transform 1 0 8352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_71
timestamp 1621261055
transform 1 0 7968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_79
timestamp 1621261055
transform 1 0 8736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_84
timestamp 1621261055
transform 1 0 9216 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input342
timestamp 1621261055
transform 1 0 9600 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input345
timestamp 1621261055
transform 1 0 10368 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input347
timestamp 1621261055
transform 1 0 11136 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_92
timestamp 1621261055
transform 1 0 9984 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_100
timestamp 1621261055
transform 1 0 10752 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _147_
timestamp 1621261055
transform 1 0 11904 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input321
timestamp 1621261055
transform 1 0 12576 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_108
timestamp 1621261055
transform 1 0 11520 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_115
timestamp 1621261055
transform 1 0 12192 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_123
timestamp 1621261055
transform 1 0 12960 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_218
timestamp 1621261055
transform 1 0 14400 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input250
timestamp 1621261055
transform 1 0 14976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input351
timestamp 1621261055
transform 1 0 13344 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_131
timestamp 1621261055
transform 1 0 13728 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_135
timestamp 1621261055
transform 1 0 14112 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_137
timestamp 1621261055
transform 1 0 14304 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_139
timestamp 1621261055
transform 1 0 14496 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_143
timestamp 1621261055
transform 1 0 14880 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input272
timestamp 1621261055
transform 1 0 15744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input283
timestamp 1621261055
transform 1 0 16512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input294
timestamp 1621261055
transform 1 0 17280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_148
timestamp 1621261055
transform 1 0 15360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_156
timestamp 1621261055
transform 1 0 16128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_164
timestamp 1621261055
transform 1 0 16896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input201
timestamp 1621261055
transform 1 0 18720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_172
timestamp 1621261055
transform 1 0 17664 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_180
timestamp 1621261055
transform 1 0 18432 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_182
timestamp 1621261055
transform 1 0 18624 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_187
timestamp 1621261055
transform 1 0 19104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_219
timestamp 1621261055
transform 1 0 19680 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input204
timestamp 1621261055
transform 1 0 20160 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input207
timestamp 1621261055
transform 1 0 20928 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_191
timestamp 1621261055
transform 1 0 19488 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_194
timestamp 1621261055
transform 1 0 19776 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_202
timestamp 1621261055
transform 1 0 20544 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_210
timestamp 1621261055
transform 1 0 21312 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input208
timestamp 1621261055
transform 1 0 21696 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input210
timestamp 1621261055
transform 1 0 22464 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input213
timestamp 1621261055
transform 1 0 23232 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_218
timestamp 1621261055
transform 1 0 22080 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_226
timestamp 1621261055
transform 1 0 22848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_220
timestamp 1621261055
transform 1 0 24960 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input215
timestamp 1621261055
transform 1 0 24000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_234
timestamp 1621261055
transform 1 0 23616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_242
timestamp 1621261055
transform 1 0 24384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_246
timestamp 1621261055
transform 1 0 24768 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_249
timestamp 1621261055
transform 1 0 25056 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input219
timestamp 1621261055
transform 1 0 25440 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input221
timestamp 1621261055
transform 1 0 26208 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input223
timestamp 1621261055
transform 1 0 26976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_257
timestamp 1621261055
transform 1 0 25824 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_265
timestamp 1621261055
transform 1 0 26592 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_273
timestamp 1621261055
transform 1 0 27360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input226
timestamp 1621261055
transform 1 0 27744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input229
timestamp 1621261055
transform 1 0 28512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input231
timestamp 1621261055
transform 1 0 29280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_281
timestamp 1621261055
transform 1 0 28128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_289
timestamp 1621261055
transform 1 0 28896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_221
timestamp 1621261055
transform 1 0 30240 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input235
timestamp 1621261055
transform 1 0 30720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_297
timestamp 1621261055
transform 1 0 29664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_301
timestamp 1621261055
transform 1 0 30048 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_304
timestamp 1621261055
transform 1 0 30336 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_312
timestamp 1621261055
transform 1 0 31104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input237
timestamp 1621261055
transform 1 0 31488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input240
timestamp 1621261055
transform 1 0 32256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input242
timestamp 1621261055
transform 1 0 33024 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_320
timestamp 1621261055
transform 1 0 31872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_328
timestamp 1621261055
transform 1 0 32640 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_336
timestamp 1621261055
transform 1 0 33408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input244
timestamp 1621261055
transform 1 0 33792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input246
timestamp 1621261055
transform 1 0 34560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_344
timestamp 1621261055
transform 1 0 34176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_352
timestamp 1621261055
transform 1 0 34944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_356
timestamp 1621261055
transform 1 0 35328 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_222
timestamp 1621261055
transform 1 0 35520 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input251
timestamp 1621261055
transform 1 0 36000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input253
timestamp 1621261055
transform 1 0 36768 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_359
timestamp 1621261055
transform 1 0 35616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_367
timestamp 1621261055
transform 1 0 36384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_375
timestamp 1621261055
transform 1 0 37152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input255
timestamp 1621261055
transform 1 0 37536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input257
timestamp 1621261055
transform 1 0 38304 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input259
timestamp 1621261055
transform 1 0 39072 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_383
timestamp 1621261055
transform 1 0 37920 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_391
timestamp 1621261055
transform 1 0 38688 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_399
timestamp 1621261055
transform 1 0 39456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_223
timestamp 1621261055
transform 1 0 40800 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input263
timestamp 1621261055
transform 1 0 39840 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input267
timestamp 1621261055
transform 1 0 41280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_407
timestamp 1621261055
transform 1 0 40224 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_411
timestamp 1621261055
transform 1 0 40608 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_414
timestamp 1621261055
transform 1 0 40896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input269
timestamp 1621261055
transform 1 0 42048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input271
timestamp 1621261055
transform 1 0 42816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_422
timestamp 1621261055
transform 1 0 41664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_430
timestamp 1621261055
transform 1 0 42432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_438
timestamp 1621261055
transform 1 0 43200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input274
timestamp 1621261055
transform 1 0 43584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input276
timestamp 1621261055
transform 1 0 44352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input278
timestamp 1621261055
transform 1 0 45120 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_446
timestamp 1621261055
transform 1 0 43968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_454
timestamp 1621261055
transform 1 0 44736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_462
timestamp 1621261055
transform 1 0 45504 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_224
timestamp 1621261055
transform 1 0 46080 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input282
timestamp 1621261055
transform 1 0 46560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input285
timestamp 1621261055
transform 1 0 47328 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_466
timestamp 1621261055
transform 1 0 45888 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_469
timestamp 1621261055
transform 1 0 46176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_477
timestamp 1621261055
transform 1 0 46944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input287
timestamp 1621261055
transform 1 0 48096 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input289
timestamp 1621261055
transform 1 0 48864 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_485
timestamp 1621261055
transform 1 0 47712 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_493
timestamp 1621261055
transform 1 0 48480 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_501
timestamp 1621261055
transform 1 0 49248 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_225
timestamp 1621261055
transform 1 0 51360 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input290
timestamp 1621261055
transform 1 0 49632 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input292
timestamp 1621261055
transform 1 0 50400 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_509
timestamp 1621261055
transform 1 0 50016 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_517
timestamp 1621261055
transform 1 0 50784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_521
timestamp 1621261055
transform 1 0 51168 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_524
timestamp 1621261055
transform 1 0 51456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input174
timestamp 1621261055
transform 1 0 52128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input175
timestamp 1621261055
transform 1 0 52896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_528
timestamp 1621261055
transform 1 0 51840 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_530
timestamp 1621261055
transform 1 0 52032 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_535
timestamp 1621261055
transform 1 0 52512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_543
timestamp 1621261055
transform 1 0 53280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _014_
timestamp 1621261055
transform -1 0 55488 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input176
timestamp 1621261055
transform 1 0 53664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input179
timestamp 1621261055
transform 1 0 54432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_23
timestamp 1621261055
transform -1 0 55200 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_551
timestamp 1621261055
transform 1 0 54048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_559
timestamp 1621261055
transform 1 0 54816 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_566
timestamp 1621261055
transform 1 0 55488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_226
timestamp 1621261055
transform 1 0 56640 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input63
timestamp 1621261055
transform 1 0 57408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input69
timestamp 1621261055
transform 1 0 55872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_574
timestamp 1621261055
transform 1 0 56256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_579
timestamp 1621261055
transform 1 0 56736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_583
timestamp 1621261055
transform 1 0 57120 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_585
timestamp 1621261055
transform 1 0 57312 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_9
timestamp 1621261055
transform -1 0 58848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_590
timestamp 1621261055
transform 1 0 57792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_594
timestamp 1621261055
transform 1 0 58176 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_596
timestamp 1621261055
transform 1 0 58368 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_10
timestamp 1621261055
transform 1 0 1152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input357
timestamp 1621261055
transform 1 0 3168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input363
timestamp 1621261055
transform 1 0 1536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input364
timestamp 1621261055
transform 1 0 2304 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_8
timestamp 1621261055
transform 1 0 1920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_16
timestamp 1621261055
transform 1 0 2688 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_20
timestamp 1621261055
transform 1 0 3072 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input359
timestamp 1621261055
transform 1 0 3936 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input361
timestamp 1621261055
transform 1 0 4704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_25
timestamp 1621261055
transform 1 0 3552 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_33
timestamp 1621261055
transform 1 0 4320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_41
timestamp 1621261055
transform 1 0 5088 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_227
timestamp 1621261055
transform 1 0 6432 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output575
timestamp 1621261055
transform 1 0 5472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output577
timestamp 1621261055
transform 1 0 6912 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_213
timestamp 1621261055
transform 1 0 6720 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_49
timestamp 1621261055
transform 1 0 5856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_53
timestamp 1621261055
transform 1 0 6240 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_56
timestamp 1621261055
transform 1 0 6528 0 1 5994
box -38 -49 230 715
use AND2X2  AND2X2
timestamp 1624074425
transform 1 0 7680 0 1 5994
box 0 -48 1152 714
use sky130_fd_sc_ls__diode_2  ANTENNA_89
timestamp 1621261055
transform 1 0 7488 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_64
timestamp 1621261055
transform 1 0 7296 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_80
timestamp 1621261055
transform 1 0 8832 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_84
timestamp 1621261055
transform 1 0 9216 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input344
timestamp 1621261055
transform 1 0 9408 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input346
timestamp 1621261055
transform 1 0 10176 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input348
timestamp 1621261055
transform 1 0 10944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_90
timestamp 1621261055
transform 1 0 9792 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_98
timestamp 1621261055
transform 1 0 10560 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_228
timestamp 1621261055
transform 1 0 11712 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input350
timestamp 1621261055
transform 1 0 12192 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input353
timestamp 1621261055
transform 1 0 12960 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_106
timestamp 1621261055
transform 1 0 11328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_111
timestamp 1621261055
transform 1 0 11808 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_119
timestamp 1621261055
transform 1 0 12576 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output444
timestamp 1621261055
transform -1 0 14112 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output494
timestamp 1621261055
transform 1 0 14496 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output505
timestamp 1621261055
transform 1 0 15264 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_96
timestamp 1621261055
transform -1 0 13728 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_147
timestamp 1621261055
transform 1 0 15072 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_127
timestamp 1621261055
transform 1 0 13344 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_135
timestamp 1621261055
transform 1 0 14112 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_143
timestamp 1621261055
transform 1 0 14880 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_229
timestamp 1621261055
transform 1 0 16992 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output527
timestamp 1621261055
transform 1 0 16032 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_111
timestamp 1621261055
transform 1 0 17280 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_151
timestamp 1621261055
transform 1 0 15648 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_159
timestamp 1621261055
transform 1 0 16416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_163
timestamp 1621261055
transform 1 0 16800 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_166
timestamp 1621261055
transform 1 0 17088 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output455
timestamp 1621261055
transform 1 0 17472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output475
timestamp 1621261055
transform 1 0 18240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output477
timestamp 1621261055
transform 1 0 19008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_174
timestamp 1621261055
transform 1 0 17856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_182
timestamp 1621261055
transform 1 0 18624 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output479
timestamp 1621261055
transform 1 0 19776 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output480
timestamp 1621261055
transform 1 0 20544 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output482
timestamp 1621261055
transform 1 0 21312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_133
timestamp 1621261055
transform 1 0 19584 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_190
timestamp 1621261055
transform 1 0 19392 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_198
timestamp 1621261055
transform 1 0 20160 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_206
timestamp 1621261055
transform 1 0 20928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_230
timestamp 1621261055
transform 1 0 22272 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output487
timestamp 1621261055
transform 1 0 22752 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_214
timestamp 1621261055
transform 1 0 21696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_218
timestamp 1621261055
transform 1 0 22080 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_221
timestamp 1621261055
transform 1 0 22368 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_229
timestamp 1621261055
transform 1 0 23136 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output489
timestamp 1621261055
transform 1 0 23520 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output491
timestamp 1621261055
transform 1 0 24288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_237
timestamp 1621261055
transform 1 0 23904 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_245
timestamp 1621261055
transform 1 0 24672 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input222
timestamp 1621261055
transform 1 0 25632 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input225
timestamp 1621261055
transform 1 0 26784 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_253
timestamp 1621261055
transform 1 0 25440 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_259
timestamp 1621261055
transform 1 0 26016 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_5_271
timestamp 1621261055
transform 1 0 27168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_231
timestamp 1621261055
transform 1 0 27552 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output501
timestamp 1621261055
transform 1 0 28032 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output504
timestamp 1621261055
transform 1 0 28800 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_143
timestamp 1621261055
transform 1 0 27840 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_145
timestamp 1621261055
transform 1 0 28608 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_276
timestamp 1621261055
transform 1 0 27648 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_284
timestamp 1621261055
transform 1 0 28416 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_292
timestamp 1621261055
transform 1 0 29184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input234
timestamp 1621261055
transform 1 0 29664 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input238
timestamp 1621261055
transform 1 0 31200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output509
timestamp 1621261055
transform 1 0 30432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_151
timestamp 1621261055
transform 1 0 30240 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_296
timestamp 1621261055
transform 1 0 29568 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_301
timestamp 1621261055
transform 1 0 30048 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_309
timestamp 1621261055
transform 1 0 30816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_317
timestamp 1621261055
transform 1 0 31584 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_155
timestamp 1621261055
transform -1 0 31968 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output513
timestamp 1621261055
transform -1 0 32352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_329
timestamp 1621261055
transform 1 0 32736 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_327
timestamp 1621261055
transform 1 0 32544 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_156
timestamp 1621261055
transform -1 0 32544 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_331
timestamp 1621261055
transform 1 0 32928 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_166
timestamp 1621261055
transform -1 0 33312 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_232
timestamp 1621261055
transform 1 0 32832 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output518
timestamp 1621261055
transform -1 0 33696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output520
timestamp 1621261055
transform 1 0 34080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output522
timestamp 1621261055
transform -1 0 35232 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_167
timestamp 1621261055
transform -1 0 33888 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_173
timestamp 1621261055
transform -1 0 34848 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_341
timestamp 1621261055
transform 1 0 33888 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_347
timestamp 1621261055
transform 1 0 34464 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_355
timestamp 1621261055
transform 1 0 35232 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input254
timestamp 1621261055
transform 1 0 36288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output529
timestamp 1621261055
transform -1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_177
timestamp 1621261055
transform -1 0 37056 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_363
timestamp 1621261055
transform 1 0 36000 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_365
timestamp 1621261055
transform 1 0 36192 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_370
timestamp 1621261055
transform 1 0 36672 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_378
timestamp 1621261055
transform 1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_233
timestamp 1621261055
transform 1 0 38112 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input262
timestamp 1621261055
transform 1 0 38880 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_382
timestamp 1621261055
transform 1 0 37824 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_384
timestamp 1621261055
transform 1 0 38016 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_386
timestamp 1621261055
transform 1 0 38208 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_390
timestamp 1621261055
transform 1 0 38592 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_392
timestamp 1621261055
transform 1 0 38784 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_5_397
timestamp 1621261055
transform 1 0 39264 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input266
timestamp 1621261055
transform 1 0 40320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output540
timestamp 1621261055
transform 1 0 41088 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_405
timestamp 1621261055
transform 1 0 40032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_407
timestamp 1621261055
transform 1 0 40224 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_412
timestamp 1621261055
transform 1 0 40704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_420
timestamp 1621261055
transform 1 0 41472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_234
timestamp 1621261055
transform 1 0 43392 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input270
timestamp 1621261055
transform 1 0 41856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output544
timestamp 1621261055
transform -1 0 43008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_181
timestamp 1621261055
transform -1 0 42624 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_428
timestamp 1621261055
transform 1 0 42240 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_436
timestamp 1621261055
transform 1 0 43008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_441
timestamp 1621261055
transform 1 0 43488 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input281
timestamp 1621261055
transform 1 0 45504 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output548
timestamp 1621261055
transform -1 0 44256 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output552
timestamp 1621261055
transform -1 0 45024 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_183
timestamp 1621261055
transform -1 0 43872 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_187
timestamp 1621261055
transform -1 0 44640 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_449
timestamp 1621261055
transform 1 0 44256 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_457
timestamp 1621261055
transform 1 0 45024 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_461
timestamp 1621261055
transform 1 0 45408 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _068_
timestamp 1621261055
transform -1 0 46560 0 1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input286
timestamp 1621261055
transform 1 0 46944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_110
timestamp 1621261055
transform -1 0 46272 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_466
timestamp 1621261055
transform 1 0 45888 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_473
timestamp 1621261055
transform 1 0 46560 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_481
timestamp 1621261055
transform 1 0 47328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_235
timestamp 1621261055
transform 1 0 48672 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input288
timestamp 1621261055
transform 1 0 47712 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input291
timestamp 1621261055
transform 1 0 49152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_489
timestamp 1621261055
transform 1 0 48096 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_493
timestamp 1621261055
transform 1 0 48480 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_496
timestamp 1621261055
transform 1 0 48768 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_504
timestamp 1621261055
transform 1 0 49536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input293
timestamp 1621261055
transform 1 0 49920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output445
timestamp 1621261055
transform 1 0 50688 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output447
timestamp 1621261055
transform -1 0 51840 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_100
timestamp 1621261055
transform -1 0 51456 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_512
timestamp 1621261055
transform 1 0 50304 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_520
timestamp 1621261055
transform 1 0 51072 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input192
timestamp 1621261055
transform 1 0 53184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output448
timestamp 1621261055
transform -1 0 52608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_102
timestamp 1621261055
transform -1 0 52224 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_528
timestamp 1621261055
transform 1 0 51840 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_536
timestamp 1621261055
transform 1 0 52608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_540
timestamp 1621261055
transform 1 0 52992 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_546
timestamp 1621261055
transform 1 0 53568 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_236
timestamp 1621261055
transform 1 0 53952 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input180
timestamp 1621261055
transform 1 0 54432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input181
timestamp 1621261055
transform 1 0 55200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_551
timestamp 1621261055
transform 1 0 54048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_559
timestamp 1621261055
transform 1 0 54816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_567
timestamp 1621261055
transform 1 0 55584 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input67
timestamp 1621261055
transform 1 0 56928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input183
timestamp 1621261055
transform 1 0 55968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_575
timestamp 1621261055
transform 1 0 56352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_579
timestamp 1621261055
transform 1 0 56736 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_585
timestamp 1621261055
transform 1 0 57312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_11
timestamp 1621261055
transform -1 0 58848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input65
timestamp 1621261055
transform 1 0 57696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_593
timestamp 1621261055
transform 1 0 58080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_12
timestamp 1621261055
transform 1 0 1152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input365
timestamp 1621261055
transform 1 0 2496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input366
timestamp 1621261055
transform 1 0 1536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_8
timestamp 1621261055
transform 1 0 1920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_12
timestamp 1621261055
transform 1 0 2304 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_18
timestamp 1621261055
transform 1 0 2880 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_237
timestamp 1621261055
transform 1 0 3840 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output598
timestamp 1621261055
transform 1 0 4320 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output601
timestamp 1621261055
transform 1 0 5088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_237
timestamp 1621261055
transform 1 0 4896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_26
timestamp 1621261055
transform 1 0 3648 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_29
timestamp 1621261055
transform 1 0 3936 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_37
timestamp 1621261055
transform 1 0 4704 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output576
timestamp 1621261055
transform 1 0 5856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output578
timestamp 1621261055
transform 1 0 6624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_215
timestamp 1621261055
transform 1 0 6432 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_45
timestamp 1621261055
transform 1 0 5472 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_53
timestamp 1621261055
transform 1 0 6240 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_61
timestamp 1621261055
transform 1 0 7008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_238
timestamp 1621261055
transform 1 0 9120 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output579
timestamp 1621261055
transform 1 0 7392 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output580
timestamp 1621261055
transform 1 0 8160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_217
timestamp 1621261055
transform 1 0 7968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_69
timestamp 1621261055
transform 1 0 7776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_77
timestamp 1621261055
transform 1 0 8544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_81
timestamp 1621261055
transform 1 0 8928 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_84
timestamp 1621261055
transform 1 0 9216 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input349
timestamp 1621261055
transform 1 0 11232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output582
timestamp 1621261055
transform 1 0 9600 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output585
timestamp 1621261055
transform 1 0 10368 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_223
timestamp 1621261055
transform 1 0 10176 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_92
timestamp 1621261055
transform 1 0 9984 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_100
timestamp 1621261055
transform 1 0 10752 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_104
timestamp 1621261055
transform 1 0 11136 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _033_
timestamp 1621261055
transform 1 0 12000 0 -1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input354
timestamp 1621261055
transform 1 0 12672 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_20
timestamp 1621261055
transform 1 0 11808 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_109
timestamp 1621261055
transform 1 0 11616 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_116
timestamp 1621261055
transform 1 0 12288 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_124
timestamp 1621261055
transform 1 0 13056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_239
timestamp 1621261055
transform 1 0 14400 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output483
timestamp 1621261055
transform 1 0 13440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output516
timestamp 1621261055
transform 1 0 14880 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_132
timestamp 1621261055
transform 1 0 13824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_136
timestamp 1621261055
transform 1 0 14208 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_139
timestamp 1621261055
transform 1 0 14496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_147
timestamp 1621261055
transform 1 0 15264 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output466
timestamp 1621261055
transform 1 0 17088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output538
timestamp 1621261055
transform 1 0 15648 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_155
timestamp 1621261055
transform 1 0 16032 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_163
timestamp 1621261055
transform 1 0 16800 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_165
timestamp 1621261055
transform 1 0 16992 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output476
timestamp 1621261055
transform 1 0 17856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output478
timestamp 1621261055
transform 1 0 18624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_129
timestamp 1621261055
transform 1 0 17664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_131
timestamp 1621261055
transform 1 0 18432 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_170
timestamp 1621261055
transform 1 0 17472 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_178
timestamp 1621261055
transform 1 0 18240 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_186
timestamp 1621261055
transform 1 0 19008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_240
timestamp 1621261055
transform 1 0 19680 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output481
timestamp 1621261055
transform 1 0 20160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output484
timestamp 1621261055
transform 1 0 20928 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_135
timestamp 1621261055
transform 1 0 19968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_190
timestamp 1621261055
transform 1 0 19392 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_192
timestamp 1621261055
transform 1 0 19584 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_194
timestamp 1621261055
transform 1 0 19776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_202
timestamp 1621261055
transform 1 0 20544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_210
timestamp 1621261055
transform 1 0 21312 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output486
timestamp 1621261055
transform 1 0 21696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output488
timestamp 1621261055
transform 1 0 22464 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output490
timestamp 1621261055
transform 1 0 23232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_137
timestamp 1621261055
transform 1 0 21504 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_218
timestamp 1621261055
transform 1 0 22080 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_226
timestamp 1621261055
transform 1 0 22848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_241
timestamp 1621261055
transform 1 0 24960 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output492
timestamp 1621261055
transform 1 0 24000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_139
timestamp 1621261055
transform 1 0 25248 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_234
timestamp 1621261055
transform 1 0 23616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_242
timestamp 1621261055
transform 1 0 24384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_246
timestamp 1621261055
transform 1 0 24768 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_249
timestamp 1621261055
transform 1 0 25056 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output496
timestamp 1621261055
transform 1 0 25440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output498
timestamp 1621261055
transform 1 0 26208 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output500
timestamp 1621261055
transform 1 0 26976 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_257
timestamp 1621261055
transform 1 0 25824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_265
timestamp 1621261055
transform 1 0 26592 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_273
timestamp 1621261055
transform 1 0 27360 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output503
timestamp 1621261055
transform 1 0 27744 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output506
timestamp 1621261055
transform 1 0 28512 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output508
timestamp 1621261055
transform 1 0 29280 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_281
timestamp 1621261055
transform 1 0 28128 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_289
timestamp 1621261055
transform 1 0 28896 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_242
timestamp 1621261055
transform 1 0 30240 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output512
timestamp 1621261055
transform 1 0 30720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_158
timestamp 1621261055
transform -1 0 31488 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_297
timestamp 1621261055
transform 1 0 29664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_301
timestamp 1621261055
transform 1 0 30048 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_304
timestamp 1621261055
transform 1 0 30336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_312
timestamp 1621261055
transform 1 0 31104 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output514
timestamp 1621261055
transform -1 0 31872 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output517
timestamp 1621261055
transform 1 0 32256 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output519
timestamp 1621261055
transform 1 0 33024 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_159
timestamp 1621261055
transform -1 0 32064 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_164
timestamp 1621261055
transform 1 0 32064 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_169
timestamp 1621261055
transform 1 0 32832 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_328
timestamp 1621261055
transform 1 0 32640 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_336
timestamp 1621261055
transform 1 0 33408 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output521
timestamp 1621261055
transform 1 0 33792 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output524
timestamp 1621261055
transform 1 0 34560 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_171
timestamp 1621261055
transform 1 0 33600 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_344
timestamp 1621261055
transform 1 0 34176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_352
timestamp 1621261055
transform 1 0 34944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_356
timestamp 1621261055
transform 1 0 35328 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_243
timestamp 1621261055
transform 1 0 35520 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output528
timestamp 1621261055
transform 1 0 36000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output531
timestamp 1621261055
transform 1 0 36768 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_359
timestamp 1621261055
transform 1 0 35616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_367
timestamp 1621261055
transform 1 0 36384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_375
timestamp 1621261055
transform 1 0 37152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output533
timestamp 1621261055
transform 1 0 37536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output534
timestamp 1621261055
transform 1 0 38304 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output535
timestamp 1621261055
transform 1 0 39072 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_383
timestamp 1621261055
transform 1 0 37920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_391
timestamp 1621261055
transform 1 0 38688 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_399
timestamp 1621261055
transform 1 0 39456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_244
timestamp 1621261055
transform 1 0 40800 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output537
timestamp 1621261055
transform 1 0 39840 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output542
timestamp 1621261055
transform 1 0 41280 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_179
timestamp 1621261055
transform 1 0 41088 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_407
timestamp 1621261055
transform 1 0 40224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_411
timestamp 1621261055
transform 1 0 40608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_414
timestamp 1621261055
transform 1 0 40896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output545
timestamp 1621261055
transform 1 0 42048 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output547
timestamp 1621261055
transform 1 0 42816 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_422
timestamp 1621261055
transform 1 0 41664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_430
timestamp 1621261055
transform 1 0 42432 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_438
timestamp 1621261055
transform 1 0 43200 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output551
timestamp 1621261055
transform 1 0 43584 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output553
timestamp 1621261055
transform -1 0 44736 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output555
timestamp 1621261055
transform 1 0 45120 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_189
timestamp 1621261055
transform -1 0 44352 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_446
timestamp 1621261055
transform 1 0 43968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_454
timestamp 1621261055
transform 1 0 44736 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_462
timestamp 1621261055
transform 1 0 45504 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_245
timestamp 1621261055
transform 1 0 46080 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output558
timestamp 1621261055
transform -1 0 46944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output561
timestamp 1621261055
transform -1 0 47712 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_195
timestamp 1621261055
transform -1 0 46560 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_198
timestamp 1621261055
transform -1 0 47328 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_466
timestamp 1621261055
transform 1 0 45888 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_469
timestamp 1621261055
transform 1 0 46176 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_477
timestamp 1621261055
transform 1 0 46944 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output563
timestamp 1621261055
transform 1 0 48096 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output565
timestamp 1621261055
transform 1 0 48864 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_485
timestamp 1621261055
transform 1 0 47712 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_493
timestamp 1621261055
transform 1 0 48480 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_501
timestamp 1621261055
transform 1 0 49248 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_246
timestamp 1621261055
transform 1 0 51360 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output446
timestamp 1621261055
transform -1 0 50496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_98
timestamp 1621261055
transform -1 0 50112 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_505
timestamp 1621261055
transform 1 0 49632 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_507
timestamp 1621261055
transform 1 0 49824 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_6_514
timestamp 1621261055
transform 1 0 50496 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_6_522
timestamp 1621261055
transform 1 0 51264 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_524
timestamp 1621261055
transform 1 0 51456 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output449
timestamp 1621261055
transform -1 0 52224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output451
timestamp 1621261055
transform 1 0 52608 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_104
timestamp 1621261055
transform -1 0 51840 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_532
timestamp 1621261055
transform 1 0 52224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_540
timestamp 1621261055
transform 1 0 52992 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input182
timestamp 1621261055
transform 1 0 54720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input184
timestamp 1621261055
transform 1 0 55488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input196
timestamp 1621261055
transform 1 0 53952 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_548
timestamp 1621261055
transform 1 0 53760 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_554
timestamp 1621261055
transform 1 0 54336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_562
timestamp 1621261055
transform 1 0 55104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_247
timestamp 1621261055
transform 1 0 56640 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_6_570
timestamp 1621261055
transform 1 0 55872 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_6_579
timestamp 1621261055
transform 1 0 56736 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_587
timestamp 1621261055
transform 1 0 57504 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_13
timestamp 1621261055
transform -1 0 58848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input66
timestamp 1621261055
transform 1 0 57696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_593
timestamp 1621261055
transform 1 0 58080 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output572
timestamp 1621261055
transform 1 0 1536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input367
timestamp 1621261055
transform 1 0 1536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_16
timestamp 1621261055
transform 1 0 1152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_14
timestamp 1621261055
transform 1 0 1152 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_8
timestamp 1621261055
transform 1 0 1920 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_207
timestamp 1621261055
transform 1 0 1920 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_221
timestamp 1621261055
transform 1 0 2112 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_209
timestamp 1621261055
transform 1 0 2112 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output584
timestamp 1621261055
transform 1 0 2304 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output573
timestamp 1621261055
transform 1 0 2304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_16
timestamp 1621261055
transform 1 0 2688 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_16
timestamp 1621261055
transform 1 0 2688 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output599
timestamp 1621261055
transform 1 0 3072 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output595
timestamp 1621261055
transform 1 0 3072 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_24
timestamp 1621261055
transform 1 0 3456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_24
timestamp 1621261055
transform 1 0 3456 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_29
timestamp 1621261055
transform 1 0 3936 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_235
timestamp 1621261055
transform 1 0 3648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output600
timestamp 1621261055
transform 1 0 3840 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_258
timestamp 1621261055
transform 1 0 3840 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_32
timestamp 1621261055
transform 1 0 4224 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output603
timestamp 1621261055
transform 1 0 4320 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_37
timestamp 1621261055
transform 1 0 4704 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_40
timestamp 1621261055
transform 1 0 4992 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output602
timestamp 1621261055
transform 1 0 4608 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_41
timestamp 1621261055
transform 1 0 5088 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_239
timestamp 1621261055
transform 1 0 5184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_49
timestamp 1621261055
transform 1 0 5856 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_43
timestamp 1621261055
transform 1 0 5280 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_48
timestamp 1621261055
transform 1 0 5760 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_2
timestamp 1621261055
transform -1 0 5568 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output604
timestamp 1621261055
transform 1 0 5376 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _001_
timestamp 1621261055
transform -1 0 5856 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_57
timestamp 1621261055
transform 1 0 6624 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_56
timestamp 1621261055
transform 1 0 6528 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_54
timestamp 1621261055
transform 1 0 6336 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_52
timestamp 1621261055
transform 1 0 6144 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_248
timestamp 1621261055
transform 1 0 6432 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_72
timestamp 1621261055
transform 1 0 8064 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_67
timestamp 1621261055
transform 1 0 7584 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_65
timestamp 1621261055
transform 1 0 7392 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_64
timestamp 1621261055
transform 1 0 7296 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_93
timestamp 1621261055
transform 1 0 7488 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output581
timestamp 1621261055
transform 1 0 7680 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_84
timestamp 1621261055
transform 1 0 9216 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_82
timestamp 1621261055
transform 1 0 9024 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_80
timestamp 1621261055
transform 1 0 8832 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_80
timestamp 1621261055
transform 1 0 8832 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_219
timestamp 1621261055
transform 1 0 9024 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output583
timestamp 1621261055
transform 1 0 9216 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_259
timestamp 1621261055
transform 1 0 9120 0 -1 8658
box -38 -49 134 715
use AOI21X1  AOI21X1
timestamp 1624074425
transform 1 0 7680 0 1 7326
box 0 -48 1152 714
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_88
timestamp 1621261055
transform 1 0 9600 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_227
timestamp 1621261055
transform -1 0 9600 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output587
timestamp 1621261055
transform -1 0 9984 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_92
timestamp 1621261055
transform 1 0 9984 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_225
timestamp 1621261055
transform 1 0 9792 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output586
timestamp 1621261055
transform 1 0 9984 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_96
timestamp 1621261055
transform 1 0 10368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output589
timestamp 1621261055
transform 1 0 10368 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_100
timestamp 1621261055
transform 1 0 10752 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output588
timestamp 1621261055
transform 1 0 10752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_104
timestamp 1621261055
transform 1 0 11136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output590
timestamp 1621261055
transform 1 0 11136 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_108
timestamp 1621261055
transform 1 0 11520 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_108
timestamp 1621261055
transform 1 0 11520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_111
timestamp 1621261055
transform 1 0 11808 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_229
timestamp 1621261055
transform -1 0 12192 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output592
timestamp 1621261055
transform 1 0 11904 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_249
timestamp 1621261055
transform 1 0 11712 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_116
timestamp 1621261055
transform 1 0 12288 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_119
timestamp 1621261055
transform 1 0 12576 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_231
timestamp 1621261055
transform 1 0 12480 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output591
timestamp 1621261055
transform -1 0 12576 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_124
timestamp 1621261055
transform 1 0 13056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output594
timestamp 1621261055
transform 1 0 12672 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output593
timestamp 1621261055
transform 1 0 12960 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_132
timestamp 1621261055
transform 1 0 13824 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_127
timestamp 1621261055
transform 1 0 13344 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_233
timestamp 1621261055
transform 1 0 13536 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output597
timestamp 1621261055
transform 1 0 13440 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output596
timestamp 1621261055
transform 1 0 13728 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_139
timestamp 1621261055
transform 1 0 14496 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_136
timestamp 1621261055
transform 1 0 14208 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_143
timestamp 1621261055
transform 1 0 14880 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_135
timestamp 1621261055
transform 1 0 14112 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_260
timestamp 1621261055
transform 1 0 14400 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_147
timestamp 1621261055
transform 1 0 15264 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_147
timestamp 1621261055
transform 1 0 15264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_155
timestamp 1621261055
transform 1 0 16032 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_185
timestamp 1621261055
transform -1 0 15648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output560
timestamp 1621261055
transform 1 0 16032 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output549
timestamp 1621261055
transform -1 0 16032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_159
timestamp 1621261055
transform 1 0 16416 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_163
timestamp 1621261055
transform 1 0 16800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output571
timestamp 1621261055
transform 1 0 16800 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_167
timestamp 1621261055
transform 1 0 17184 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_166
timestamp 1621261055
transform 1 0 17088 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_250
timestamp 1621261055
transform 1 0 16992 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_7_174
timestamp 1621261055
transform 1 0 17856 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_182
timestamp 1621261055
transform 1 0 18624 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_175
timestamp 1621261055
transform 1 0 17952 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_183
timestamp 1621261055
transform 1 0 18720 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_194
timestamp 1621261055
transform 1 0 19776 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_191
timestamp 1621261055
transform 1 0 19488 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_190
timestamp 1621261055
transform 1 0 19392 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_261
timestamp 1621261055
transform 1 0 19680 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_202
timestamp 1621261055
transform 1 0 20544 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_202
timestamp 1621261055
transform 1 0 20544 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_198
timestamp 1621261055
transform 1 0 20160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output485
timestamp 1621261055
transform 1 0 20736 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_210
timestamp 1621261055
transform 1 0 21312 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_208
timestamp 1621261055
transform 1 0 21120 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_251
timestamp 1621261055
transform 1 0 22272 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_216
timestamp 1621261055
transform 1 0 21888 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_221
timestamp 1621261055
transform 1 0 22368 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_229
timestamp 1621261055
transform 1 0 23136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_218
timestamp 1621261055
transform 1 0 22080 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_226
timestamp 1621261055
transform 1 0 22848 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_234
timestamp 1621261055
transform 1 0 23616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_239
timestamp 1621261055
transform 1 0 24096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_233
timestamp 1621261055
transform 1 0 23520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output493
timestamp 1621261055
transform 1 0 23712 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_246
timestamp 1621261055
transform 1 0 24768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_242
timestamp 1621261055
transform 1 0 24384 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_247
timestamp 1621261055
transform 1 0 24864 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output495
timestamp 1621261055
transform 1 0 24480 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_262
timestamp 1621261055
transform 1 0 24960 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_249
timestamp 1621261055
transform 1 0 25056 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output497
timestamp 1621261055
transform 1 0 25248 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output499
timestamp 1621261055
transform -1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output502
timestamp 1621261055
transform 1 0 26784 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_141
timestamp 1621261055
transform -1 0 26016 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_255
timestamp 1621261055
transform 1 0 25632 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_263
timestamp 1621261055
transform 1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_271
timestamp 1621261055
transform 1 0 27168 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_257
timestamp 1621261055
transform 1 0 25824 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_265
timestamp 1621261055
transform 1 0 26592 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_273
timestamp 1621261055
transform 1 0 27360 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_281
timestamp 1621261055
transform 1 0 28128 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_278
timestamp 1621261055
transform 1 0 27840 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_276
timestamp 1621261055
transform 1 0 27648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_149
timestamp 1621261055
transform -1 0 28128 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output507
timestamp 1621261055
transform -1 0 28512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_252
timestamp 1621261055
transform 1 0 27552 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_289
timestamp 1621261055
transform 1 0 28896 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_289
timestamp 1621261055
transform 1 0 28896 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_285
timestamp 1621261055
transform 1 0 28512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_153
timestamp 1621261055
transform 1 0 28992 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_293
timestamp 1621261055
transform 1 0 29280 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output510
timestamp 1621261055
transform 1 0 29184 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_299
timestamp 1621261055
transform 1 0 29856 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_295
timestamp 1621261055
transform 1 0 29472 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_296
timestamp 1621261055
transform 1 0 29568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output511
timestamp 1621261055
transform 1 0 29952 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _177_
timestamp 1621261055
transform 1 0 29568 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_311
timestamp 1621261055
transform 1 0 31008 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_8_304
timestamp 1621261055
transform 1 0 30336 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_308
timestamp 1621261055
transform 1 0 30720 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_304
timestamp 1621261055
transform 1 0 30336 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_161
timestamp 1621261055
transform -1 0 31008 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output515
timestamp 1621261055
transform -1 0 31392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_263
timestamp 1621261055
transform 1 0 30240 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _119_
timestamp 1621261055
transform 1 0 30720 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_162
timestamp 1621261055
transform -1 0 31584 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_253
timestamp 1621261055
transform 1 0 32832 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_7_317
timestamp 1621261055
transform 1 0 31584 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_325
timestamp 1621261055
transform 1 0 32352 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_329
timestamp 1621261055
transform 1 0 32736 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_331
timestamp 1621261055
transform 1 0 32928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_335
timestamp 1621261055
transform 1 0 33312 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_319
timestamp 1621261055
transform 1 0 31776 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_327
timestamp 1621261055
transform 1 0 32544 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_335
timestamp 1621261055
transform 1 0 33312 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_337
timestamp 1621261055
transform 1 0 33504 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output523
timestamp 1621261055
transform 1 0 33600 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_343
timestamp 1621261055
transform 1 0 34080 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_342
timestamp 1621261055
transform 1 0 33984 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_175
timestamp 1621261055
transform 1 0 34176 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _096_
timestamp 1621261055
transform 1 0 34176 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_8_347
timestamp 1621261055
transform 1 0 34464 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_350
timestamp 1621261055
transform 1 0 34752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output525
timestamp 1621261055
transform 1 0 34368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_354
timestamp 1621261055
transform 1 0 35136 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output526
timestamp 1621261055
transform 1 0 35136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _124_
timestamp 1621261055
transform 1 0 34848 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_264
timestamp 1621261055
transform 1 0 35520 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output530
timestamp 1621261055
transform 1 0 35904 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output532
timestamp 1621261055
transform 1 0 36672 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_358
timestamp 1621261055
transform 1 0 35520 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_366
timestamp 1621261055
transform 1 0 36288 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_374
timestamp 1621261055
transform 1 0 37056 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_359
timestamp 1621261055
transform 1 0 35616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_367
timestamp 1621261055
transform 1 0 36384 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_375
timestamp 1621261055
transform 1 0 37152 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_383
timestamp 1621261055
transform 1 0 37920 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_386
timestamp 1621261055
transform 1 0 38208 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_384
timestamp 1621261055
transform 1 0 38016 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_382
timestamp 1621261055
transform 1 0 37824 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_254
timestamp 1621261055
transform 1 0 38112 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_391
timestamp 1621261055
transform 1 0 38688 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_394
timestamp 1621261055
transform 1 0 38976 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output536
timestamp 1621261055
transform 1 0 38592 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_399
timestamp 1621261055
transform 1 0 39456 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output539
timestamp 1621261055
transform 1 0 39360 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_265
timestamp 1621261055
transform 1 0 40800 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output541
timestamp 1621261055
transform 1 0 40128 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output543
timestamp 1621261055
transform 1 0 40896 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_402
timestamp 1621261055
transform 1 0 39744 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_410
timestamp 1621261055
transform 1 0 40512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_418
timestamp 1621261055
transform 1 0 41280 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_407
timestamp 1621261055
transform 1 0 40224 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_411
timestamp 1621261055
transform 1 0 40608 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_414
timestamp 1621261055
transform 1 0 40896 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_422
timestamp 1621261055
transform 1 0 41664 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_426
timestamp 1621261055
transform 1 0 42048 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output546
timestamp 1621261055
transform 1 0 41664 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_430
timestamp 1621261055
transform 1 0 42432 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_434
timestamp 1621261055
transform 1 0 42816 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output550
timestamp 1621261055
transform 1 0 42432 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_438
timestamp 1621261055
transform 1 0 43200 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_441
timestamp 1621261055
transform 1 0 43488 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_438
timestamp 1621261055
transform 1 0 43200 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_255
timestamp 1621261055
transform 1 0 43392 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_446
timestamp 1621261055
transform 1 0 43968 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_449
timestamp 1621261055
transform 1 0 44256 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output554
timestamp 1621261055
transform 1 0 43872 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_454
timestamp 1621261055
transform 1 0 44736 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_457
timestamp 1621261055
transform 1 0 45024 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_191
timestamp 1621261055
transform -1 0 44640 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output556
timestamp 1621261055
transform -1 0 45024 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_462
timestamp 1621261055
transform 1 0 45504 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_193
timestamp 1621261055
transform -1 0 45408 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output557
timestamp 1621261055
transform -1 0 45792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_469
timestamp 1621261055
transform 1 0 46176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_466
timestamp 1621261055
transform 1 0 45888 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_465
timestamp 1621261055
transform 1 0 45792 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_197
timestamp 1621261055
transform -1 0 46176 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output559
timestamp 1621261055
transform -1 0 46560 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_266
timestamp 1621261055
transform 1 0 46080 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_477
timestamp 1621261055
transform 1 0 46944 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_473
timestamp 1621261055
transform 1 0 46560 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_199
timestamp 1621261055
transform -1 0 46944 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output562
timestamp 1621261055
transform -1 0 47328 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_481
timestamp 1621261055
transform 1 0 47328 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_200
timestamp 1621261055
transform -1 0 47712 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_485
timestamp 1621261055
transform 1 0 47712 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_202
timestamp 1621261055
transform -1 0 48000 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output566
timestamp 1621261055
transform -1 0 48384 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output564
timestamp 1621261055
transform -1 0 48096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_492
timestamp 1621261055
transform 1 0 48384 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_489
timestamp 1621261055
transform 1 0 48096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_496
timestamp 1621261055
transform 1 0 48768 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_493
timestamp 1621261055
transform 1 0 48480 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_205
timestamp 1621261055
transform -1 0 48768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output568
timestamp 1621261055
transform -1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_256
timestamp 1621261055
transform 1 0 48672 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_500
timestamp 1621261055
transform 1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_204
timestamp 1621261055
transform -1 0 49152 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output567
timestamp 1621261055
transform -1 0 49536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_504
timestamp 1621261055
transform 1 0 49536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output570
timestamp 1621261055
transform 1 0 49536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_508
timestamp 1621261055
transform 1 0 49920 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output569
timestamp 1621261055
transform 1 0 49920 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_512
timestamp 1621261055
transform 1 0 50304 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_512
timestamp 1621261055
transform 1 0 50304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_516
timestamp 1621261055
transform 1 0 50688 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_10
timestamp 1621261055
transform -1 0 50688 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output473
timestamp 1621261055
transform 1 0 50880 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _029_
timestamp 1621261055
transform -1 0 50976 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_8_519
timestamp 1621261055
transform 1 0 50976 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_522
timestamp 1621261055
transform 1 0 51264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_267
timestamp 1621261055
transform 1 0 51360 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_524
timestamp 1621261055
transform 1 0 51456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_106
timestamp 1621261055
transform -1 0 51648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_530
timestamp 1621261055
transform 1 0 52032 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_528
timestamp 1621261055
transform 1 0 51840 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_530
timestamp 1621261055
transform 1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output450
timestamp 1621261055
transform -1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_126
timestamp 1621261055
transform -1 0 52320 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output472
timestamp 1621261055
transform -1 0 52704 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output452
timestamp 1621261055
transform 1 0 52416 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_537
timestamp 1621261055
transform 1 0 52704 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_538
timestamp 1621261055
transform 1 0 52800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_109
timestamp 1621261055
transform -1 0 53088 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_108
timestamp 1621261055
transform -1 0 53184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output454
timestamp 1621261055
transform -1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output453
timestamp 1621261055
transform -1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_545
timestamp 1621261055
transform 1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_546
timestamp 1621261055
transform 1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_553
timestamp 1621261055
transform 1 0 54240 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_551
timestamp 1621261055
transform 1 0 54048 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output456
timestamp 1621261055
transform 1 0 53856 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_257
timestamp 1621261055
transform 1 0 53952 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_561
timestamp 1621261055
transform 1 0 55008 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_559
timestamp 1621261055
transform 1 0 54816 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input197
timestamp 1621261055
transform 1 0 55104 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input194
timestamp 1621261055
transform 1 0 55008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_566
timestamp 1621261055
transform 1 0 55488 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_565
timestamp 1621261055
transform 1 0 55392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_574
timestamp 1621261055
transform 1 0 56256 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_573
timestamp 1621261055
transform 1 0 56160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input193
timestamp 1621261055
transform 1 0 55872 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input185
timestamp 1621261055
transform 1 0 55776 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_579
timestamp 1621261055
transform 1 0 56736 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_581
timestamp 1621261055
transform 1 0 56928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input188
timestamp 1621261055
transform 1 0 57120 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input186
timestamp 1621261055
transform 1 0 56544 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_268
timestamp 1621261055
transform 1 0 56640 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_587
timestamp 1621261055
transform 1 0 57504 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input187
timestamp 1621261055
transform 1 0 57312 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_15
timestamp 1621261055
transform -1 0 58848 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_17
timestamp 1621261055
transform -1 0 58848 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_589
timestamp 1621261055
transform 1 0 57696 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_595
timestamp 1621261055
transform 1 0 58272 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_18
timestamp 1621261055
transform 1 0 1152 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_4
timestamp 1621261055
transform 1 0 1536 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_12
timestamp 1621261055
transform 1 0 2304 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_20
timestamp 1621261055
transform 1 0 3072 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _144_
timestamp 1621261055
transform 1 0 4512 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_9_28
timestamp 1621261055
transform 1 0 3840 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_32
timestamp 1621261055
transform 1 0 4224 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_34
timestamp 1621261055
transform 1 0 4416 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_38
timestamp 1621261055
transform 1 0 4800 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_269
timestamp 1621261055
transform 1 0 6432 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_46
timestamp 1621261055
transform 1 0 5568 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_9_54
timestamp 1621261055
transform 1 0 6336 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_56
timestamp 1621261055
transform 1 0 6528 0 1 8658
box -38 -49 806 715
use AOI22X1  AOI22X1
timestamp 1624074425
transform 1 0 7680 0 1 8658
box 0 -48 1440 714
use sky130_fd_sc_ls__diode_2  ANTENNA_43
timestamp 1621261055
transform 1 0 7488 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_64
timestamp 1621261055
transform 1 0 7296 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_83
timestamp 1621261055
transform 1 0 9120 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_91
timestamp 1621261055
transform 1 0 9888 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_99
timestamp 1621261055
transform 1 0 10656 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_270
timestamp 1621261055
transform 1 0 11712 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_107
timestamp 1621261055
transform 1 0 11424 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_109
timestamp 1621261055
transform 1 0 11616 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_111
timestamp 1621261055
transform 1 0 11808 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_119
timestamp 1621261055
transform 1 0 12576 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_127
timestamp 1621261055
transform 1 0 13344 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_135
timestamp 1621261055
transform 1 0 14112 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_143
timestamp 1621261055
transform 1 0 14880 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_271
timestamp 1621261055
transform 1 0 16992 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_151
timestamp 1621261055
transform 1 0 15648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_159
timestamp 1621261055
transform 1 0 16416 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_163
timestamp 1621261055
transform 1 0 16800 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_166
timestamp 1621261055
transform 1 0 17088 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_174
timestamp 1621261055
transform 1 0 17856 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_182
timestamp 1621261055
transform 1 0 18624 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_190
timestamp 1621261055
transform 1 0 19392 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_198
timestamp 1621261055
transform 1 0 20160 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_206
timestamp 1621261055
transform 1 0 20928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_272
timestamp 1621261055
transform 1 0 22272 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_214
timestamp 1621261055
transform 1 0 21696 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_218
timestamp 1621261055
transform 1 0 22080 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_221
timestamp 1621261055
transform 1 0 22368 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_229
timestamp 1621261055
transform 1 0 23136 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_237
timestamp 1621261055
transform 1 0 23904 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_245
timestamp 1621261055
transform 1 0 24672 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_253
timestamp 1621261055
transform 1 0 25440 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_261
timestamp 1621261055
transform 1 0 26208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_269
timestamp 1621261055
transform 1 0 26976 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_273
timestamp 1621261055
transform 1 0 27360 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_273
timestamp 1621261055
transform 1 0 27552 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_276
timestamp 1621261055
transform 1 0 27648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_284
timestamp 1621261055
transform 1 0 28416 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_292
timestamp 1621261055
transform 1 0 29184 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_300
timestamp 1621261055
transform 1 0 29952 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_308
timestamp 1621261055
transform 1 0 30720 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_274
timestamp 1621261055
transform 1 0 32832 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_316
timestamp 1621261055
transform 1 0 31488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_324
timestamp 1621261055
transform 1 0 32256 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_328
timestamp 1621261055
transform 1 0 32640 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_331
timestamp 1621261055
transform 1 0 32928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_339
timestamp 1621261055
transform 1 0 33696 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_347
timestamp 1621261055
transform 1 0 34464 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_355
timestamp 1621261055
transform 1 0 35232 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_363
timestamp 1621261055
transform 1 0 36000 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_371
timestamp 1621261055
transform 1 0 36768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _185_
timestamp 1621261055
transform 1 0 39360 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_275
timestamp 1621261055
transform 1 0 38112 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_379
timestamp 1621261055
transform 1 0 37536 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_383
timestamp 1621261055
transform 1 0 37920 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_386
timestamp 1621261055
transform 1 0 38208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_394
timestamp 1621261055
transform 1 0 38976 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_401
timestamp 1621261055
transform 1 0 39648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_409
timestamp 1621261055
transform 1 0 40416 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_417
timestamp 1621261055
transform 1 0 41184 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_276
timestamp 1621261055
transform 1 0 43392 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_425
timestamp 1621261055
transform 1 0 41952 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_433
timestamp 1621261055
transform 1 0 42720 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_437
timestamp 1621261055
transform 1 0 43104 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_439
timestamp 1621261055
transform 1 0 43296 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_441
timestamp 1621261055
transform 1 0 43488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_449
timestamp 1621261055
transform 1 0 44256 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_457
timestamp 1621261055
transform 1 0 45024 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_465
timestamp 1621261055
transform 1 0 45792 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_473
timestamp 1621261055
transform 1 0 46560 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_481
timestamp 1621261055
transform 1 0 47328 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_277
timestamp 1621261055
transform 1 0 48672 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_489
timestamp 1621261055
transform 1 0 48096 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_493
timestamp 1621261055
transform 1 0 48480 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_496
timestamp 1621261055
transform 1 0 48768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_504
timestamp 1621261055
transform 1 0 49536 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _113_
timestamp 1621261055
transform 1 0 50496 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _166_
timestamp 1621261055
transform 1 0 49728 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_9_509
timestamp 1621261055
transform 1 0 50016 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_513
timestamp 1621261055
transform 1 0 50400 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_517
timestamp 1621261055
transform 1 0 50784 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_525
timestamp 1621261055
transform 1 0 51552 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _067_
timestamp 1621261055
transform 1 0 51936 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output469
timestamp 1621261055
transform 1 0 53184 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_532
timestamp 1621261055
transform 1 0 52224 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_540
timestamp 1621261055
transform 1 0 52992 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_9_546
timestamp 1621261055
transform 1 0 53568 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_278
timestamp 1621261055
transform 1 0 53952 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output457
timestamp 1621261055
transform 1 0 54432 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output459
timestamp 1621261055
transform -1 0 55584 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_113
timestamp 1621261055
transform -1 0 55200 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_9_551
timestamp 1621261055
transform 1 0 54048 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_559
timestamp 1621261055
transform 1 0 54816 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_567
timestamp 1621261055
transform 1 0 55584 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input190
timestamp 1621261055
transform 1 0 57216 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input195
timestamp 1621261055
transform 1 0 56448 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_575
timestamp 1621261055
transform 1 0 56352 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_580
timestamp 1621261055
transform 1 0 56832 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_588
timestamp 1621261055
transform 1 0 57600 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_19
timestamp 1621261055
transform -1 0 58848 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_596
timestamp 1621261055
transform 1 0 58368 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_20
timestamp 1621261055
transform 1 0 1152 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_4
timestamp 1621261055
transform 1 0 1536 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_12
timestamp 1621261055
transform 1 0 2304 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_20
timestamp 1621261055
transform 1 0 3072 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_279
timestamp 1621261055
transform 1 0 3840 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_29
timestamp 1621261055
transform 1 0 3936 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_37
timestamp 1621261055
transform 1 0 4704 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_45
timestamp 1621261055
transform 1 0 5472 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_53
timestamp 1621261055
transform 1 0 6240 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_61
timestamp 1621261055
transform 1 0 7008 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_280
timestamp 1621261055
transform 1 0 9120 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_69
timestamp 1621261055
transform 1 0 7776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_77
timestamp 1621261055
transform 1 0 8544 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_81
timestamp 1621261055
transform 1 0 8928 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_84
timestamp 1621261055
transform 1 0 9216 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_92
timestamp 1621261055
transform 1 0 9984 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_100
timestamp 1621261055
transform 1 0 10752 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_108
timestamp 1621261055
transform 1 0 11520 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_116
timestamp 1621261055
transform 1 0 12288 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_124
timestamp 1621261055
transform 1 0 13056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_281
timestamp 1621261055
transform 1 0 14400 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_132
timestamp 1621261055
transform 1 0 13824 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_136
timestamp 1621261055
transform 1 0 14208 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_139
timestamp 1621261055
transform 1 0 14496 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_147
timestamp 1621261055
transform 1 0 15264 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_155
timestamp 1621261055
transform 1 0 16032 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_163
timestamp 1621261055
transform 1 0 16800 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_171
timestamp 1621261055
transform 1 0 17568 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_179
timestamp 1621261055
transform 1 0 18336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_187
timestamp 1621261055
transform 1 0 19104 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_282
timestamp 1621261055
transform 1 0 19680 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_191
timestamp 1621261055
transform 1 0 19488 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_194
timestamp 1621261055
transform 1 0 19776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_202
timestamp 1621261055
transform 1 0 20544 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_210
timestamp 1621261055
transform 1 0 21312 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_218
timestamp 1621261055
transform 1 0 22080 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_226
timestamp 1621261055
transform 1 0 22848 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _059_
timestamp 1621261055
transform 1 0 24288 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_283
timestamp 1621261055
transform 1 0 24960 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_80
timestamp 1621261055
transform 1 0 24096 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_10_234
timestamp 1621261055
transform 1 0 23616 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_238
timestamp 1621261055
transform 1 0 24000 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_244
timestamp 1621261055
transform 1 0 24576 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_249
timestamp 1621261055
transform 1 0 25056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_257
timestamp 1621261055
transform 1 0 25824 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_265
timestamp 1621261055
transform 1 0 26592 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_273
timestamp 1621261055
transform 1 0 27360 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_281
timestamp 1621261055
transform 1 0 28128 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_289
timestamp 1621261055
transform 1 0 28896 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_284
timestamp 1621261055
transform 1 0 30240 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_297
timestamp 1621261055
transform 1 0 29664 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_301
timestamp 1621261055
transform 1 0 30048 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_304
timestamp 1621261055
transform 1 0 30336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_312
timestamp 1621261055
transform 1 0 31104 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_320
timestamp 1621261055
transform 1 0 31872 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_328
timestamp 1621261055
transform 1 0 32640 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_336
timestamp 1621261055
transform 1 0 33408 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_344
timestamp 1621261055
transform 1 0 34176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_352
timestamp 1621261055
transform 1 0 34944 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_356
timestamp 1621261055
transform 1 0 35328 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_285
timestamp 1621261055
transform 1 0 35520 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_359
timestamp 1621261055
transform 1 0 35616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_367
timestamp 1621261055
transform 1 0 36384 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_375
timestamp 1621261055
transform 1 0 37152 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_383
timestamp 1621261055
transform 1 0 37920 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_391
timestamp 1621261055
transform 1 0 38688 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_399
timestamp 1621261055
transform 1 0 39456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_286
timestamp 1621261055
transform 1 0 40800 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_407
timestamp 1621261055
transform 1 0 40224 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_411
timestamp 1621261055
transform 1 0 40608 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_414
timestamp 1621261055
transform 1 0 40896 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_422
timestamp 1621261055
transform 1 0 41664 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_430
timestamp 1621261055
transform 1 0 42432 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_438
timestamp 1621261055
transform 1 0 43200 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_446
timestamp 1621261055
transform 1 0 43968 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_454
timestamp 1621261055
transform 1 0 44736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_462
timestamp 1621261055
transform 1 0 45504 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_287
timestamp 1621261055
transform 1 0 46080 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_466
timestamp 1621261055
transform 1 0 45888 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_469
timestamp 1621261055
transform 1 0 46176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_477
timestamp 1621261055
transform 1 0 46944 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_485
timestamp 1621261055
transform 1 0 47712 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_493
timestamp 1621261055
transform 1 0 48480 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_501
timestamp 1621261055
transform 1 0 49248 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _122_
timestamp 1621261055
transform 1 0 50112 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_288
timestamp 1621261055
transform 1 0 51360 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_10_509
timestamp 1621261055
transform 1 0 50016 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_513
timestamp 1621261055
transform 1 0 50400 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_521
timestamp 1621261055
transform 1 0 51168 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_524
timestamp 1621261055
transform 1 0 51456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _075_
timestamp 1621261055
transform 1 0 52416 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_532
timestamp 1621261055
transform 1 0 52224 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_537
timestamp 1621261055
transform 1 0 52704 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_545
timestamp 1621261055
transform 1 0 53472 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output458
timestamp 1621261055
transform 1 0 54240 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output460
timestamp 1621261055
transform -1 0 55392 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_114
timestamp 1621261055
transform -1 0 55008 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_116
timestamp 1621261055
transform -1 0 55776 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_557
timestamp 1621261055
transform 1 0 54624 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_565
timestamp 1621261055
transform 1 0 55392 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_289
timestamp 1621261055
transform 1 0 56640 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input191
timestamp 1621261055
transform 1 0 57600 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output461
timestamp 1621261055
transform -1 0 56160 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_117
timestamp 1621261055
transform -1 0 56352 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_575
timestamp 1621261055
transform 1 0 56352 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_577
timestamp 1621261055
transform 1 0 56544 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_579
timestamp 1621261055
transform 1 0 56736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_10_587
timestamp 1621261055
transform 1 0 57504 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_21
timestamp 1621261055
transform -1 0 58848 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_592
timestamp 1621261055
transform 1 0 57984 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_596
timestamp 1621261055
transform 1 0 58368 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_22
timestamp 1621261055
transform 1 0 1152 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_4
timestamp 1621261055
transform 1 0 1536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_12
timestamp 1621261055
transform 1 0 2304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_20
timestamp 1621261055
transform 1 0 3072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_28
timestamp 1621261055
transform 1 0 3840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_36
timestamp 1621261055
transform 1 0 4608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_290
timestamp 1621261055
transform 1 0 6432 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_44
timestamp 1621261055
transform 1 0 5376 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_52
timestamp 1621261055
transform 1 0 6144 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_54
timestamp 1621261055
transform 1 0 6336 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_56
timestamp 1621261055
transform 1 0 6528 0 1 9990
box -38 -49 806 715
use BUFX2  BUFX2
timestamp 1624074425
transform 1 0 7680 0 1 9990
box 0 -48 864 714
use sky130_fd_sc_ls__diode_2  ANTENNA_47
timestamp 1621261055
transform 1 0 7488 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_64
timestamp 1621261055
transform 1 0 7296 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_77
timestamp 1621261055
transform 1 0 8544 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_85
timestamp 1621261055
transform 1 0 9312 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_93
timestamp 1621261055
transform 1 0 10080 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_101
timestamp 1621261055
transform 1 0 10848 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_291
timestamp 1621261055
transform 1 0 11712 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_11_109
timestamp 1621261055
transform 1 0 11616 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_111
timestamp 1621261055
transform 1 0 11808 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_119
timestamp 1621261055
transform 1 0 12576 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_127
timestamp 1621261055
transform 1 0 13344 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_135
timestamp 1621261055
transform 1 0 14112 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_143
timestamp 1621261055
transform 1 0 14880 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_292
timestamp 1621261055
transform 1 0 16992 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_151
timestamp 1621261055
transform 1 0 15648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_159
timestamp 1621261055
transform 1 0 16416 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_163
timestamp 1621261055
transform 1 0 16800 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_166
timestamp 1621261055
transform 1 0 17088 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_174
timestamp 1621261055
transform 1 0 17856 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_182
timestamp 1621261055
transform 1 0 18624 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_190
timestamp 1621261055
transform 1 0 19392 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_198
timestamp 1621261055
transform 1 0 20160 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_206
timestamp 1621261055
transform 1 0 20928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_293
timestamp 1621261055
transform 1 0 22272 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_214
timestamp 1621261055
transform 1 0 21696 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_218
timestamp 1621261055
transform 1 0 22080 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_221
timestamp 1621261055
transform 1 0 22368 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_229
timestamp 1621261055
transform 1 0 23136 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_237
timestamp 1621261055
transform 1 0 23904 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_245
timestamp 1621261055
transform 1 0 24672 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_253
timestamp 1621261055
transform 1 0 25440 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_261
timestamp 1621261055
transform 1 0 26208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_269
timestamp 1621261055
transform 1 0 26976 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_273
timestamp 1621261055
transform 1 0 27360 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_294
timestamp 1621261055
transform 1 0 27552 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_276
timestamp 1621261055
transform 1 0 27648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_284
timestamp 1621261055
transform 1 0 28416 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_292
timestamp 1621261055
transform 1 0 29184 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_300
timestamp 1621261055
transform 1 0 29952 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_308
timestamp 1621261055
transform 1 0 30720 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_295
timestamp 1621261055
transform 1 0 32832 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_316
timestamp 1621261055
transform 1 0 31488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_324
timestamp 1621261055
transform 1 0 32256 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_328
timestamp 1621261055
transform 1 0 32640 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_331
timestamp 1621261055
transform 1 0 32928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_339
timestamp 1621261055
transform 1 0 33696 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_347
timestamp 1621261055
transform 1 0 34464 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_355
timestamp 1621261055
transform 1 0 35232 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_363
timestamp 1621261055
transform 1 0 36000 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_371
timestamp 1621261055
transform 1 0 36768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _160_
timestamp 1621261055
transform 1 0 39360 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_296
timestamp 1621261055
transform 1 0 38112 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_379
timestamp 1621261055
transform 1 0 37536 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_383
timestamp 1621261055
transform 1 0 37920 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_386
timestamp 1621261055
transform 1 0 38208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_394
timestamp 1621261055
transform 1 0 38976 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_401
timestamp 1621261055
transform 1 0 39648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_409
timestamp 1621261055
transform 1 0 40416 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_417
timestamp 1621261055
transform 1 0 41184 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_297
timestamp 1621261055
transform 1 0 43392 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_425
timestamp 1621261055
transform 1 0 41952 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_433
timestamp 1621261055
transform 1 0 42720 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_437
timestamp 1621261055
transform 1 0 43104 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_439
timestamp 1621261055
transform 1 0 43296 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_441
timestamp 1621261055
transform 1 0 43488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_449
timestamp 1621261055
transform 1 0 44256 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_457
timestamp 1621261055
transform 1 0 45024 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_465
timestamp 1621261055
transform 1 0 45792 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_473
timestamp 1621261055
transform 1 0 46560 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_481
timestamp 1621261055
transform 1 0 47328 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_298
timestamp 1621261055
transform 1 0 48672 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_489
timestamp 1621261055
transform 1 0 48096 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_493
timestamp 1621261055
transform 1 0 48480 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_496
timestamp 1621261055
transform 1 0 48768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_504
timestamp 1621261055
transform 1 0 49536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_512
timestamp 1621261055
transform 1 0 50304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_520
timestamp 1621261055
transform 1 0 51072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_528
timestamp 1621261055
transform 1 0 51840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_536
timestamp 1621261055
transform 1 0 52608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_544
timestamp 1621261055
transform 1 0 53376 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_299
timestamp 1621261055
transform 1 0 53952 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output471
timestamp 1621261055
transform -1 0 55296 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_125
timestamp 1621261055
transform -1 0 54912 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_548
timestamp 1621261055
transform 1 0 53760 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_551
timestamp 1621261055
transform 1 0 54048 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_555
timestamp 1621261055
transform 1 0 54432 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_557
timestamp 1621261055
transform 1 0 54624 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_564
timestamp 1621261055
transform 1 0 55296 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output462
timestamp 1621261055
transform 1 0 55680 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output463
timestamp 1621261055
transform 1 0 56448 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output464
timestamp 1621261055
transform 1 0 57216 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_119
timestamp 1621261055
transform 1 0 56256 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_572
timestamp 1621261055
transform 1 0 56064 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_580
timestamp 1621261055
transform 1 0 56832 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_588
timestamp 1621261055
transform 1 0 57600 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_23
timestamp 1621261055
transform -1 0 58848 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_596
timestamp 1621261055
transform 1 0 58368 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_24
timestamp 1621261055
transform 1 0 1152 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_12_4
timestamp 1621261055
transform 1 0 1536 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_12
timestamp 1621261055
transform 1 0 2304 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_20
timestamp 1621261055
transform 1 0 3072 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_300
timestamp 1621261055
transform 1 0 3840 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_29
timestamp 1621261055
transform 1 0 3936 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_37
timestamp 1621261055
transform 1 0 4704 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_45
timestamp 1621261055
transform 1 0 5472 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_53
timestamp 1621261055
transform 1 0 6240 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_61
timestamp 1621261055
transform 1 0 7008 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _153_
timestamp 1621261055
transform 1 0 7872 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_301
timestamp 1621261055
transform 1 0 9120 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_12_69
timestamp 1621261055
transform 1 0 7776 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_73
timestamp 1621261055
transform 1 0 8160 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_81
timestamp 1621261055
transform 1 0 8928 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_12_84
timestamp 1621261055
transform 1 0 9216 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _064_
timestamp 1621261055
transform 1 0 9696 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_12_88
timestamp 1621261055
transform 1 0 9600 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_92
timestamp 1621261055
transform 1 0 9984 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_100
timestamp 1621261055
transform 1 0 10752 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_108
timestamp 1621261055
transform 1 0 11520 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_116
timestamp 1621261055
transform 1 0 12288 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_124
timestamp 1621261055
transform 1 0 13056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_302
timestamp 1621261055
transform 1 0 14400 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_132
timestamp 1621261055
transform 1 0 13824 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_136
timestamp 1621261055
transform 1 0 14208 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_139
timestamp 1621261055
transform 1 0 14496 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_147
timestamp 1621261055
transform 1 0 15264 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_155
timestamp 1621261055
transform 1 0 16032 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_163
timestamp 1621261055
transform 1 0 16800 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _215_
timestamp 1621261055
transform -1 0 19296 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_16
timestamp 1621261055
transform -1 0 19008 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_171
timestamp 1621261055
transform 1 0 17568 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_179
timestamp 1621261055
transform 1 0 18336 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_12_183
timestamp 1621261055
transform 1 0 18720 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_189
timestamp 1621261055
transform 1 0 19296 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_303
timestamp 1621261055
transform 1 0 19680 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_194
timestamp 1621261055
transform 1 0 19776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_202
timestamp 1621261055
transform 1 0 20544 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_210
timestamp 1621261055
transform 1 0 21312 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_218
timestamp 1621261055
transform 1 0 22080 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_226
timestamp 1621261055
transform 1 0 22848 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_304
timestamp 1621261055
transform 1 0 24960 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_234
timestamp 1621261055
transform 1 0 23616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_242
timestamp 1621261055
transform 1 0 24384 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_246
timestamp 1621261055
transform 1 0 24768 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_249
timestamp 1621261055
transform 1 0 25056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_257
timestamp 1621261055
transform 1 0 25824 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_265
timestamp 1621261055
transform 1 0 26592 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_273
timestamp 1621261055
transform 1 0 27360 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _107_
timestamp 1621261055
transform 1 0 29184 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_281
timestamp 1621261055
transform 1 0 28128 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_289
timestamp 1621261055
transform 1 0 28896 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_291
timestamp 1621261055
transform 1 0 29088 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_305
timestamp 1621261055
transform 1 0 30240 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_295
timestamp 1621261055
transform 1 0 29472 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_304
timestamp 1621261055
transform 1 0 30336 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_312
timestamp 1621261055
transform 1 0 31104 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _080_
timestamp 1621261055
transform 1 0 32256 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_12_320
timestamp 1621261055
transform 1 0 31872 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_12_327
timestamp 1621261055
transform 1 0 32544 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_335
timestamp 1621261055
transform 1 0 33312 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_343
timestamp 1621261055
transform 1 0 34080 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_351
timestamp 1621261055
transform 1 0 34848 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_355
timestamp 1621261055
transform 1 0 35232 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_357
timestamp 1621261055
transform 1 0 35424 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_306
timestamp 1621261055
transform 1 0 35520 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_359
timestamp 1621261055
transform 1 0 35616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_367
timestamp 1621261055
transform 1 0 36384 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_375
timestamp 1621261055
transform 1 0 37152 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_383
timestamp 1621261055
transform 1 0 37920 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_391
timestamp 1621261055
transform 1 0 38688 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_399
timestamp 1621261055
transform 1 0 39456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_307
timestamp 1621261055
transform 1 0 40800 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_407
timestamp 1621261055
transform 1 0 40224 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_411
timestamp 1621261055
transform 1 0 40608 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_414
timestamp 1621261055
transform 1 0 40896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_422
timestamp 1621261055
transform 1 0 41664 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_430
timestamp 1621261055
transform 1 0 42432 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_438
timestamp 1621261055
transform 1 0 43200 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_446
timestamp 1621261055
transform 1 0 43968 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_454
timestamp 1621261055
transform 1 0 44736 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_462
timestamp 1621261055
transform 1 0 45504 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_308
timestamp 1621261055
transform 1 0 46080 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_466
timestamp 1621261055
transform 1 0 45888 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_469
timestamp 1621261055
transform 1 0 46176 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_477
timestamp 1621261055
transform 1 0 46944 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _047_
timestamp 1621261055
transform -1 0 49056 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_49
timestamp 1621261055
transform -1 0 48768 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_485
timestamp 1621261055
transform 1 0 47712 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_12_493
timestamp 1621261055
transform 1 0 48480 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_499
timestamp 1621261055
transform 1 0 49056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_309
timestamp 1621261055
transform 1 0 51360 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_507
timestamp 1621261055
transform 1 0 49824 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_515
timestamp 1621261055
transform 1 0 50592 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_524
timestamp 1621261055
transform 1 0 51456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_532
timestamp 1621261055
transform 1 0 52224 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_540
timestamp 1621261055
transform 1 0 52992 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _110_
timestamp 1621261055
transform 1 0 54432 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_12_548
timestamp 1621261055
transform 1 0 53760 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_552
timestamp 1621261055
transform 1 0 54144 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_554
timestamp 1621261055
transform 1 0 54336 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_558
timestamp 1621261055
transform 1 0 54720 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_566
timestamp 1621261055
transform 1 0 55488 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_310
timestamp 1621261055
transform 1 0 56640 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output465
timestamp 1621261055
transform -1 0 57504 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output470
timestamp 1621261055
transform 1 0 55872 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_120
timestamp 1621261055
transform -1 0 57120 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_12_574
timestamp 1621261055
transform 1 0 56256 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_579
timestamp 1621261055
transform 1 0 56736 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_587
timestamp 1621261055
transform 1 0 57504 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_25
timestamp 1621261055
transform -1 0 58848 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_595
timestamp 1621261055
transform 1 0 58272 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_26
timestamp 1621261055
transform 1 0 1152 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_4
timestamp 1621261055
transform 1 0 1536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_12
timestamp 1621261055
transform 1 0 2304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_20
timestamp 1621261055
transform 1 0 3072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_28
timestamp 1621261055
transform 1 0 3840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_36
timestamp 1621261055
transform 1 0 4608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_311
timestamp 1621261055
transform 1 0 6432 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_44
timestamp 1621261055
transform 1 0 5376 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_52
timestamp 1621261055
transform 1 0 6144 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_54
timestamp 1621261055
transform 1 0 6336 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_56
timestamp 1621261055
transform 1 0 6528 0 1 11322
box -38 -49 806 715
use INV  INV
timestamp 1624074425
transform 1 0 7680 0 1 11322
box 0 -48 576 714
use sky130_fd_sc_ls__diode_2  ANTENNA_51
timestamp 1621261055
transform 1 0 7488 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_64
timestamp 1621261055
transform 1 0 7296 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_74
timestamp 1621261055
transform 1 0 8256 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_82
timestamp 1621261055
transform 1 0 9024 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_90
timestamp 1621261055
transform 1 0 9792 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_98
timestamp 1621261055
transform 1 0 10560 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_312
timestamp 1621261055
transform 1 0 11712 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_106
timestamp 1621261055
transform 1 0 11328 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_111
timestamp 1621261055
transform 1 0 11808 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_119
timestamp 1621261055
transform 1 0 12576 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_127
timestamp 1621261055
transform 1 0 13344 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_135
timestamp 1621261055
transform 1 0 14112 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_143
timestamp 1621261055
transform 1 0 14880 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_313
timestamp 1621261055
transform 1 0 16992 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_151
timestamp 1621261055
transform 1 0 15648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_159
timestamp 1621261055
transform 1 0 16416 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_163
timestamp 1621261055
transform 1 0 16800 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_166
timestamp 1621261055
transform 1 0 17088 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_174
timestamp 1621261055
transform 1 0 17856 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_182
timestamp 1621261055
transform 1 0 18624 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_190
timestamp 1621261055
transform 1 0 19392 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_198
timestamp 1621261055
transform 1 0 20160 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_206
timestamp 1621261055
transform 1 0 20928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_314
timestamp 1621261055
transform 1 0 22272 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_214
timestamp 1621261055
transform 1 0 21696 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_218
timestamp 1621261055
transform 1 0 22080 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_221
timestamp 1621261055
transform 1 0 22368 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_229
timestamp 1621261055
transform 1 0 23136 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _126_
timestamp 1621261055
transform 1 0 23712 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_233
timestamp 1621261055
transform 1 0 23520 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_238
timestamp 1621261055
transform 1 0 24000 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_246
timestamp 1621261055
transform 1 0 24768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_254
timestamp 1621261055
transform 1 0 25536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_262
timestamp 1621261055
transform 1 0 26304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_270
timestamp 1621261055
transform 1 0 27072 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_315
timestamp 1621261055
transform 1 0 27552 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_13_274
timestamp 1621261055
transform 1 0 27456 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_276
timestamp 1621261055
transform 1 0 27648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_284
timestamp 1621261055
transform 1 0 28416 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_292
timestamp 1621261055
transform 1 0 29184 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_300
timestamp 1621261055
transform 1 0 29952 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_308
timestamp 1621261055
transform 1 0 30720 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_316
timestamp 1621261055
transform 1 0 32832 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_316
timestamp 1621261055
transform 1 0 31488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_324
timestamp 1621261055
transform 1 0 32256 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_328
timestamp 1621261055
transform 1 0 32640 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_331
timestamp 1621261055
transform 1 0 32928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_339
timestamp 1621261055
transform 1 0 33696 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_347
timestamp 1621261055
transform 1 0 34464 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_355
timestamp 1621261055
transform 1 0 35232 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_363
timestamp 1621261055
transform 1 0 36000 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_371
timestamp 1621261055
transform 1 0 36768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_317
timestamp 1621261055
transform 1 0 38112 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_379
timestamp 1621261055
transform 1 0 37536 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_383
timestamp 1621261055
transform 1 0 37920 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_386
timestamp 1621261055
transform 1 0 38208 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_394
timestamp 1621261055
transform 1 0 38976 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_402
timestamp 1621261055
transform 1 0 39744 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_410
timestamp 1621261055
transform 1 0 40512 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_418
timestamp 1621261055
transform 1 0 41280 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_318
timestamp 1621261055
transform 1 0 43392 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_426
timestamp 1621261055
transform 1 0 42048 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_434
timestamp 1621261055
transform 1 0 42816 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_438
timestamp 1621261055
transform 1 0 43200 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_441
timestamp 1621261055
transform 1 0 43488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_449
timestamp 1621261055
transform 1 0 44256 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_457
timestamp 1621261055
transform 1 0 45024 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_465
timestamp 1621261055
transform 1 0 45792 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_473
timestamp 1621261055
transform 1 0 46560 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_481
timestamp 1621261055
transform 1 0 47328 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_319
timestamp 1621261055
transform 1 0 48672 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_489
timestamp 1621261055
transform 1 0 48096 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_493
timestamp 1621261055
transform 1 0 48480 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_496
timestamp 1621261055
transform 1 0 48768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_504
timestamp 1621261055
transform 1 0 49536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_512
timestamp 1621261055
transform 1 0 50304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_520
timestamp 1621261055
transform 1 0 51072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_528
timestamp 1621261055
transform 1 0 51840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_536
timestamp 1621261055
transform 1 0 52608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_544
timestamp 1621261055
transform 1 0 53376 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_320
timestamp 1621261055
transform 1 0 53952 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_548
timestamp 1621261055
transform 1 0 53760 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_551
timestamp 1621261055
transform 1 0 54048 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_559
timestamp 1621261055
transform 1 0 54816 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_13_567
timestamp 1621261055
transform 1 0 55584 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _207_
timestamp 1621261055
transform 1 0 55680 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output467
timestamp 1621261055
transform -1 0 57504 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output474
timestamp 1621261055
transform -1 0 56736 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_121
timestamp 1621261055
transform -1 0 57120 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_127
timestamp 1621261055
transform -1 0 56352 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_571
timestamp 1621261055
transform 1 0 55968 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_579
timestamp 1621261055
transform 1 0 56736 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_587
timestamp 1621261055
transform 1 0 57504 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_27
timestamp 1621261055
transform -1 0 58848 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_595
timestamp 1621261055
transform 1 0 58272 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _208_
timestamp 1621261055
transform 1 0 1920 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_28
timestamp 1621261055
transform 1 0 1152 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_14_4
timestamp 1621261055
transform 1 0 1536 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_14_11
timestamp 1621261055
transform 1 0 2208 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_19
timestamp 1621261055
transform 1 0 2976 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_321
timestamp 1621261055
transform 1 0 3840 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_14_27
timestamp 1621261055
transform 1 0 3744 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_29
timestamp 1621261055
transform 1 0 3936 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_37
timestamp 1621261055
transform 1 0 4704 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _164_
timestamp 1621261055
transform 1 0 6336 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_14_45
timestamp 1621261055
transform 1 0 5472 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_14_53
timestamp 1621261055
transform 1 0 6240 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_57
timestamp 1621261055
transform 1 0 6624 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_322
timestamp 1621261055
transform 1 0 9120 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_65
timestamp 1621261055
transform 1 0 7392 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_73
timestamp 1621261055
transform 1 0 8160 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_81
timestamp 1621261055
transform 1 0 8928 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_84
timestamp 1621261055
transform 1 0 9216 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_92
timestamp 1621261055
transform 1 0 9984 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_100
timestamp 1621261055
transform 1 0 10752 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_108
timestamp 1621261055
transform 1 0 11520 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_116
timestamp 1621261055
transform 1 0 12288 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_124
timestamp 1621261055
transform 1 0 13056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_323
timestamp 1621261055
transform 1 0 14400 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_132
timestamp 1621261055
transform 1 0 13824 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_136
timestamp 1621261055
transform 1 0 14208 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_139
timestamp 1621261055
transform 1 0 14496 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_147
timestamp 1621261055
transform 1 0 15264 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_155
timestamp 1621261055
transform 1 0 16032 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_163
timestamp 1621261055
transform 1 0 16800 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_171
timestamp 1621261055
transform 1 0 17568 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_179
timestamp 1621261055
transform 1 0 18336 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_187
timestamp 1621261055
transform 1 0 19104 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_324
timestamp 1621261055
transform 1 0 19680 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_191
timestamp 1621261055
transform 1 0 19488 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_194
timestamp 1621261055
transform 1 0 19776 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_202
timestamp 1621261055
transform 1 0 20544 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_210
timestamp 1621261055
transform 1 0 21312 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_218
timestamp 1621261055
transform 1 0 22080 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_226
timestamp 1621261055
transform 1 0 22848 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_325
timestamp 1621261055
transform 1 0 24960 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_234
timestamp 1621261055
transform 1 0 23616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_242
timestamp 1621261055
transform 1 0 24384 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_246
timestamp 1621261055
transform 1 0 24768 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_249
timestamp 1621261055
transform 1 0 25056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_257
timestamp 1621261055
transform 1 0 25824 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_265
timestamp 1621261055
transform 1 0 26592 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_273
timestamp 1621261055
transform 1 0 27360 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_281
timestamp 1621261055
transform 1 0 28128 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_289
timestamp 1621261055
transform 1 0 28896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_326
timestamp 1621261055
transform 1 0 30240 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_297
timestamp 1621261055
transform 1 0 29664 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_301
timestamp 1621261055
transform 1 0 30048 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_304
timestamp 1621261055
transform 1 0 30336 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_312
timestamp 1621261055
transform 1 0 31104 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_320
timestamp 1621261055
transform 1 0 31872 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_328
timestamp 1621261055
transform 1 0 32640 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_336
timestamp 1621261055
transform 1 0 33408 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_344
timestamp 1621261055
transform 1 0 34176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_352
timestamp 1621261055
transform 1 0 34944 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_356
timestamp 1621261055
transform 1 0 35328 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_327
timestamp 1621261055
transform 1 0 35520 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_25
timestamp 1621261055
transform -1 0 37536 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_359
timestamp 1621261055
transform 1 0 35616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_367
timestamp 1621261055
transform 1 0 36384 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_375
timestamp 1621261055
transform 1 0 37152 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _015_
timestamp 1621261055
transform -1 0 37824 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_14_382
timestamp 1621261055
transform 1 0 37824 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_390
timestamp 1621261055
transform 1 0 38592 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_398
timestamp 1621261055
transform 1 0 39360 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_328
timestamp 1621261055
transform 1 0 40800 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_406
timestamp 1621261055
transform 1 0 40128 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_410
timestamp 1621261055
transform 1 0 40512 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_14_412
timestamp 1621261055
transform 1 0 40704 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_414
timestamp 1621261055
transform 1 0 40896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_422
timestamp 1621261055
transform 1 0 41664 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_430
timestamp 1621261055
transform 1 0 42432 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_438
timestamp 1621261055
transform 1 0 43200 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_446
timestamp 1621261055
transform 1 0 43968 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_454
timestamp 1621261055
transform 1 0 44736 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_462
timestamp 1621261055
transform 1 0 45504 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_329
timestamp 1621261055
transform 1 0 46080 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_466
timestamp 1621261055
transform 1 0 45888 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_469
timestamp 1621261055
transform 1 0 46176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_477
timestamp 1621261055
transform 1 0 46944 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _041_
timestamp 1621261055
transform -1 0 49440 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_91
timestamp 1621261055
transform -1 0 49152 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_485
timestamp 1621261055
transform 1 0 47712 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_493
timestamp 1621261055
transform 1 0 48480 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_14_497
timestamp 1621261055
transform 1 0 48864 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_503
timestamp 1621261055
transform 1 0 49440 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_330
timestamp 1621261055
transform 1 0 51360 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_511
timestamp 1621261055
transform 1 0 50208 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_519
timestamp 1621261055
transform 1 0 50976 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_14_524
timestamp 1621261055
transform 1 0 51456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_532
timestamp 1621261055
transform 1 0 52224 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_540
timestamp 1621261055
transform 1 0 52992 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_548
timestamp 1621261055
transform 1 0 53760 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_556
timestamp 1621261055
transform 1 0 54528 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_564
timestamp 1621261055
transform 1 0 55296 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_331
timestamp 1621261055
transform 1 0 56640 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output468
timestamp 1621261055
transform -1 0 57888 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_123
timestamp 1621261055
transform -1 0 57504 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_572
timestamp 1621261055
transform 1 0 56064 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_576
timestamp 1621261055
transform 1 0 56448 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_579
timestamp 1621261055
transform 1 0 56736 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_583
timestamp 1621261055
transform 1 0 57120 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_29
timestamp 1621261055
transform -1 0 58848 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_124
timestamp 1621261055
transform -1 0 58080 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_593
timestamp 1621261055
transform 1 0 58080 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_30
timestamp 1621261055
transform 1 0 1152 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_32
timestamp 1621261055
transform 1 0 1152 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_4
timestamp 1621261055
transform 1 0 1536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_12
timestamp 1621261055
transform 1 0 2304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_20
timestamp 1621261055
transform 1 0 3072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_4
timestamp 1621261055
transform 1 0 1536 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_12
timestamp 1621261055
transform 1 0 2304 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_20
timestamp 1621261055
transform 1 0 3072 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_342
timestamp 1621261055
transform 1 0 3840 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_28
timestamp 1621261055
transform 1 0 3840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_36
timestamp 1621261055
transform 1 0 4608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_29
timestamp 1621261055
transform 1 0 3936 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_37
timestamp 1621261055
transform 1 0 4704 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_332
timestamp 1621261055
transform 1 0 6432 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_44
timestamp 1621261055
transform 1 0 5376 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_52
timestamp 1621261055
transform 1 0 6144 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_15_54
timestamp 1621261055
transform 1 0 6336 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_56
timestamp 1621261055
transform 1 0 6528 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_45
timestamp 1621261055
transform 1 0 5472 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_53
timestamp 1621261055
transform 1 0 6240 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_61
timestamp 1621261055
transform 1 0 7008 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_69
timestamp 1621261055
transform 1 0 7776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_64
timestamp 1621261055
transform 1 0 7296 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_57
timestamp 1621261055
transform 1 0 7488 0 1 12654
box -38 -49 230 715
use INVX1  INVX1
timestamp 1624074425
transform 1 0 7680 0 1 12654
box 0 -48 576 714
use sky130_fd_sc_ls__decap_4  FILLER_16_77
timestamp 1621261055
transform 1 0 8544 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_74
timestamp 1621261055
transform 1 0 8256 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_84
timestamp 1621261055
transform 1 0 9216 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_81
timestamp 1621261055
transform 1 0 8928 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_82
timestamp 1621261055
transform 1 0 9024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_343
timestamp 1621261055
transform 1 0 9120 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _179_
timestamp 1621261055
transform 1 0 11232 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_15_90
timestamp 1621261055
transform 1 0 9792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_98
timestamp 1621261055
transform 1 0 10560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_92
timestamp 1621261055
transform 1 0 9984 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_100
timestamp 1621261055
transform 1 0 10752 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_16_104
timestamp 1621261055
transform 1 0 11136 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_333
timestamp 1621261055
transform 1 0 11712 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_106
timestamp 1621261055
transform 1 0 11328 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_111
timestamp 1621261055
transform 1 0 11808 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_119
timestamp 1621261055
transform 1 0 12576 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_108
timestamp 1621261055
transform 1 0 11520 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_116
timestamp 1621261055
transform 1 0 12288 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_124
timestamp 1621261055
transform 1 0 13056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_344
timestamp 1621261055
transform 1 0 14400 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_127
timestamp 1621261055
transform 1 0 13344 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_135
timestamp 1621261055
transform 1 0 14112 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_143
timestamp 1621261055
transform 1 0 14880 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_132
timestamp 1621261055
transform 1 0 13824 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_136
timestamp 1621261055
transform 1 0 14208 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_139
timestamp 1621261055
transform 1 0 14496 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_147
timestamp 1621261055
transform 1 0 15264 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_151
timestamp 1621261055
transform 1 0 15648 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_151
timestamp 1621261055
transform 1 0 15648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_39
timestamp 1621261055
transform 1 0 15840 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _042_
timestamp 1621261055
transform 1 0 16032 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_158
timestamp 1621261055
transform 1 0 16320 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_163
timestamp 1621261055
transform 1 0 16800 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_159
timestamp 1621261055
transform 1 0 16416 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_166
timestamp 1621261055
transform 1 0 17088 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_166
timestamp 1621261055
transform 1 0 17088 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_334
timestamp 1621261055
transform 1 0 16992 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_174
timestamp 1621261055
transform 1 0 17856 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_182
timestamp 1621261055
transform 1 0 18624 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_174
timestamp 1621261055
transform 1 0 17856 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_182
timestamp 1621261055
transform 1 0 18624 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_345
timestamp 1621261055
transform 1 0 19680 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_190
timestamp 1621261055
transform 1 0 19392 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_198
timestamp 1621261055
transform 1 0 20160 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_206
timestamp 1621261055
transform 1 0 20928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_190
timestamp 1621261055
transform 1 0 19392 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_16_192
timestamp 1621261055
transform 1 0 19584 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_194
timestamp 1621261055
transform 1 0 19776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_202
timestamp 1621261055
transform 1 0 20544 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_210
timestamp 1621261055
transform 1 0 21312 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_335
timestamp 1621261055
transform 1 0 22272 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_214
timestamp 1621261055
transform 1 0 21696 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_218
timestamp 1621261055
transform 1 0 22080 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_221
timestamp 1621261055
transform 1 0 22368 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_229
timestamp 1621261055
transform 1 0 23136 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_218
timestamp 1621261055
transform 1 0 22080 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_226
timestamp 1621261055
transform 1 0 22848 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_346
timestamp 1621261055
transform 1 0 24960 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_237
timestamp 1621261055
transform 1 0 23904 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_245
timestamp 1621261055
transform 1 0 24672 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_234
timestamp 1621261055
transform 1 0 23616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_242
timestamp 1621261055
transform 1 0 24384 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_246
timestamp 1621261055
transform 1 0 24768 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_249
timestamp 1621261055
transform 1 0 25056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_253
timestamp 1621261055
transform 1 0 25440 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_261
timestamp 1621261055
transform 1 0 26208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_269
timestamp 1621261055
transform 1 0 26976 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_273
timestamp 1621261055
transform 1 0 27360 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_257
timestamp 1621261055
transform 1 0 25824 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_265
timestamp 1621261055
transform 1 0 26592 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_273
timestamp 1621261055
transform 1 0 27360 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_336
timestamp 1621261055
transform 1 0 27552 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_276
timestamp 1621261055
transform 1 0 27648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_284
timestamp 1621261055
transform 1 0 28416 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_292
timestamp 1621261055
transform 1 0 29184 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_281
timestamp 1621261055
transform 1 0 28128 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_289
timestamp 1621261055
transform 1 0 28896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_347
timestamp 1621261055
transform 1 0 30240 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_300
timestamp 1621261055
transform 1 0 29952 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_308
timestamp 1621261055
transform 1 0 30720 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_297
timestamp 1621261055
transform 1 0 29664 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_301
timestamp 1621261055
transform 1 0 30048 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_304
timestamp 1621261055
transform 1 0 30336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_312
timestamp 1621261055
transform 1 0 31104 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_337
timestamp 1621261055
transform 1 0 32832 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_316
timestamp 1621261055
transform 1 0 31488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_324
timestamp 1621261055
transform 1 0 32256 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_328
timestamp 1621261055
transform 1 0 32640 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_331
timestamp 1621261055
transform 1 0 32928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_320
timestamp 1621261055
transform 1 0 31872 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_328
timestamp 1621261055
transform 1 0 32640 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_336
timestamp 1621261055
transform 1 0 33408 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_339
timestamp 1621261055
transform 1 0 33696 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_347
timestamp 1621261055
transform 1 0 34464 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_355
timestamp 1621261055
transform 1 0 35232 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_344
timestamp 1621261055
transform 1 0 34176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_352
timestamp 1621261055
transform 1 0 34944 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_356
timestamp 1621261055
transform 1 0 35328 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_348
timestamp 1621261055
transform 1 0 35520 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_363
timestamp 1621261055
transform 1 0 36000 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_371
timestamp 1621261055
transform 1 0 36768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_359
timestamp 1621261055
transform 1 0 35616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_367
timestamp 1621261055
transform 1 0 36384 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_375
timestamp 1621261055
transform 1 0 37152 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_338
timestamp 1621261055
transform 1 0 38112 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_379
timestamp 1621261055
transform 1 0 37536 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_383
timestamp 1621261055
transform 1 0 37920 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_386
timestamp 1621261055
transform 1 0 38208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_394
timestamp 1621261055
transform 1 0 38976 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_383
timestamp 1621261055
transform 1 0 37920 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_391
timestamp 1621261055
transform 1 0 38688 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_399
timestamp 1621261055
transform 1 0 39456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_349
timestamp 1621261055
transform 1 0 40800 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_402
timestamp 1621261055
transform 1 0 39744 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_410
timestamp 1621261055
transform 1 0 40512 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_418
timestamp 1621261055
transform 1 0 41280 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_407
timestamp 1621261055
transform 1 0 40224 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_411
timestamp 1621261055
transform 1 0 40608 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_414
timestamp 1621261055
transform 1 0 40896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_339
timestamp 1621261055
transform 1 0 43392 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_426
timestamp 1621261055
transform 1 0 42048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_434
timestamp 1621261055
transform 1 0 42816 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_438
timestamp 1621261055
transform 1 0 43200 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_441
timestamp 1621261055
transform 1 0 43488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_422
timestamp 1621261055
transform 1 0 41664 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_430
timestamp 1621261055
transform 1 0 42432 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_438
timestamp 1621261055
transform 1 0 43200 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _187_
timestamp 1621261055
transform 1 0 44928 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_15_449
timestamp 1621261055
transform 1 0 44256 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_457
timestamp 1621261055
transform 1 0 45024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_446
timestamp 1621261055
transform 1 0 43968 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_454
timestamp 1621261055
transform 1 0 44736 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_459
timestamp 1621261055
transform 1 0 45216 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_350
timestamp 1621261055
transform 1 0 46080 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_465
timestamp 1621261055
transform 1 0 45792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_473
timestamp 1621261055
transform 1 0 46560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_481
timestamp 1621261055
transform 1 0 47328 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_16_467
timestamp 1621261055
transform 1 0 45984 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_469
timestamp 1621261055
transform 1 0 46176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_477
timestamp 1621261055
transform 1 0 46944 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_340
timestamp 1621261055
transform 1 0 48672 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_489
timestamp 1621261055
transform 1 0 48096 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_493
timestamp 1621261055
transform 1 0 48480 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_496
timestamp 1621261055
transform 1 0 48768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_504
timestamp 1621261055
transform 1 0 49536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_485
timestamp 1621261055
transform 1 0 47712 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_493
timestamp 1621261055
transform 1 0 48480 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_501
timestamp 1621261055
transform 1 0 49248 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_351
timestamp 1621261055
transform 1 0 51360 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_512
timestamp 1621261055
transform 1 0 50304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_520
timestamp 1621261055
transform 1 0 51072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_509
timestamp 1621261055
transform 1 0 50016 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_517
timestamp 1621261055
transform 1 0 50784 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_521
timestamp 1621261055
transform 1 0 51168 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_524
timestamp 1621261055
transform 1 0 51456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_528
timestamp 1621261055
transform 1 0 51840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_536
timestamp 1621261055
transform 1 0 52608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_544
timestamp 1621261055
transform 1 0 53376 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_532
timestamp 1621261055
transform 1 0 52224 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_540
timestamp 1621261055
transform 1 0 52992 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_341
timestamp 1621261055
transform 1 0 53952 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_548
timestamp 1621261055
transform 1 0 53760 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_551
timestamp 1621261055
transform 1 0 54048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_559
timestamp 1621261055
transform 1 0 54816 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_567
timestamp 1621261055
transform 1 0 55584 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_548
timestamp 1621261055
transform 1 0 53760 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_556
timestamp 1621261055
transform 1 0 54528 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_564
timestamp 1621261055
transform 1 0 55296 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_576
timestamp 1621261055
transform 1 0 56448 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_572
timestamp 1621261055
transform 1 0 56064 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_15_575
timestamp 1621261055
transform 1 0 56352 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_579
timestamp 1621261055
transform 1 0 56736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_584
timestamp 1621261055
transform 1 0 57216 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_18
timestamp 1621261055
transform 1 0 56736 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_352
timestamp 1621261055
transform 1 0 56640 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _011_
timestamp 1621261055
transform 1 0 56928 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_587
timestamp 1621261055
transform 1 0 57504 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _180_
timestamp 1621261055
transform 1 0 57600 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_31
timestamp 1621261055
transform -1 0 58848 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_33
timestamp 1621261055
transform -1 0 58848 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_15_591
timestamp 1621261055
transform 1 0 57888 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_595
timestamp 1621261055
transform 1 0 58272 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_595
timestamp 1621261055
transform 1 0 58272 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_34
timestamp 1621261055
transform 1 0 1152 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_4
timestamp 1621261055
transform 1 0 1536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_12
timestamp 1621261055
transform 1 0 2304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_20
timestamp 1621261055
transform 1 0 3072 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_28
timestamp 1621261055
transform 1 0 3840 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_36
timestamp 1621261055
transform 1 0 4608 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_353
timestamp 1621261055
transform 1 0 6432 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_44
timestamp 1621261055
transform 1 0 5376 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_52
timestamp 1621261055
transform 1 0 6144 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_54
timestamp 1621261055
transform 1 0 6336 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_56
timestamp 1621261055
transform 1 0 6528 0 1 13986
box -38 -49 806 715
use INVX2  INVX2
timestamp 1624074425
transform 1 0 7680 0 1 13986
box 0 -48 576 714
use sky130_fd_sc_ls__diode_2  ANTENNA_61
timestamp 1621261055
transform 1 0 7488 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_64
timestamp 1621261055
transform 1 0 7296 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_74
timestamp 1621261055
transform 1 0 8256 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_82
timestamp 1621261055
transform 1 0 9024 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_90
timestamp 1621261055
transform 1 0 9792 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_98
timestamp 1621261055
transform 1 0 10560 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_354
timestamp 1621261055
transform 1 0 11712 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_106
timestamp 1621261055
transform 1 0 11328 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_111
timestamp 1621261055
transform 1 0 11808 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_119
timestamp 1621261055
transform 1 0 12576 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_127
timestamp 1621261055
transform 1 0 13344 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_135
timestamp 1621261055
transform 1 0 14112 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_143
timestamp 1621261055
transform 1 0 14880 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_355
timestamp 1621261055
transform 1 0 16992 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_151
timestamp 1621261055
transform 1 0 15648 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_159
timestamp 1621261055
transform 1 0 16416 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_163
timestamp 1621261055
transform 1 0 16800 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_166
timestamp 1621261055
transform 1 0 17088 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_174
timestamp 1621261055
transform 1 0 17856 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_182
timestamp 1621261055
transform 1 0 18624 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_190
timestamp 1621261055
transform 1 0 19392 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_198
timestamp 1621261055
transform 1 0 20160 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_206
timestamp 1621261055
transform 1 0 20928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_356
timestamp 1621261055
transform 1 0 22272 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_214
timestamp 1621261055
transform 1 0 21696 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_218
timestamp 1621261055
transform 1 0 22080 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_221
timestamp 1621261055
transform 1 0 22368 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_229
timestamp 1621261055
transform 1 0 23136 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_237
timestamp 1621261055
transform 1 0 23904 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_245
timestamp 1621261055
transform 1 0 24672 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_253
timestamp 1621261055
transform 1 0 25440 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_261
timestamp 1621261055
transform 1 0 26208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_269
timestamp 1621261055
transform 1 0 26976 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_273
timestamp 1621261055
transform 1 0 27360 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_357
timestamp 1621261055
transform 1 0 27552 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_276
timestamp 1621261055
transform 1 0 27648 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_284
timestamp 1621261055
transform 1 0 28416 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_292
timestamp 1621261055
transform 1 0 29184 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_300
timestamp 1621261055
transform 1 0 29952 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_308
timestamp 1621261055
transform 1 0 30720 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_358
timestamp 1621261055
transform 1 0 32832 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_316
timestamp 1621261055
transform 1 0 31488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_324
timestamp 1621261055
transform 1 0 32256 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_328
timestamp 1621261055
transform 1 0 32640 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_331
timestamp 1621261055
transform 1 0 32928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_339
timestamp 1621261055
transform 1 0 33696 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_347
timestamp 1621261055
transform 1 0 34464 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_355
timestamp 1621261055
transform 1 0 35232 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_363
timestamp 1621261055
transform 1 0 36000 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_371
timestamp 1621261055
transform 1 0 36768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_359
timestamp 1621261055
transform 1 0 38112 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_379
timestamp 1621261055
transform 1 0 37536 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_383
timestamp 1621261055
transform 1 0 37920 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_386
timestamp 1621261055
transform 1 0 38208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_394
timestamp 1621261055
transform 1 0 38976 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_402
timestamp 1621261055
transform 1 0 39744 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_410
timestamp 1621261055
transform 1 0 40512 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_418
timestamp 1621261055
transform 1 0 41280 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_360
timestamp 1621261055
transform 1 0 43392 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_426
timestamp 1621261055
transform 1 0 42048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_434
timestamp 1621261055
transform 1 0 42816 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_438
timestamp 1621261055
transform 1 0 43200 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_17_441
timestamp 1621261055
transform 1 0 43488 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _176_
timestamp 1621261055
transform 1 0 44160 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_445
timestamp 1621261055
transform 1 0 43872 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_447
timestamp 1621261055
transform 1 0 44064 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_451
timestamp 1621261055
transform 1 0 44448 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_459
timestamp 1621261055
transform 1 0 45216 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_467
timestamp 1621261055
transform 1 0 45984 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_475
timestamp 1621261055
transform 1 0 46752 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_483
timestamp 1621261055
transform 1 0 47520 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_361
timestamp 1621261055
transform 1 0 48672 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_491
timestamp 1621261055
transform 1 0 48288 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_496
timestamp 1621261055
transform 1 0 48768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_504
timestamp 1621261055
transform 1 0 49536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _128_
timestamp 1621261055
transform 1 0 50976 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_17_512
timestamp 1621261055
transform 1 0 50304 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_516
timestamp 1621261055
transform 1 0 50688 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_518
timestamp 1621261055
transform 1 0 50880 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_522
timestamp 1621261055
transform 1 0 51264 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_530
timestamp 1621261055
transform 1 0 52032 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_538
timestamp 1621261055
transform 1 0 52800 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_546
timestamp 1621261055
transform 1 0 53568 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_362
timestamp 1621261055
transform 1 0 53952 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_551
timestamp 1621261055
transform 1 0 54048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_559
timestamp 1621261055
transform 1 0 54816 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_567
timestamp 1621261055
transform 1 0 55584 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_575
timestamp 1621261055
transform 1 0 56352 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_583
timestamp 1621261055
transform 1 0 57120 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_35
timestamp 1621261055
transform -1 0 58848 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_17_591
timestamp 1621261055
transform 1 0 57888 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_595
timestamp 1621261055
transform 1 0 58272 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_36
timestamp 1621261055
transform 1 0 1152 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_18_4
timestamp 1621261055
transform 1 0 1536 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_12
timestamp 1621261055
transform 1 0 2304 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_20
timestamp 1621261055
transform 1 0 3072 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_363
timestamp 1621261055
transform 1 0 3840 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_29
timestamp 1621261055
transform 1 0 3936 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_37
timestamp 1621261055
transform 1 0 4704 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_45
timestamp 1621261055
transform 1 0 5472 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_53
timestamp 1621261055
transform 1 0 6240 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_61
timestamp 1621261055
transform 1 0 7008 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_364
timestamp 1621261055
transform 1 0 9120 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_69
timestamp 1621261055
transform 1 0 7776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_77
timestamp 1621261055
transform 1 0 8544 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_81
timestamp 1621261055
transform 1 0 8928 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_84
timestamp 1621261055
transform 1 0 9216 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_92
timestamp 1621261055
transform 1 0 9984 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_100
timestamp 1621261055
transform 1 0 10752 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_108
timestamp 1621261055
transform 1 0 11520 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_116
timestamp 1621261055
transform 1 0 12288 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_124
timestamp 1621261055
transform 1 0 13056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _069_
timestamp 1621261055
transform 1 0 14880 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_365
timestamp 1621261055
transform 1 0 14400 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_132
timestamp 1621261055
transform 1 0 13824 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_136
timestamp 1621261055
transform 1 0 14208 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_18_139
timestamp 1621261055
transform 1 0 14496 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_18_146
timestamp 1621261055
transform 1 0 15168 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_154
timestamp 1621261055
transform 1 0 15936 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_162
timestamp 1621261055
transform 1 0 16704 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _084_
timestamp 1621261055
transform 1 0 18048 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_18_170
timestamp 1621261055
transform 1 0 17472 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_174
timestamp 1621261055
transform 1 0 17856 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_179
timestamp 1621261055
transform 1 0 18336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_187
timestamp 1621261055
transform 1 0 19104 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_366
timestamp 1621261055
transform 1 0 19680 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_191
timestamp 1621261055
transform 1 0 19488 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_194
timestamp 1621261055
transform 1 0 19776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_202
timestamp 1621261055
transform 1 0 20544 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_210
timestamp 1621261055
transform 1 0 21312 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_218
timestamp 1621261055
transform 1 0 22080 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_226
timestamp 1621261055
transform 1 0 22848 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_367
timestamp 1621261055
transform 1 0 24960 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_234
timestamp 1621261055
transform 1 0 23616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_242
timestamp 1621261055
transform 1 0 24384 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_246
timestamp 1621261055
transform 1 0 24768 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_249
timestamp 1621261055
transform 1 0 25056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_257
timestamp 1621261055
transform 1 0 25824 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_265
timestamp 1621261055
transform 1 0 26592 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_273
timestamp 1621261055
transform 1 0 27360 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_281
timestamp 1621261055
transform 1 0 28128 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_289
timestamp 1621261055
transform 1 0 28896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_368
timestamp 1621261055
transform 1 0 30240 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_297
timestamp 1621261055
transform 1 0 29664 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_301
timestamp 1621261055
transform 1 0 30048 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_304
timestamp 1621261055
transform 1 0 30336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_312
timestamp 1621261055
transform 1 0 31104 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_320
timestamp 1621261055
transform 1 0 31872 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_328
timestamp 1621261055
transform 1 0 32640 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_336
timestamp 1621261055
transform 1 0 33408 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_344
timestamp 1621261055
transform 1 0 34176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_352
timestamp 1621261055
transform 1 0 34944 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_356
timestamp 1621261055
transform 1 0 35328 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_369
timestamp 1621261055
transform 1 0 35520 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_359
timestamp 1621261055
transform 1 0 35616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_367
timestamp 1621261055
transform 1 0 36384 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_375
timestamp 1621261055
transform 1 0 37152 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_383
timestamp 1621261055
transform 1 0 37920 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_391
timestamp 1621261055
transform 1 0 38688 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_399
timestamp 1621261055
transform 1 0 39456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_370
timestamp 1621261055
transform 1 0 40800 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_407
timestamp 1621261055
transform 1 0 40224 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_411
timestamp 1621261055
transform 1 0 40608 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_414
timestamp 1621261055
transform 1 0 40896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_422
timestamp 1621261055
transform 1 0 41664 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_430
timestamp 1621261055
transform 1 0 42432 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_438
timestamp 1621261055
transform 1 0 43200 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_446
timestamp 1621261055
transform 1 0 43968 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_454
timestamp 1621261055
transform 1 0 44736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_462
timestamp 1621261055
transform 1 0 45504 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_371
timestamp 1621261055
transform 1 0 46080 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_466
timestamp 1621261055
transform 1 0 45888 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_469
timestamp 1621261055
transform 1 0 46176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_477
timestamp 1621261055
transform 1 0 46944 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_485
timestamp 1621261055
transform 1 0 47712 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_493
timestamp 1621261055
transform 1 0 48480 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_501
timestamp 1621261055
transform 1 0 49248 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_372
timestamp 1621261055
transform 1 0 51360 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_509
timestamp 1621261055
transform 1 0 50016 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_517
timestamp 1621261055
transform 1 0 50784 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_521
timestamp 1621261055
transform 1 0 51168 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_524
timestamp 1621261055
transform 1 0 51456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_532
timestamp 1621261055
transform 1 0 52224 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_540
timestamp 1621261055
transform 1 0 52992 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_548
timestamp 1621261055
transform 1 0 53760 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_556
timestamp 1621261055
transform 1 0 54528 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_564
timestamp 1621261055
transform 1 0 55296 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_373
timestamp 1621261055
transform 1 0 56640 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_572
timestamp 1621261055
transform 1 0 56064 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_576
timestamp 1621261055
transform 1 0 56448 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_579
timestamp 1621261055
transform 1 0 56736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_587
timestamp 1621261055
transform 1 0 57504 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_37
timestamp 1621261055
transform -1 0 58848 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_595
timestamp 1621261055
transform 1 0 58272 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_38
timestamp 1621261055
transform 1 0 1152 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_4
timestamp 1621261055
transform 1 0 1536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_12
timestamp 1621261055
transform 1 0 2304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_20
timestamp 1621261055
transform 1 0 3072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_28
timestamp 1621261055
transform 1 0 3840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_36
timestamp 1621261055
transform 1 0 4608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_374
timestamp 1621261055
transform 1 0 6432 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_44
timestamp 1621261055
transform 1 0 5376 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_52
timestamp 1621261055
transform 1 0 6144 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_54
timestamp 1621261055
transform 1 0 6336 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_56
timestamp 1621261055
transform 1 0 6528 0 1 15318
box -38 -49 806 715
use INVX4  INVX4
timestamp 1624074425
transform 1 0 7680 0 1 15318
box 0 -48 864 714
use sky130_fd_sc_ls__diode_2  ANTENNA_65
timestamp 1621261055
transform 1 0 7488 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_64
timestamp 1621261055
transform 1 0 7296 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_77
timestamp 1621261055
transform 1 0 8544 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_85
timestamp 1621261055
transform 1 0 9312 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_93
timestamp 1621261055
transform 1 0 10080 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_101
timestamp 1621261055
transform 1 0 10848 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_375
timestamp 1621261055
transform 1 0 11712 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_19_109
timestamp 1621261055
transform 1 0 11616 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_111
timestamp 1621261055
transform 1 0 11808 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_119
timestamp 1621261055
transform 1 0 12576 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_127
timestamp 1621261055
transform 1 0 13344 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_135
timestamp 1621261055
transform 1 0 14112 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_143
timestamp 1621261055
transform 1 0 14880 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_376
timestamp 1621261055
transform 1 0 16992 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_151
timestamp 1621261055
transform 1 0 15648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_159
timestamp 1621261055
transform 1 0 16416 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_163
timestamp 1621261055
transform 1 0 16800 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_166
timestamp 1621261055
transform 1 0 17088 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _003_
timestamp 1621261055
transform -1 0 19584 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_8
timestamp 1621261055
transform -1 0 19296 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_174
timestamp 1621261055
transform 1 0 17856 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_182
timestamp 1621261055
transform 1 0 18624 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_19_186
timestamp 1621261055
transform 1 0 19008 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_192
timestamp 1621261055
transform 1 0 19584 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_200
timestamp 1621261055
transform 1 0 20352 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_208
timestamp 1621261055
transform 1 0 21120 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_377
timestamp 1621261055
transform 1 0 22272 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_216
timestamp 1621261055
transform 1 0 21888 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_221
timestamp 1621261055
transform 1 0 22368 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_229
timestamp 1621261055
transform 1 0 23136 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_237
timestamp 1621261055
transform 1 0 23904 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_245
timestamp 1621261055
transform 1 0 24672 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_253
timestamp 1621261055
transform 1 0 25440 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_261
timestamp 1621261055
transform 1 0 26208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_269
timestamp 1621261055
transform 1 0 26976 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_273
timestamp 1621261055
transform 1 0 27360 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_378
timestamp 1621261055
transform 1 0 27552 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_276
timestamp 1621261055
transform 1 0 27648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_284
timestamp 1621261055
transform 1 0 28416 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_292
timestamp 1621261055
transform 1 0 29184 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_300
timestamp 1621261055
transform 1 0 29952 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_308
timestamp 1621261055
transform 1 0 30720 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_379
timestamp 1621261055
transform 1 0 32832 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_316
timestamp 1621261055
transform 1 0 31488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_324
timestamp 1621261055
transform 1 0 32256 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_328
timestamp 1621261055
transform 1 0 32640 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_331
timestamp 1621261055
transform 1 0 32928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_339
timestamp 1621261055
transform 1 0 33696 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_347
timestamp 1621261055
transform 1 0 34464 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_355
timestamp 1621261055
transform 1 0 35232 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_363
timestamp 1621261055
transform 1 0 36000 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_371
timestamp 1621261055
transform 1 0 36768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_380
timestamp 1621261055
transform 1 0 38112 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_379
timestamp 1621261055
transform 1 0 37536 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_383
timestamp 1621261055
transform 1 0 37920 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_386
timestamp 1621261055
transform 1 0 38208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_394
timestamp 1621261055
transform 1 0 38976 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_402
timestamp 1621261055
transform 1 0 39744 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_410
timestamp 1621261055
transform 1 0 40512 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_418
timestamp 1621261055
transform 1 0 41280 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_381
timestamp 1621261055
transform 1 0 43392 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_426
timestamp 1621261055
transform 1 0 42048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_434
timestamp 1621261055
transform 1 0 42816 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_438
timestamp 1621261055
transform 1 0 43200 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_441
timestamp 1621261055
transform 1 0 43488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_449
timestamp 1621261055
transform 1 0 44256 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_457
timestamp 1621261055
transform 1 0 45024 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_465
timestamp 1621261055
transform 1 0 45792 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_473
timestamp 1621261055
transform 1 0 46560 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_481
timestamp 1621261055
transform 1 0 47328 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_382
timestamp 1621261055
transform 1 0 48672 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_489
timestamp 1621261055
transform 1 0 48096 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_493
timestamp 1621261055
transform 1 0 48480 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_496
timestamp 1621261055
transform 1 0 48768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_504
timestamp 1621261055
transform 1 0 49536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_512
timestamp 1621261055
transform 1 0 50304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_520
timestamp 1621261055
transform 1 0 51072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_528
timestamp 1621261055
transform 1 0 51840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_536
timestamp 1621261055
transform 1 0 52608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_544
timestamp 1621261055
transform 1 0 53376 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _044_
timestamp 1621261055
transform -1 0 55776 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_383
timestamp 1621261055
transform 1 0 53952 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_41
timestamp 1621261055
transform -1 0 55488 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_548
timestamp 1621261055
transform 1 0 53760 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_551
timestamp 1621261055
transform 1 0 54048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_559
timestamp 1621261055
transform 1 0 54816 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_19_563
timestamp 1621261055
transform 1 0 55200 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_569
timestamp 1621261055
transform 1 0 55776 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_577
timestamp 1621261055
transform 1 0 56544 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_585
timestamp 1621261055
transform 1 0 57312 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_39
timestamp 1621261055
transform -1 0 58848 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_19_593
timestamp 1621261055
transform 1 0 58080 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_40
timestamp 1621261055
transform 1 0 1152 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_20_4
timestamp 1621261055
transform 1 0 1536 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_12
timestamp 1621261055
transform 1 0 2304 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_20
timestamp 1621261055
transform 1 0 3072 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_384
timestamp 1621261055
transform 1 0 3840 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_29
timestamp 1621261055
transform 1 0 3936 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_37
timestamp 1621261055
transform 1 0 4704 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_45
timestamp 1621261055
transform 1 0 5472 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_53
timestamp 1621261055
transform 1 0 6240 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_61
timestamp 1621261055
transform 1 0 7008 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_385
timestamp 1621261055
transform 1 0 9120 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_69
timestamp 1621261055
transform 1 0 7776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_77
timestamp 1621261055
transform 1 0 8544 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_81
timestamp 1621261055
transform 1 0 8928 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_84
timestamp 1621261055
transform 1 0 9216 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_92
timestamp 1621261055
transform 1 0 9984 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_100
timestamp 1621261055
transform 1 0 10752 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_108
timestamp 1621261055
transform 1 0 11520 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_116
timestamp 1621261055
transform 1 0 12288 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_124
timestamp 1621261055
transform 1 0 13056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_386
timestamp 1621261055
transform 1 0 14400 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_132
timestamp 1621261055
transform 1 0 13824 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_136
timestamp 1621261055
transform 1 0 14208 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_139
timestamp 1621261055
transform 1 0 14496 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_147
timestamp 1621261055
transform 1 0 15264 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_155
timestamp 1621261055
transform 1 0 16032 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_163
timestamp 1621261055
transform 1 0 16800 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_171
timestamp 1621261055
transform 1 0 17568 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_179
timestamp 1621261055
transform 1 0 18336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_187
timestamp 1621261055
transform 1 0 19104 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_387
timestamp 1621261055
transform 1 0 19680 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_191
timestamp 1621261055
transform 1 0 19488 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_194
timestamp 1621261055
transform 1 0 19776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_202
timestamp 1621261055
transform 1 0 20544 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_210
timestamp 1621261055
transform 1 0 21312 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_218
timestamp 1621261055
transform 1 0 22080 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_226
timestamp 1621261055
transform 1 0 22848 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_388
timestamp 1621261055
transform 1 0 24960 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_234
timestamp 1621261055
transform 1 0 23616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_242
timestamp 1621261055
transform 1 0 24384 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_246
timestamp 1621261055
transform 1 0 24768 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_249
timestamp 1621261055
transform 1 0 25056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_257
timestamp 1621261055
transform 1 0 25824 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_265
timestamp 1621261055
transform 1 0 26592 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_273
timestamp 1621261055
transform 1 0 27360 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_281
timestamp 1621261055
transform 1 0 28128 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_289
timestamp 1621261055
transform 1 0 28896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_389
timestamp 1621261055
transform 1 0 30240 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_297
timestamp 1621261055
transform 1 0 29664 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_301
timestamp 1621261055
transform 1 0 30048 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_304
timestamp 1621261055
transform 1 0 30336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_312
timestamp 1621261055
transform 1 0 31104 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_320
timestamp 1621261055
transform 1 0 31872 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_328
timestamp 1621261055
transform 1 0 32640 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_336
timestamp 1621261055
transform 1 0 33408 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_344
timestamp 1621261055
transform 1 0 34176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_352
timestamp 1621261055
transform 1 0 34944 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_356
timestamp 1621261055
transform 1 0 35328 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_390
timestamp 1621261055
transform 1 0 35520 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_359
timestamp 1621261055
transform 1 0 35616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_367
timestamp 1621261055
transform 1 0 36384 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_375
timestamp 1621261055
transform 1 0 37152 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_383
timestamp 1621261055
transform 1 0 37920 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_391
timestamp 1621261055
transform 1 0 38688 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_399
timestamp 1621261055
transform 1 0 39456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_391
timestamp 1621261055
transform 1 0 40800 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_407
timestamp 1621261055
transform 1 0 40224 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_411
timestamp 1621261055
transform 1 0 40608 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_414
timestamp 1621261055
transform 1 0 40896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_422
timestamp 1621261055
transform 1 0 41664 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_430
timestamp 1621261055
transform 1 0 42432 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_438
timestamp 1621261055
transform 1 0 43200 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_446
timestamp 1621261055
transform 1 0 43968 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_454
timestamp 1621261055
transform 1 0 44736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_462
timestamp 1621261055
transform 1 0 45504 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_392
timestamp 1621261055
transform 1 0 46080 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_466
timestamp 1621261055
transform 1 0 45888 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_469
timestamp 1621261055
transform 1 0 46176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_477
timestamp 1621261055
transform 1 0 46944 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_485
timestamp 1621261055
transform 1 0 47712 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_493
timestamp 1621261055
transform 1 0 48480 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_501
timestamp 1621261055
transform 1 0 49248 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_393
timestamp 1621261055
transform 1 0 51360 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_509
timestamp 1621261055
transform 1 0 50016 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_517
timestamp 1621261055
transform 1 0 50784 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_521
timestamp 1621261055
transform 1 0 51168 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_524
timestamp 1621261055
transform 1 0 51456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_532
timestamp 1621261055
transform 1 0 52224 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_540
timestamp 1621261055
transform 1 0 52992 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_548
timestamp 1621261055
transform 1 0 53760 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_556
timestamp 1621261055
transform 1 0 54528 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_564
timestamp 1621261055
transform 1 0 55296 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_394
timestamp 1621261055
transform 1 0 56640 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_572
timestamp 1621261055
transform 1 0 56064 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_576
timestamp 1621261055
transform 1 0 56448 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_579
timestamp 1621261055
transform 1 0 56736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_587
timestamp 1621261055
transform 1 0 57504 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_41
timestamp 1621261055
transform -1 0 58848 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_595
timestamp 1621261055
transform 1 0 58272 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_42
timestamp 1621261055
transform 1 0 1152 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_21_4
timestamp 1621261055
transform 1 0 1536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_12
timestamp 1621261055
transform 1 0 2304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_20
timestamp 1621261055
transform 1 0 3072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_28
timestamp 1621261055
transform 1 0 3840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_36
timestamp 1621261055
transform 1 0 4608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_395
timestamp 1621261055
transform 1 0 6432 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_44
timestamp 1621261055
transform 1 0 5376 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_52
timestamp 1621261055
transform 1 0 6144 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_21_54
timestamp 1621261055
transform 1 0 6336 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_56
timestamp 1621261055
transform 1 0 6528 0 1 16650
box -38 -49 806 715
use INVX8  INVX8
timestamp 1624074425
transform 1 0 7680 0 1 16650
box 0 -48 1440 714
use sky130_fd_sc_ls__diode_2  ANTENNA_68
timestamp 1621261055
transform 1 0 7488 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_64
timestamp 1621261055
transform 1 0 7296 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_83
timestamp 1621261055
transform 1 0 9120 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_91
timestamp 1621261055
transform 1 0 9888 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_99
timestamp 1621261055
transform 1 0 10656 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_396
timestamp 1621261055
transform 1 0 11712 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_107
timestamp 1621261055
transform 1 0 11424 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_21_109
timestamp 1621261055
transform 1 0 11616 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_111
timestamp 1621261055
transform 1 0 11808 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_119
timestamp 1621261055
transform 1 0 12576 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_127
timestamp 1621261055
transform 1 0 13344 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_135
timestamp 1621261055
transform 1 0 14112 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_143
timestamp 1621261055
transform 1 0 14880 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_397
timestamp 1621261055
transform 1 0 16992 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_151
timestamp 1621261055
transform 1 0 15648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_159
timestamp 1621261055
transform 1 0 16416 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_163
timestamp 1621261055
transform 1 0 16800 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_166
timestamp 1621261055
transform 1 0 17088 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_174
timestamp 1621261055
transform 1 0 17856 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_182
timestamp 1621261055
transform 1 0 18624 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_190
timestamp 1621261055
transform 1 0 19392 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_198
timestamp 1621261055
transform 1 0 20160 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_206
timestamp 1621261055
transform 1 0 20928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_398
timestamp 1621261055
transform 1 0 22272 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_214
timestamp 1621261055
transform 1 0 21696 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_218
timestamp 1621261055
transform 1 0 22080 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_221
timestamp 1621261055
transform 1 0 22368 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_229
timestamp 1621261055
transform 1 0 23136 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_237
timestamp 1621261055
transform 1 0 23904 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_245
timestamp 1621261055
transform 1 0 24672 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_253
timestamp 1621261055
transform 1 0 25440 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_261
timestamp 1621261055
transform 1 0 26208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_269
timestamp 1621261055
transform 1 0 26976 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_273
timestamp 1621261055
transform 1 0 27360 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_399
timestamp 1621261055
transform 1 0 27552 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_276
timestamp 1621261055
transform 1 0 27648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_284
timestamp 1621261055
transform 1 0 28416 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_292
timestamp 1621261055
transform 1 0 29184 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _081_
timestamp 1621261055
transform 1 0 30240 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_300
timestamp 1621261055
transform 1 0 29952 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_21_302
timestamp 1621261055
transform 1 0 30144 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_306
timestamp 1621261055
transform 1 0 30528 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_314
timestamp 1621261055
transform 1 0 31296 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_400
timestamp 1621261055
transform 1 0 32832 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_322
timestamp 1621261055
transform 1 0 32064 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_331
timestamp 1621261055
transform 1 0 32928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_339
timestamp 1621261055
transform 1 0 33696 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_347
timestamp 1621261055
transform 1 0 34464 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_355
timestamp 1621261055
transform 1 0 35232 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_363
timestamp 1621261055
transform 1 0 36000 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_371
timestamp 1621261055
transform 1 0 36768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_401
timestamp 1621261055
transform 1 0 38112 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_379
timestamp 1621261055
transform 1 0 37536 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_383
timestamp 1621261055
transform 1 0 37920 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_386
timestamp 1621261055
transform 1 0 38208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_394
timestamp 1621261055
transform 1 0 38976 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_402
timestamp 1621261055
transform 1 0 39744 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_410
timestamp 1621261055
transform 1 0 40512 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_418
timestamp 1621261055
transform 1 0 41280 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_402
timestamp 1621261055
transform 1 0 43392 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_426
timestamp 1621261055
transform 1 0 42048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_434
timestamp 1621261055
transform 1 0 42816 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_438
timestamp 1621261055
transform 1 0 43200 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_441
timestamp 1621261055
transform 1 0 43488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_449
timestamp 1621261055
transform 1 0 44256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_457
timestamp 1621261055
transform 1 0 45024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_465
timestamp 1621261055
transform 1 0 45792 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_473
timestamp 1621261055
transform 1 0 46560 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_481
timestamp 1621261055
transform 1 0 47328 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_403
timestamp 1621261055
transform 1 0 48672 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_489
timestamp 1621261055
transform 1 0 48096 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_493
timestamp 1621261055
transform 1 0 48480 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_496
timestamp 1621261055
transform 1 0 48768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_504
timestamp 1621261055
transform 1 0 49536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_512
timestamp 1621261055
transform 1 0 50304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_520
timestamp 1621261055
transform 1 0 51072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_528
timestamp 1621261055
transform 1 0 51840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_536
timestamp 1621261055
transform 1 0 52608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_544
timestamp 1621261055
transform 1 0 53376 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_404
timestamp 1621261055
transform 1 0 53952 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_548
timestamp 1621261055
transform 1 0 53760 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_551
timestamp 1621261055
transform 1 0 54048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_559
timestamp 1621261055
transform 1 0 54816 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_567
timestamp 1621261055
transform 1 0 55584 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_575
timestamp 1621261055
transform 1 0 56352 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_583
timestamp 1621261055
transform 1 0 57120 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_43
timestamp 1621261055
transform -1 0 58848 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_21_591
timestamp 1621261055
transform 1 0 57888 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_595
timestamp 1621261055
transform 1 0 58272 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _151_
timestamp 1621261055
transform 1 0 1536 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_44
timestamp 1621261055
transform 1 0 1152 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_22_7
timestamp 1621261055
transform 1 0 1824 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_15
timestamp 1621261055
transform 1 0 2592 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_405
timestamp 1621261055
transform 1 0 3840 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_23
timestamp 1621261055
transform 1 0 3360 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_22_27
timestamp 1621261055
transform 1 0 3744 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_29
timestamp 1621261055
transform 1 0 3936 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_37
timestamp 1621261055
transform 1 0 4704 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_45
timestamp 1621261055
transform 1 0 5472 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_53
timestamp 1621261055
transform 1 0 6240 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_61
timestamp 1621261055
transform 1 0 7008 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_406
timestamp 1621261055
transform 1 0 9120 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_69
timestamp 1621261055
transform 1 0 7776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_77
timestamp 1621261055
transform 1 0 8544 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_81
timestamp 1621261055
transform 1 0 8928 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_84
timestamp 1621261055
transform 1 0 9216 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_92
timestamp 1621261055
transform 1 0 9984 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_100
timestamp 1621261055
transform 1 0 10752 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_108
timestamp 1621261055
transform 1 0 11520 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_116
timestamp 1621261055
transform 1 0 12288 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_124
timestamp 1621261055
transform 1 0 13056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_407
timestamp 1621261055
transform 1 0 14400 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_132
timestamp 1621261055
transform 1 0 13824 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_136
timestamp 1621261055
transform 1 0 14208 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_139
timestamp 1621261055
transform 1 0 14496 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_147
timestamp 1621261055
transform 1 0 15264 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_155
timestamp 1621261055
transform 1 0 16032 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_163
timestamp 1621261055
transform 1 0 16800 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_171
timestamp 1621261055
transform 1 0 17568 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_179
timestamp 1621261055
transform 1 0 18336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_187
timestamp 1621261055
transform 1 0 19104 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_408
timestamp 1621261055
transform 1 0 19680 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_191
timestamp 1621261055
transform 1 0 19488 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_194
timestamp 1621261055
transform 1 0 19776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_202
timestamp 1621261055
transform 1 0 20544 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_210
timestamp 1621261055
transform 1 0 21312 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_218
timestamp 1621261055
transform 1 0 22080 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_226
timestamp 1621261055
transform 1 0 22848 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_409
timestamp 1621261055
transform 1 0 24960 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_234
timestamp 1621261055
transform 1 0 23616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_242
timestamp 1621261055
transform 1 0 24384 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_246
timestamp 1621261055
transform 1 0 24768 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_249
timestamp 1621261055
transform 1 0 25056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_257
timestamp 1621261055
transform 1 0 25824 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_265
timestamp 1621261055
transform 1 0 26592 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_273
timestamp 1621261055
transform 1 0 27360 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_281
timestamp 1621261055
transform 1 0 28128 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_289
timestamp 1621261055
transform 1 0 28896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_410
timestamp 1621261055
transform 1 0 30240 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_297
timestamp 1621261055
transform 1 0 29664 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_301
timestamp 1621261055
transform 1 0 30048 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_304
timestamp 1621261055
transform 1 0 30336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_312
timestamp 1621261055
transform 1 0 31104 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_320
timestamp 1621261055
transform 1 0 31872 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_328
timestamp 1621261055
transform 1 0 32640 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_336
timestamp 1621261055
transform 1 0 33408 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_344
timestamp 1621261055
transform 1 0 34176 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_352
timestamp 1621261055
transform 1 0 34944 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_356
timestamp 1621261055
transform 1 0 35328 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_411
timestamp 1621261055
transform 1 0 35520 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_359
timestamp 1621261055
transform 1 0 35616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_367
timestamp 1621261055
transform 1 0 36384 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_375
timestamp 1621261055
transform 1 0 37152 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_383
timestamp 1621261055
transform 1 0 37920 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_391
timestamp 1621261055
transform 1 0 38688 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_399
timestamp 1621261055
transform 1 0 39456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_412
timestamp 1621261055
transform 1 0 40800 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_407
timestamp 1621261055
transform 1 0 40224 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_411
timestamp 1621261055
transform 1 0 40608 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_414
timestamp 1621261055
transform 1 0 40896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_422
timestamp 1621261055
transform 1 0 41664 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_430
timestamp 1621261055
transform 1 0 42432 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_438
timestamp 1621261055
transform 1 0 43200 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_446
timestamp 1621261055
transform 1 0 43968 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_454
timestamp 1621261055
transform 1 0 44736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_462
timestamp 1621261055
transform 1 0 45504 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_413
timestamp 1621261055
transform 1 0 46080 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_466
timestamp 1621261055
transform 1 0 45888 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_469
timestamp 1621261055
transform 1 0 46176 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_477
timestamp 1621261055
transform 1 0 46944 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_485
timestamp 1621261055
transform 1 0 47712 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_493
timestamp 1621261055
transform 1 0 48480 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_501
timestamp 1621261055
transform 1 0 49248 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_414
timestamp 1621261055
transform 1 0 51360 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_509
timestamp 1621261055
transform 1 0 50016 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_517
timestamp 1621261055
transform 1 0 50784 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_521
timestamp 1621261055
transform 1 0 51168 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_524
timestamp 1621261055
transform 1 0 51456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_532
timestamp 1621261055
transform 1 0 52224 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_540
timestamp 1621261055
transform 1 0 52992 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_548
timestamp 1621261055
transform 1 0 53760 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_556
timestamp 1621261055
transform 1 0 54528 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_564
timestamp 1621261055
transform 1 0 55296 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_415
timestamp 1621261055
transform 1 0 56640 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_572
timestamp 1621261055
transform 1 0 56064 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_576
timestamp 1621261055
transform 1 0 56448 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_579
timestamp 1621261055
transform 1 0 56736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_587
timestamp 1621261055
transform 1 0 57504 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_45
timestamp 1621261055
transform -1 0 58848 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_595
timestamp 1621261055
transform 1 0 58272 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_46
timestamp 1621261055
transform 1 0 1152 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_48
timestamp 1621261055
transform 1 0 1152 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_4
timestamp 1621261055
transform 1 0 1536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_12
timestamp 1621261055
transform 1 0 2304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_20
timestamp 1621261055
transform 1 0 3072 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_4
timestamp 1621261055
transform 1 0 1536 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_12
timestamp 1621261055
transform 1 0 2304 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_20
timestamp 1621261055
transform 1 0 3072 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_426
timestamp 1621261055
transform 1 0 3840 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_28
timestamp 1621261055
transform 1 0 3840 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_36
timestamp 1621261055
transform 1 0 4608 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_29
timestamp 1621261055
transform 1 0 3936 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_37
timestamp 1621261055
transform 1 0 4704 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_416
timestamp 1621261055
transform 1 0 6432 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_44
timestamp 1621261055
transform 1 0 5376 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_52
timestamp 1621261055
transform 1 0 6144 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_23_54
timestamp 1621261055
transform 1 0 6336 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_56
timestamp 1621261055
transform 1 0 6528 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_45
timestamp 1621261055
transform 1 0 5472 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_53
timestamp 1621261055
transform 1 0 6240 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_61
timestamp 1621261055
transform 1 0 7008 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_69
timestamp 1621261055
transform 1 0 7776 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_64
timestamp 1621261055
transform 1 0 7296 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_73
timestamp 1621261055
transform 1 0 7488 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _077_
timestamp 1621261055
transform 1 0 8160 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_84
timestamp 1621261055
transform 1 0 9216 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_24_82
timestamp 1621261055
transform 1 0 9024 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_80
timestamp 1621261055
transform 1 0 8832 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_76
timestamp 1621261055
transform 1 0 8448 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_427
timestamp 1621261055
transform 1 0 9120 0 -1 19314
box -38 -49 134 715
use MUX2X1  MUX2X1
timestamp 1624074425
transform 1 0 7680 0 1 17982
box 0 -48 1728 714
use sky130_fd_sc_ls__decap_8  FILLER_23_86
timestamp 1621261055
transform 1 0 9408 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_94
timestamp 1621261055
transform 1 0 10176 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_102
timestamp 1621261055
transform 1 0 10944 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_92
timestamp 1621261055
transform 1 0 9984 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_100
timestamp 1621261055
transform 1 0 10752 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_417
timestamp 1621261055
transform 1 0 11712 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_111
timestamp 1621261055
transform 1 0 11808 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_119
timestamp 1621261055
transform 1 0 12576 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_108
timestamp 1621261055
transform 1 0 11520 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_116
timestamp 1621261055
transform 1 0 12288 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_124
timestamp 1621261055
transform 1 0 13056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_428
timestamp 1621261055
transform 1 0 14400 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_127
timestamp 1621261055
transform 1 0 13344 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_135
timestamp 1621261055
transform 1 0 14112 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_143
timestamp 1621261055
transform 1 0 14880 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_132
timestamp 1621261055
transform 1 0 13824 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_136
timestamp 1621261055
transform 1 0 14208 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_139
timestamp 1621261055
transform 1 0 14496 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_147
timestamp 1621261055
transform 1 0 15264 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_418
timestamp 1621261055
transform 1 0 16992 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_151
timestamp 1621261055
transform 1 0 15648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_159
timestamp 1621261055
transform 1 0 16416 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_163
timestamp 1621261055
transform 1 0 16800 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_166
timestamp 1621261055
transform 1 0 17088 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_155
timestamp 1621261055
transform 1 0 16032 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_163
timestamp 1621261055
transform 1 0 16800 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_174
timestamp 1621261055
transform 1 0 17856 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_182
timestamp 1621261055
transform 1 0 18624 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_171
timestamp 1621261055
transform 1 0 17568 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_179
timestamp 1621261055
transform 1 0 18336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_187
timestamp 1621261055
transform 1 0 19104 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_194
timestamp 1621261055
transform 1 0 19776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_191
timestamp 1621261055
transform 1 0 19488 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_190
timestamp 1621261055
transform 1 0 19392 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_429
timestamp 1621261055
transform 1 0 19680 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_202
timestamp 1621261055
transform 1 0 20544 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_204
timestamp 1621261055
transform 1 0 20736 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_200
timestamp 1621261055
transform 1 0 20352 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_198
timestamp 1621261055
transform 1 0 20160 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _206_
timestamp 1621261055
transform 1 0 20448 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_210
timestamp 1621261055
transform 1 0 21312 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_419
timestamp 1621261055
transform 1 0 22272 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_212
timestamp 1621261055
transform 1 0 21504 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_221
timestamp 1621261055
transform 1 0 22368 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_229
timestamp 1621261055
transform 1 0 23136 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_218
timestamp 1621261055
transform 1 0 22080 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_226
timestamp 1621261055
transform 1 0 22848 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _049_
timestamp 1621261055
transform 1 0 24480 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_430
timestamp 1621261055
transform 1 0 24960 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_59
timestamp 1621261055
transform 1 0 24288 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_237
timestamp 1621261055
transform 1 0 23904 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_246
timestamp 1621261055
transform 1 0 24768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_234
timestamp 1621261055
transform 1 0 23616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_242
timestamp 1621261055
transform 1 0 24384 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_246
timestamp 1621261055
transform 1 0 24768 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_249
timestamp 1621261055
transform 1 0 25056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_254
timestamp 1621261055
transform 1 0 25536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_262
timestamp 1621261055
transform 1 0 26304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_270
timestamp 1621261055
transform 1 0 27072 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_257
timestamp 1621261055
transform 1 0 25824 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_265
timestamp 1621261055
transform 1 0 26592 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_273
timestamp 1621261055
transform 1 0 27360 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_420
timestamp 1621261055
transform 1 0 27552 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_23_274
timestamp 1621261055
transform 1 0 27456 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_276
timestamp 1621261055
transform 1 0 27648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_284
timestamp 1621261055
transform 1 0 28416 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_292
timestamp 1621261055
transform 1 0 29184 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_281
timestamp 1621261055
transform 1 0 28128 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_289
timestamp 1621261055
transform 1 0 28896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_431
timestamp 1621261055
transform 1 0 30240 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_300
timestamp 1621261055
transform 1 0 29952 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_308
timestamp 1621261055
transform 1 0 30720 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_297
timestamp 1621261055
transform 1 0 29664 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_301
timestamp 1621261055
transform 1 0 30048 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_304
timestamp 1621261055
transform 1 0 30336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_312
timestamp 1621261055
transform 1 0 31104 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_421
timestamp 1621261055
transform 1 0 32832 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_316
timestamp 1621261055
transform 1 0 31488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_324
timestamp 1621261055
transform 1 0 32256 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_328
timestamp 1621261055
transform 1 0 32640 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_331
timestamp 1621261055
transform 1 0 32928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_320
timestamp 1621261055
transform 1 0 31872 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_328
timestamp 1621261055
transform 1 0 32640 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_336
timestamp 1621261055
transform 1 0 33408 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_339
timestamp 1621261055
transform 1 0 33696 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_347
timestamp 1621261055
transform 1 0 34464 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_355
timestamp 1621261055
transform 1 0 35232 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_344
timestamp 1621261055
transform 1 0 34176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_352
timestamp 1621261055
transform 1 0 34944 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_356
timestamp 1621261055
transform 1 0 35328 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_432
timestamp 1621261055
transform 1 0 35520 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_363
timestamp 1621261055
transform 1 0 36000 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_371
timestamp 1621261055
transform 1 0 36768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_359
timestamp 1621261055
transform 1 0 35616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_367
timestamp 1621261055
transform 1 0 36384 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_375
timestamp 1621261055
transform 1 0 37152 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_422
timestamp 1621261055
transform 1 0 38112 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_23_379
timestamp 1621261055
transform 1 0 37536 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_383
timestamp 1621261055
transform 1 0 37920 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_386
timestamp 1621261055
transform 1 0 38208 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_394
timestamp 1621261055
transform 1 0 38976 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_383
timestamp 1621261055
transform 1 0 37920 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_391
timestamp 1621261055
transform 1 0 38688 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_399
timestamp 1621261055
transform 1 0 39456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_433
timestamp 1621261055
transform 1 0 40800 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_402
timestamp 1621261055
transform 1 0 39744 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_410
timestamp 1621261055
transform 1 0 40512 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_418
timestamp 1621261055
transform 1 0 41280 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_407
timestamp 1621261055
transform 1 0 40224 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_411
timestamp 1621261055
transform 1 0 40608 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_414
timestamp 1621261055
transform 1 0 40896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_423
timestamp 1621261055
transform 1 0 43392 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_426
timestamp 1621261055
transform 1 0 42048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_434
timestamp 1621261055
transform 1 0 42816 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_438
timestamp 1621261055
transform 1 0 43200 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_441
timestamp 1621261055
transform 1 0 43488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_422
timestamp 1621261055
transform 1 0 41664 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_430
timestamp 1621261055
transform 1 0 42432 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_438
timestamp 1621261055
transform 1 0 43200 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_449
timestamp 1621261055
transform 1 0 44256 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_457
timestamp 1621261055
transform 1 0 45024 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_446
timestamp 1621261055
transform 1 0 43968 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_454
timestamp 1621261055
transform 1 0 44736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_462
timestamp 1621261055
transform 1 0 45504 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_434
timestamp 1621261055
transform 1 0 46080 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_465
timestamp 1621261055
transform 1 0 45792 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_473
timestamp 1621261055
transform 1 0 46560 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_481
timestamp 1621261055
transform 1 0 47328 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_466
timestamp 1621261055
transform 1 0 45888 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_469
timestamp 1621261055
transform 1 0 46176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_477
timestamp 1621261055
transform 1 0 46944 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_424
timestamp 1621261055
transform 1 0 48672 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_23_489
timestamp 1621261055
transform 1 0 48096 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_493
timestamp 1621261055
transform 1 0 48480 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_496
timestamp 1621261055
transform 1 0 48768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_504
timestamp 1621261055
transform 1 0 49536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_485
timestamp 1621261055
transform 1 0 47712 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_493
timestamp 1621261055
transform 1 0 48480 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_501
timestamp 1621261055
transform 1 0 49248 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _152_
timestamp 1621261055
transform 1 0 51456 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_435
timestamp 1621261055
transform 1 0 51360 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_512
timestamp 1621261055
transform 1 0 50304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_520
timestamp 1621261055
transform 1 0 51072 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_509
timestamp 1621261055
transform 1 0 50016 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_517
timestamp 1621261055
transform 1 0 50784 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_521
timestamp 1621261055
transform 1 0 51168 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_524
timestamp 1621261055
transform 1 0 51456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_527
timestamp 1621261055
transform 1 0 51744 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_535
timestamp 1621261055
transform 1 0 52512 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_543
timestamp 1621261055
transform 1 0 53280 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_532
timestamp 1621261055
transform 1 0 52224 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_540
timestamp 1621261055
transform 1 0 52992 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_425
timestamp 1621261055
transform 1 0 53952 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_547
timestamp 1621261055
transform 1 0 53664 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_23_549
timestamp 1621261055
transform 1 0 53856 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_551
timestamp 1621261055
transform 1 0 54048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_559
timestamp 1621261055
transform 1 0 54816 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_567
timestamp 1621261055
transform 1 0 55584 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_548
timestamp 1621261055
transform 1 0 53760 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_556
timestamp 1621261055
transform 1 0 54528 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_564
timestamp 1621261055
transform 1 0 55296 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_436
timestamp 1621261055
transform 1 0 56640 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_575
timestamp 1621261055
transform 1 0 56352 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_583
timestamp 1621261055
transform 1 0 57120 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_572
timestamp 1621261055
transform 1 0 56064 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_576
timestamp 1621261055
transform 1 0 56448 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_579
timestamp 1621261055
transform 1 0 56736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_587
timestamp 1621261055
transform 1 0 57504 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_47
timestamp 1621261055
transform -1 0 58848 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_49
timestamp 1621261055
transform -1 0 58848 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_23_591
timestamp 1621261055
transform 1 0 57888 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_595
timestamp 1621261055
transform 1 0 58272 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_595
timestamp 1621261055
transform 1 0 58272 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_50
timestamp 1621261055
transform 1 0 1152 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_4
timestamp 1621261055
transform 1 0 1536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_12
timestamp 1621261055
transform 1 0 2304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_20
timestamp 1621261055
transform 1 0 3072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_28
timestamp 1621261055
transform 1 0 3840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_36
timestamp 1621261055
transform 1 0 4608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_437
timestamp 1621261055
transform 1 0 6432 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_44
timestamp 1621261055
transform 1 0 5376 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_52
timestamp 1621261055
transform 1 0 6144 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_54
timestamp 1621261055
transform 1 0 6336 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_56
timestamp 1621261055
transform 1 0 6528 0 1 19314
box -38 -49 806 715
use NAND2X1  NAND2X1
timestamp 1624074425
transform 1 0 7680 0 1 19314
box 0 -48 864 714
use sky130_fd_sc_ls__diode_2  ANTENNA_77
timestamp 1621261055
transform 1 0 7488 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_64
timestamp 1621261055
transform 1 0 7296 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_77
timestamp 1621261055
transform 1 0 8544 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_85
timestamp 1621261055
transform 1 0 9312 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_93
timestamp 1621261055
transform 1 0 10080 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_101
timestamp 1621261055
transform 1 0 10848 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_438
timestamp 1621261055
transform 1 0 11712 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_25_109
timestamp 1621261055
transform 1 0 11616 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_111
timestamp 1621261055
transform 1 0 11808 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_119
timestamp 1621261055
transform 1 0 12576 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_127
timestamp 1621261055
transform 1 0 13344 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_135
timestamp 1621261055
transform 1 0 14112 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_143
timestamp 1621261055
transform 1 0 14880 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_439
timestamp 1621261055
transform 1 0 16992 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_151
timestamp 1621261055
transform 1 0 15648 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_159
timestamp 1621261055
transform 1 0 16416 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_163
timestamp 1621261055
transform 1 0 16800 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_166
timestamp 1621261055
transform 1 0 17088 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_174
timestamp 1621261055
transform 1 0 17856 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_182
timestamp 1621261055
transform 1 0 18624 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_190
timestamp 1621261055
transform 1 0 19392 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_198
timestamp 1621261055
transform 1 0 20160 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_206
timestamp 1621261055
transform 1 0 20928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_440
timestamp 1621261055
transform 1 0 22272 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_214
timestamp 1621261055
transform 1 0 21696 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_218
timestamp 1621261055
transform 1 0 22080 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_221
timestamp 1621261055
transform 1 0 22368 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_229
timestamp 1621261055
transform 1 0 23136 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_237
timestamp 1621261055
transform 1 0 23904 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_245
timestamp 1621261055
transform 1 0 24672 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_253
timestamp 1621261055
transform 1 0 25440 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_261
timestamp 1621261055
transform 1 0 26208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_269
timestamp 1621261055
transform 1 0 26976 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_273
timestamp 1621261055
transform 1 0 27360 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_441
timestamp 1621261055
transform 1 0 27552 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_276
timestamp 1621261055
transform 1 0 27648 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_284
timestamp 1621261055
transform 1 0 28416 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_292
timestamp 1621261055
transform 1 0 29184 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_300
timestamp 1621261055
transform 1 0 29952 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_308
timestamp 1621261055
transform 1 0 30720 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_442
timestamp 1621261055
transform 1 0 32832 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_316
timestamp 1621261055
transform 1 0 31488 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_324
timestamp 1621261055
transform 1 0 32256 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_328
timestamp 1621261055
transform 1 0 32640 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_331
timestamp 1621261055
transform 1 0 32928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_339
timestamp 1621261055
transform 1 0 33696 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_347
timestamp 1621261055
transform 1 0 34464 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_355
timestamp 1621261055
transform 1 0 35232 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_363
timestamp 1621261055
transform 1 0 36000 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_371
timestamp 1621261055
transform 1 0 36768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_443
timestamp 1621261055
transform 1 0 38112 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_379
timestamp 1621261055
transform 1 0 37536 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_383
timestamp 1621261055
transform 1 0 37920 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_386
timestamp 1621261055
transform 1 0 38208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_394
timestamp 1621261055
transform 1 0 38976 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_402
timestamp 1621261055
transform 1 0 39744 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_410
timestamp 1621261055
transform 1 0 40512 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_418
timestamp 1621261055
transform 1 0 41280 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_444
timestamp 1621261055
transform 1 0 43392 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_426
timestamp 1621261055
transform 1 0 42048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_434
timestamp 1621261055
transform 1 0 42816 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_438
timestamp 1621261055
transform 1 0 43200 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_25_441
timestamp 1621261055
transform 1 0 43488 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _089_
timestamp 1621261055
transform 1 0 43872 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_25_448
timestamp 1621261055
transform 1 0 44160 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_456
timestamp 1621261055
transform 1 0 44928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_464
timestamp 1621261055
transform 1 0 45696 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_472
timestamp 1621261055
transform 1 0 46464 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_480
timestamp 1621261055
transform 1 0 47232 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_445
timestamp 1621261055
transform 1 0 48672 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_488
timestamp 1621261055
transform 1 0 48000 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_492
timestamp 1621261055
transform 1 0 48384 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_494
timestamp 1621261055
transform 1 0 48576 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_496
timestamp 1621261055
transform 1 0 48768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_504
timestamp 1621261055
transform 1 0 49536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_512
timestamp 1621261055
transform 1 0 50304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_520
timestamp 1621261055
transform 1 0 51072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_528
timestamp 1621261055
transform 1 0 51840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_536
timestamp 1621261055
transform 1 0 52608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_544
timestamp 1621261055
transform 1 0 53376 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_446
timestamp 1621261055
transform 1 0 53952 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_548
timestamp 1621261055
transform 1 0 53760 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_551
timestamp 1621261055
transform 1 0 54048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_559
timestamp 1621261055
transform 1 0 54816 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_567
timestamp 1621261055
transform 1 0 55584 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_575
timestamp 1621261055
transform 1 0 56352 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_583
timestamp 1621261055
transform 1 0 57120 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_51
timestamp 1621261055
transform -1 0 58848 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_25_591
timestamp 1621261055
transform 1 0 57888 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_595
timestamp 1621261055
transform 1 0 58272 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_52
timestamp 1621261055
transform 1 0 1152 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_26_4
timestamp 1621261055
transform 1 0 1536 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_12
timestamp 1621261055
transform 1 0 2304 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_20
timestamp 1621261055
transform 1 0 3072 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_447
timestamp 1621261055
transform 1 0 3840 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_29
timestamp 1621261055
transform 1 0 3936 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_37
timestamp 1621261055
transform 1 0 4704 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_45
timestamp 1621261055
transform 1 0 5472 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_53
timestamp 1621261055
transform 1 0 6240 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_61
timestamp 1621261055
transform 1 0 7008 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_448
timestamp 1621261055
transform 1 0 9120 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_69
timestamp 1621261055
transform 1 0 7776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_77
timestamp 1621261055
transform 1 0 8544 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_81
timestamp 1621261055
transform 1 0 8928 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_84
timestamp 1621261055
transform 1 0 9216 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_92
timestamp 1621261055
transform 1 0 9984 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_100
timestamp 1621261055
transform 1 0 10752 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_108
timestamp 1621261055
transform 1 0 11520 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_116
timestamp 1621261055
transform 1 0 12288 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_124
timestamp 1621261055
transform 1 0 13056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_449
timestamp 1621261055
transform 1 0 14400 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_132
timestamp 1621261055
transform 1 0 13824 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_136
timestamp 1621261055
transform 1 0 14208 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_139
timestamp 1621261055
transform 1 0 14496 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_147
timestamp 1621261055
transform 1 0 15264 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_155
timestamp 1621261055
transform 1 0 16032 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_163
timestamp 1621261055
transform 1 0 16800 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_171
timestamp 1621261055
transform 1 0 17568 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_179
timestamp 1621261055
transform 1 0 18336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_187
timestamp 1621261055
transform 1 0 19104 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_450
timestamp 1621261055
transform 1 0 19680 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_191
timestamp 1621261055
transform 1 0 19488 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_194
timestamp 1621261055
transform 1 0 19776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_202
timestamp 1621261055
transform 1 0 20544 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_210
timestamp 1621261055
transform 1 0 21312 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_218
timestamp 1621261055
transform 1 0 22080 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_226
timestamp 1621261055
transform 1 0 22848 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_451
timestamp 1621261055
transform 1 0 24960 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_234
timestamp 1621261055
transform 1 0 23616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_242
timestamp 1621261055
transform 1 0 24384 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_246
timestamp 1621261055
transform 1 0 24768 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_249
timestamp 1621261055
transform 1 0 25056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _181_
timestamp 1621261055
transform 1 0 26880 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_257
timestamp 1621261055
transform 1 0 25824 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_265
timestamp 1621261055
transform 1 0 26592 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_267
timestamp 1621261055
transform 1 0 26784 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_271
timestamp 1621261055
transform 1 0 27168 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_279
timestamp 1621261055
transform 1 0 27936 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_287
timestamp 1621261055
transform 1 0 28704 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_452
timestamp 1621261055
transform 1 0 30240 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_295
timestamp 1621261055
transform 1 0 29472 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_304
timestamp 1621261055
transform 1 0 30336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_312
timestamp 1621261055
transform 1 0 31104 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_320
timestamp 1621261055
transform 1 0 31872 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_328
timestamp 1621261055
transform 1 0 32640 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_336
timestamp 1621261055
transform 1 0 33408 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_344
timestamp 1621261055
transform 1 0 34176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_352
timestamp 1621261055
transform 1 0 34944 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_356
timestamp 1621261055
transform 1 0 35328 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_453
timestamp 1621261055
transform 1 0 35520 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_359
timestamp 1621261055
transform 1 0 35616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_367
timestamp 1621261055
transform 1 0 36384 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_375
timestamp 1621261055
transform 1 0 37152 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _004_
timestamp 1621261055
transform 1 0 37920 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_386
timestamp 1621261055
transform 1 0 38208 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_394
timestamp 1621261055
transform 1 0 38976 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_454
timestamp 1621261055
transform 1 0 40800 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_402
timestamp 1621261055
transform 1 0 39744 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_410
timestamp 1621261055
transform 1 0 40512 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_412
timestamp 1621261055
transform 1 0 40704 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_414
timestamp 1621261055
transform 1 0 40896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_422
timestamp 1621261055
transform 1 0 41664 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_430
timestamp 1621261055
transform 1 0 42432 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_438
timestamp 1621261055
transform 1 0 43200 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_446
timestamp 1621261055
transform 1 0 43968 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_454
timestamp 1621261055
transform 1 0 44736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_462
timestamp 1621261055
transform 1 0 45504 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_455
timestamp 1621261055
transform 1 0 46080 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_466
timestamp 1621261055
transform 1 0 45888 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_469
timestamp 1621261055
transform 1 0 46176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_477
timestamp 1621261055
transform 1 0 46944 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_485
timestamp 1621261055
transform 1 0 47712 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_493
timestamp 1621261055
transform 1 0 48480 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_501
timestamp 1621261055
transform 1 0 49248 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_456
timestamp 1621261055
transform 1 0 51360 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_509
timestamp 1621261055
transform 1 0 50016 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_517
timestamp 1621261055
transform 1 0 50784 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_521
timestamp 1621261055
transform 1 0 51168 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_524
timestamp 1621261055
transform 1 0 51456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _138_
timestamp 1621261055
transform 1 0 52800 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_26_532
timestamp 1621261055
transform 1 0 52224 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_536
timestamp 1621261055
transform 1 0 52608 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_541
timestamp 1621261055
transform 1 0 53088 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_549
timestamp 1621261055
transform 1 0 53856 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_557
timestamp 1621261055
transform 1 0 54624 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_565
timestamp 1621261055
transform 1 0 55392 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_457
timestamp 1621261055
transform 1 0 56640 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_573
timestamp 1621261055
transform 1 0 56160 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_26_577
timestamp 1621261055
transform 1 0 56544 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_579
timestamp 1621261055
transform 1 0 56736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_587
timestamp 1621261055
transform 1 0 57504 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_53
timestamp 1621261055
transform -1 0 58848 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_595
timestamp 1621261055
transform 1 0 58272 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_54
timestamp 1621261055
transform 1 0 1152 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_4
timestamp 1621261055
transform 1 0 1536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_12
timestamp 1621261055
transform 1 0 2304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_20
timestamp 1621261055
transform 1 0 3072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_28
timestamp 1621261055
transform 1 0 3840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_36
timestamp 1621261055
transform 1 0 4608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_458
timestamp 1621261055
transform 1 0 6432 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_44
timestamp 1621261055
transform 1 0 5376 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_52
timestamp 1621261055
transform 1 0 6144 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_54
timestamp 1621261055
transform 1 0 6336 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_56
timestamp 1621261055
transform 1 0 6528 0 1 20646
box -38 -49 806 715
use NAND3X1  NAND3X1
timestamp 1624074425
transform 1 0 7680 0 1 20646
box 0 -48 1152 714
use sky130_fd_sc_ls__diode_2  ANTENNA_83
timestamp 1621261055
transform 1 0 7488 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_64
timestamp 1621261055
transform 1 0 7296 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_80
timestamp 1621261055
transform 1 0 8832 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_88
timestamp 1621261055
transform 1 0 9600 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_96
timestamp 1621261055
transform 1 0 10368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_104
timestamp 1621261055
transform 1 0 11136 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_459
timestamp 1621261055
transform 1 0 11712 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_108
timestamp 1621261055
transform 1 0 11520 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_111
timestamp 1621261055
transform 1 0 11808 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_119
timestamp 1621261055
transform 1 0 12576 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_127
timestamp 1621261055
transform 1 0 13344 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_135
timestamp 1621261055
transform 1 0 14112 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_143
timestamp 1621261055
transform 1 0 14880 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_147
timestamp 1621261055
transform 1 0 15264 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _210_
timestamp 1621261055
transform 1 0 15552 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_460
timestamp 1621261055
transform 1 0 16992 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_27_149
timestamp 1621261055
transform 1 0 15456 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_153
timestamp 1621261055
transform 1 0 15840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_161
timestamp 1621261055
transform 1 0 16608 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_166
timestamp 1621261055
transform 1 0 17088 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_174
timestamp 1621261055
transform 1 0 17856 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_182
timestamp 1621261055
transform 1 0 18624 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_190
timestamp 1621261055
transform 1 0 19392 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_198
timestamp 1621261055
transform 1 0 20160 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_206
timestamp 1621261055
transform 1 0 20928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_461
timestamp 1621261055
transform 1 0 22272 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_214
timestamp 1621261055
transform 1 0 21696 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_218
timestamp 1621261055
transform 1 0 22080 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_221
timestamp 1621261055
transform 1 0 22368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_229
timestamp 1621261055
transform 1 0 23136 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_237
timestamp 1621261055
transform 1 0 23904 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_245
timestamp 1621261055
transform 1 0 24672 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_253
timestamp 1621261055
transform 1 0 25440 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_261
timestamp 1621261055
transform 1 0 26208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_269
timestamp 1621261055
transform 1 0 26976 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_273
timestamp 1621261055
transform 1 0 27360 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _148_
timestamp 1621261055
transform 1 0 28032 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_462
timestamp 1621261055
transform 1 0 27552 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_276
timestamp 1621261055
transform 1 0 27648 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_283
timestamp 1621261055
transform 1 0 28320 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_291
timestamp 1621261055
transform 1 0 29088 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_299
timestamp 1621261055
transform 1 0 29856 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_307
timestamp 1621261055
transform 1 0 30624 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_315
timestamp 1621261055
transform 1 0 31392 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_463
timestamp 1621261055
transform 1 0 32832 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_323
timestamp 1621261055
transform 1 0 32160 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_327
timestamp 1621261055
transform 1 0 32544 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_329
timestamp 1621261055
transform 1 0 32736 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_331
timestamp 1621261055
transform 1 0 32928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_339
timestamp 1621261055
transform 1 0 33696 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_347
timestamp 1621261055
transform 1 0 34464 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_355
timestamp 1621261055
transform 1 0 35232 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_363
timestamp 1621261055
transform 1 0 36000 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_371
timestamp 1621261055
transform 1 0 36768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_464
timestamp 1621261055
transform 1 0 38112 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_379
timestamp 1621261055
transform 1 0 37536 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_383
timestamp 1621261055
transform 1 0 37920 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_386
timestamp 1621261055
transform 1 0 38208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_394
timestamp 1621261055
transform 1 0 38976 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_402
timestamp 1621261055
transform 1 0 39744 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_410
timestamp 1621261055
transform 1 0 40512 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_418
timestamp 1621261055
transform 1 0 41280 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_465
timestamp 1621261055
transform 1 0 43392 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_426
timestamp 1621261055
transform 1 0 42048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_434
timestamp 1621261055
transform 1 0 42816 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_438
timestamp 1621261055
transform 1 0 43200 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_441
timestamp 1621261055
transform 1 0 43488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_449
timestamp 1621261055
transform 1 0 44256 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_457
timestamp 1621261055
transform 1 0 45024 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_465
timestamp 1621261055
transform 1 0 45792 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_473
timestamp 1621261055
transform 1 0 46560 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_481
timestamp 1621261055
transform 1 0 47328 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_466
timestamp 1621261055
transform 1 0 48672 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_489
timestamp 1621261055
transform 1 0 48096 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_493
timestamp 1621261055
transform 1 0 48480 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_496
timestamp 1621261055
transform 1 0 48768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_504
timestamp 1621261055
transform 1 0 49536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_512
timestamp 1621261055
transform 1 0 50304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_520
timestamp 1621261055
transform 1 0 51072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_528
timestamp 1621261055
transform 1 0 51840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_536
timestamp 1621261055
transform 1 0 52608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_544
timestamp 1621261055
transform 1 0 53376 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_467
timestamp 1621261055
transform 1 0 53952 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_548
timestamp 1621261055
transform 1 0 53760 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_551
timestamp 1621261055
transform 1 0 54048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_559
timestamp 1621261055
transform 1 0 54816 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_567
timestamp 1621261055
transform 1 0 55584 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_575
timestamp 1621261055
transform 1 0 56352 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_583
timestamp 1621261055
transform 1 0 57120 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_55
timestamp 1621261055
transform -1 0 58848 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_27_591
timestamp 1621261055
transform 1 0 57888 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_595
timestamp 1621261055
transform 1 0 58272 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_56
timestamp 1621261055
transform 1 0 1152 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_28_4
timestamp 1621261055
transform 1 0 1536 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_12
timestamp 1621261055
transform 1 0 2304 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_20
timestamp 1621261055
transform 1 0 3072 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_468
timestamp 1621261055
transform 1 0 3840 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_29
timestamp 1621261055
transform 1 0 3936 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_37
timestamp 1621261055
transform 1 0 4704 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_45
timestamp 1621261055
transform 1 0 5472 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_53
timestamp 1621261055
transform 1 0 6240 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_61
timestamp 1621261055
transform 1 0 7008 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_469
timestamp 1621261055
transform 1 0 9120 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_69
timestamp 1621261055
transform 1 0 7776 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_77
timestamp 1621261055
transform 1 0 8544 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_81
timestamp 1621261055
transform 1 0 8928 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_28_84
timestamp 1621261055
transform 1 0 9216 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _174_
timestamp 1621261055
transform 1 0 9600 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_28_91
timestamp 1621261055
transform 1 0 9888 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_99
timestamp 1621261055
transform 1 0 10656 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_107
timestamp 1621261055
transform 1 0 11424 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_115
timestamp 1621261055
transform 1 0 12192 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_123
timestamp 1621261055
transform 1 0 12960 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_470
timestamp 1621261055
transform 1 0 14400 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_131
timestamp 1621261055
transform 1 0 13728 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_135
timestamp 1621261055
transform 1 0 14112 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_28_137
timestamp 1621261055
transform 1 0 14304 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_139
timestamp 1621261055
transform 1 0 14496 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_147
timestamp 1621261055
transform 1 0 15264 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_155
timestamp 1621261055
transform 1 0 16032 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_163
timestamp 1621261055
transform 1 0 16800 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_171
timestamp 1621261055
transform 1 0 17568 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_179
timestamp 1621261055
transform 1 0 18336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_187
timestamp 1621261055
transform 1 0 19104 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _025_
timestamp 1621261055
transform 1 0 20640 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_471
timestamp 1621261055
transform 1 0 19680 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_4
timestamp 1621261055
transform 1 0 20448 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_191
timestamp 1621261055
transform 1 0 19488 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_28_194
timestamp 1621261055
transform 1 0 19776 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_198
timestamp 1621261055
transform 1 0 20160 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_28_200
timestamp 1621261055
transform 1 0 20352 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_206
timestamp 1621261055
transform 1 0 20928 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_214
timestamp 1621261055
transform 1 0 21696 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_222
timestamp 1621261055
transform 1 0 22464 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_230
timestamp 1621261055
transform 1 0 23232 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_472
timestamp 1621261055
transform 1 0 24960 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_238
timestamp 1621261055
transform 1 0 24000 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_246
timestamp 1621261055
transform 1 0 24768 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_249
timestamp 1621261055
transform 1 0 25056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_257
timestamp 1621261055
transform 1 0 25824 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_265
timestamp 1621261055
transform 1 0 26592 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_273
timestamp 1621261055
transform 1 0 27360 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_281
timestamp 1621261055
transform 1 0 28128 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_289
timestamp 1621261055
transform 1 0 28896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_473
timestamp 1621261055
transform 1 0 30240 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_297
timestamp 1621261055
transform 1 0 29664 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_301
timestamp 1621261055
transform 1 0 30048 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_304
timestamp 1621261055
transform 1 0 30336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_312
timestamp 1621261055
transform 1 0 31104 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_320
timestamp 1621261055
transform 1 0 31872 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_328
timestamp 1621261055
transform 1 0 32640 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_336
timestamp 1621261055
transform 1 0 33408 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_344
timestamp 1621261055
transform 1 0 34176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_352
timestamp 1621261055
transform 1 0 34944 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_356
timestamp 1621261055
transform 1 0 35328 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_474
timestamp 1621261055
transform 1 0 35520 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_359
timestamp 1621261055
transform 1 0 35616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_367
timestamp 1621261055
transform 1 0 36384 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_375
timestamp 1621261055
transform 1 0 37152 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_383
timestamp 1621261055
transform 1 0 37920 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_391
timestamp 1621261055
transform 1 0 38688 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_399
timestamp 1621261055
transform 1 0 39456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_475
timestamp 1621261055
transform 1 0 40800 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_407
timestamp 1621261055
transform 1 0 40224 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_411
timestamp 1621261055
transform 1 0 40608 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_414
timestamp 1621261055
transform 1 0 40896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_422
timestamp 1621261055
transform 1 0 41664 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_430
timestamp 1621261055
transform 1 0 42432 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_438
timestamp 1621261055
transform 1 0 43200 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_446
timestamp 1621261055
transform 1 0 43968 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_454
timestamp 1621261055
transform 1 0 44736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_462
timestamp 1621261055
transform 1 0 45504 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_476
timestamp 1621261055
transform 1 0 46080 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_466
timestamp 1621261055
transform 1 0 45888 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_469
timestamp 1621261055
transform 1 0 46176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_477
timestamp 1621261055
transform 1 0 46944 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_485
timestamp 1621261055
transform 1 0 47712 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_493
timestamp 1621261055
transform 1 0 48480 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_501
timestamp 1621261055
transform 1 0 49248 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_477
timestamp 1621261055
transform 1 0 51360 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_509
timestamp 1621261055
transform 1 0 50016 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_517
timestamp 1621261055
transform 1 0 50784 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_521
timestamp 1621261055
transform 1 0 51168 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_524
timestamp 1621261055
transform 1 0 51456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_532
timestamp 1621261055
transform 1 0 52224 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_540
timestamp 1621261055
transform 1 0 52992 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_548
timestamp 1621261055
transform 1 0 53760 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_556
timestamp 1621261055
transform 1 0 54528 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_564
timestamp 1621261055
transform 1 0 55296 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_478
timestamp 1621261055
transform 1 0 56640 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_572
timestamp 1621261055
transform 1 0 56064 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_576
timestamp 1621261055
transform 1 0 56448 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_579
timestamp 1621261055
transform 1 0 56736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_587
timestamp 1621261055
transform 1 0 57504 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_57
timestamp 1621261055
transform -1 0 58848 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_595
timestamp 1621261055
transform 1 0 58272 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_58
timestamp 1621261055
transform 1 0 1152 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_29_4
timestamp 1621261055
transform 1 0 1536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_12
timestamp 1621261055
transform 1 0 2304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_20
timestamp 1621261055
transform 1 0 3072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_28
timestamp 1621261055
transform 1 0 3840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_36
timestamp 1621261055
transform 1 0 4608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_479
timestamp 1621261055
transform 1 0 6432 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_44
timestamp 1621261055
transform 1 0 5376 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_52
timestamp 1621261055
transform 1 0 6144 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_54
timestamp 1621261055
transform 1 0 6336 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_56
timestamp 1621261055
transform 1 0 6528 0 1 21978
box -38 -49 806 715
use NOR2X1  NOR2X1
timestamp 1624074425
transform 1 0 7680 0 1 21978
box 0 -48 864 714
use sky130_fd_sc_ls__conb_1  _094_
timestamp 1621261055
transform 1 0 8928 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_29_64
timestamp 1621261055
transform 1 0 7296 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_29_77
timestamp 1621261055
transform 1 0 8544 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_29_84
timestamp 1621261055
transform 1 0 9216 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_92
timestamp 1621261055
transform 1 0 9984 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_100
timestamp 1621261055
transform 1 0 10752 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_480
timestamp 1621261055
transform 1 0 11712 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_108
timestamp 1621261055
transform 1 0 11520 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_111
timestamp 1621261055
transform 1 0 11808 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_119
timestamp 1621261055
transform 1 0 12576 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_127
timestamp 1621261055
transform 1 0 13344 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_135
timestamp 1621261055
transform 1 0 14112 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_143
timestamp 1621261055
transform 1 0 14880 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_481
timestamp 1621261055
transform 1 0 16992 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_151
timestamp 1621261055
transform 1 0 15648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_159
timestamp 1621261055
transform 1 0 16416 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_163
timestamp 1621261055
transform 1 0 16800 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_166
timestamp 1621261055
transform 1 0 17088 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_174
timestamp 1621261055
transform 1 0 17856 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_182
timestamp 1621261055
transform 1 0 18624 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_190
timestamp 1621261055
transform 1 0 19392 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_198
timestamp 1621261055
transform 1 0 20160 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_206
timestamp 1621261055
transform 1 0 20928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_482
timestamp 1621261055
transform 1 0 22272 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_214
timestamp 1621261055
transform 1 0 21696 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_218
timestamp 1621261055
transform 1 0 22080 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_221
timestamp 1621261055
transform 1 0 22368 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_229
timestamp 1621261055
transform 1 0 23136 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_237
timestamp 1621261055
transform 1 0 23904 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_245
timestamp 1621261055
transform 1 0 24672 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_253
timestamp 1621261055
transform 1 0 25440 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_261
timestamp 1621261055
transform 1 0 26208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_269
timestamp 1621261055
transform 1 0 26976 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_273
timestamp 1621261055
transform 1 0 27360 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_483
timestamp 1621261055
transform 1 0 27552 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_276
timestamp 1621261055
transform 1 0 27648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_284
timestamp 1621261055
transform 1 0 28416 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_292
timestamp 1621261055
transform 1 0 29184 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_300
timestamp 1621261055
transform 1 0 29952 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_308
timestamp 1621261055
transform 1 0 30720 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_484
timestamp 1621261055
transform 1 0 32832 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_316
timestamp 1621261055
transform 1 0 31488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_324
timestamp 1621261055
transform 1 0 32256 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_328
timestamp 1621261055
transform 1 0 32640 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_331
timestamp 1621261055
transform 1 0 32928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _191_
timestamp 1621261055
transform 1 0 34752 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_29_339
timestamp 1621261055
transform 1 0 33696 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_347
timestamp 1621261055
transform 1 0 34464 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_349
timestamp 1621261055
transform 1 0 34656 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_353
timestamp 1621261055
transform 1 0 35040 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _117_
timestamp 1621261055
transform 1 0 36288 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_29_361
timestamp 1621261055
transform 1 0 35808 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_29_365
timestamp 1621261055
transform 1 0 36192 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_369
timestamp 1621261055
transform 1 0 36576 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_377
timestamp 1621261055
transform 1 0 37344 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_485
timestamp 1621261055
transform 1 0 38112 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_386
timestamp 1621261055
transform 1 0 38208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_394
timestamp 1621261055
transform 1 0 38976 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_402
timestamp 1621261055
transform 1 0 39744 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_410
timestamp 1621261055
transform 1 0 40512 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_418
timestamp 1621261055
transform 1 0 41280 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_486
timestamp 1621261055
transform 1 0 43392 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_426
timestamp 1621261055
transform 1 0 42048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_434
timestamp 1621261055
transform 1 0 42816 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_438
timestamp 1621261055
transform 1 0 43200 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_441
timestamp 1621261055
transform 1 0 43488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_449
timestamp 1621261055
transform 1 0 44256 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_457
timestamp 1621261055
transform 1 0 45024 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_465
timestamp 1621261055
transform 1 0 45792 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_473
timestamp 1621261055
transform 1 0 46560 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_481
timestamp 1621261055
transform 1 0 47328 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_487
timestamp 1621261055
transform 1 0 48672 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_489
timestamp 1621261055
transform 1 0 48096 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_493
timestamp 1621261055
transform 1 0 48480 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_496
timestamp 1621261055
transform 1 0 48768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_504
timestamp 1621261055
transform 1 0 49536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_512
timestamp 1621261055
transform 1 0 50304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_520
timestamp 1621261055
transform 1 0 51072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_528
timestamp 1621261055
transform 1 0 51840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_536
timestamp 1621261055
transform 1 0 52608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_544
timestamp 1621261055
transform 1 0 53376 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_488
timestamp 1621261055
transform 1 0 53952 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_548
timestamp 1621261055
transform 1 0 53760 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_551
timestamp 1621261055
transform 1 0 54048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_559
timestamp 1621261055
transform 1 0 54816 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_567
timestamp 1621261055
transform 1 0 55584 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_575
timestamp 1621261055
transform 1 0 56352 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_583
timestamp 1621261055
transform 1 0 57120 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_59
timestamp 1621261055
transform -1 0 58848 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_29_591
timestamp 1621261055
transform 1 0 57888 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_595
timestamp 1621261055
transform 1 0 58272 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_60
timestamp 1621261055
transform 1 0 1152 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_62
timestamp 1621261055
transform 1 0 1152 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_4
timestamp 1621261055
transform 1 0 1536 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_12
timestamp 1621261055
transform 1 0 2304 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_20
timestamp 1621261055
transform 1 0 3072 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_4
timestamp 1621261055
transform 1 0 1536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_12
timestamp 1621261055
transform 1 0 2304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_20
timestamp 1621261055
transform 1 0 3072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_489
timestamp 1621261055
transform 1 0 3840 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_29
timestamp 1621261055
transform 1 0 3936 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_37
timestamp 1621261055
transform 1 0 4704 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_28
timestamp 1621261055
transform 1 0 3840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_36
timestamp 1621261055
transform 1 0 4608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_500
timestamp 1621261055
transform 1 0 6432 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_45
timestamp 1621261055
transform 1 0 5472 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_53
timestamp 1621261055
transform 1 0 6240 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_61
timestamp 1621261055
transform 1 0 7008 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_44
timestamp 1621261055
transform 1 0 5376 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_52
timestamp 1621261055
transform 1 0 6144 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_31_54
timestamp 1621261055
transform 1 0 6336 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_56
timestamp 1621261055
transform 1 0 6528 0 1 23310
box -38 -49 806 715
use OAI21X1  OAI21X1
timestamp 1624074425
transform 1 0 7680 0 1 23310
box 0 -48 1152 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_490
timestamp 1621261055
transform 1 0 9120 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_69
timestamp 1621261055
transform 1 0 7776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_77
timestamp 1621261055
transform 1 0 8544 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_81
timestamp 1621261055
transform 1 0 8928 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_84
timestamp 1621261055
transform 1 0 9216 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_64
timestamp 1621261055
transform 1 0 7296 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_80
timestamp 1621261055
transform 1 0 8832 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_92
timestamp 1621261055
transform 1 0 9984 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_100
timestamp 1621261055
transform 1 0 10752 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_88
timestamp 1621261055
transform 1 0 9600 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_96
timestamp 1621261055
transform 1 0 10368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_104
timestamp 1621261055
transform 1 0 11136 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _163_
timestamp 1621261055
transform 1 0 12192 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _201_
timestamp 1621261055
transform 1 0 13056 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_501
timestamp 1621261055
transform 1 0 11712 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_108
timestamp 1621261055
transform 1 0 11520 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_116
timestamp 1621261055
transform 1 0 12288 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_108
timestamp 1621261055
transform 1 0 11520 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_111
timestamp 1621261055
transform 1 0 11808 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_118
timestamp 1621261055
transform 1 0 12480 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_126
timestamp 1621261055
transform 1 0 13248 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_491
timestamp 1621261055
transform 1 0 14400 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_127
timestamp 1621261055
transform 1 0 13344 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_135
timestamp 1621261055
transform 1 0 14112 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_30_137
timestamp 1621261055
transform 1 0 14304 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_139
timestamp 1621261055
transform 1 0 14496 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_147
timestamp 1621261055
transform 1 0 15264 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_134
timestamp 1621261055
transform 1 0 14016 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_142
timestamp 1621261055
transform 1 0 14784 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_502
timestamp 1621261055
transform 1 0 16992 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_155
timestamp 1621261055
transform 1 0 16032 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_163
timestamp 1621261055
transform 1 0 16800 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_150
timestamp 1621261055
transform 1 0 15552 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_158
timestamp 1621261055
transform 1 0 16320 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_162
timestamp 1621261055
transform 1 0 16704 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_31_164
timestamp 1621261055
transform 1 0 16896 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_166
timestamp 1621261055
transform 1 0 17088 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_171
timestamp 1621261055
transform 1 0 17568 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_179
timestamp 1621261055
transform 1 0 18336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_187
timestamp 1621261055
transform 1 0 19104 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_174
timestamp 1621261055
transform 1 0 17856 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_182
timestamp 1621261055
transform 1 0 18624 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_492
timestamp 1621261055
transform 1 0 19680 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_191
timestamp 1621261055
transform 1 0 19488 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_194
timestamp 1621261055
transform 1 0 19776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_202
timestamp 1621261055
transform 1 0 20544 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_210
timestamp 1621261055
transform 1 0 21312 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_190
timestamp 1621261055
transform 1 0 19392 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_198
timestamp 1621261055
transform 1 0 20160 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_206
timestamp 1621261055
transform 1 0 20928 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_210
timestamp 1621261055
transform 1 0 21312 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _118_
timestamp 1621261055
transform 1 0 21504 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_503
timestamp 1621261055
transform 1 0 22272 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_218
timestamp 1621261055
transform 1 0 22080 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_226
timestamp 1621261055
transform 1 0 22848 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_215
timestamp 1621261055
transform 1 0 21792 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_31_219
timestamp 1621261055
transform 1 0 22176 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_221
timestamp 1621261055
transform 1 0 22368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_229
timestamp 1621261055
transform 1 0 23136 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_493
timestamp 1621261055
transform 1 0 24960 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_234
timestamp 1621261055
transform 1 0 23616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_242
timestamp 1621261055
transform 1 0 24384 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_246
timestamp 1621261055
transform 1 0 24768 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_249
timestamp 1621261055
transform 1 0 25056 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_237
timestamp 1621261055
transform 1 0 23904 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_245
timestamp 1621261055
transform 1 0 24672 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_257
timestamp 1621261055
transform 1 0 25824 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_265
timestamp 1621261055
transform 1 0 26592 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_273
timestamp 1621261055
transform 1 0 27360 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_253
timestamp 1621261055
transform 1 0 25440 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_261
timestamp 1621261055
transform 1 0 26208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_269
timestamp 1621261055
transform 1 0 26976 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_273
timestamp 1621261055
transform 1 0 27360 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_504
timestamp 1621261055
transform 1 0 27552 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_281
timestamp 1621261055
transform 1 0 28128 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_289
timestamp 1621261055
transform 1 0 28896 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_276
timestamp 1621261055
transform 1 0 27648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_284
timestamp 1621261055
transform 1 0 28416 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_292
timestamp 1621261055
transform 1 0 29184 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_494
timestamp 1621261055
transform 1 0 30240 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_297
timestamp 1621261055
transform 1 0 29664 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_301
timestamp 1621261055
transform 1 0 30048 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_304
timestamp 1621261055
transform 1 0 30336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_312
timestamp 1621261055
transform 1 0 31104 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_300
timestamp 1621261055
transform 1 0 29952 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_308
timestamp 1621261055
transform 1 0 30720 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_505
timestamp 1621261055
transform 1 0 32832 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_320
timestamp 1621261055
transform 1 0 31872 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_328
timestamp 1621261055
transform 1 0 32640 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_336
timestamp 1621261055
transform 1 0 33408 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_316
timestamp 1621261055
transform 1 0 31488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_324
timestamp 1621261055
transform 1 0 32256 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_328
timestamp 1621261055
transform 1 0 32640 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_331
timestamp 1621261055
transform 1 0 32928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _018_
timestamp 1621261055
transform 1 0 35232 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_29
timestamp 1621261055
transform 1 0 35040 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_344
timestamp 1621261055
transform 1 0 34176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_352
timestamp 1621261055
transform 1 0 34944 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_356
timestamp 1621261055
transform 1 0 35328 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_339
timestamp 1621261055
transform 1 0 33696 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_347
timestamp 1621261055
transform 1 0 34464 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_351
timestamp 1621261055
transform 1 0 34848 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_495
timestamp 1621261055
transform 1 0 35520 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_359
timestamp 1621261055
transform 1 0 35616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_367
timestamp 1621261055
transform 1 0 36384 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_375
timestamp 1621261055
transform 1 0 37152 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_358
timestamp 1621261055
transform 1 0 35520 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_366
timestamp 1621261055
transform 1 0 36288 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_374
timestamp 1621261055
transform 1 0 37056 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_506
timestamp 1621261055
transform 1 0 38112 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_383
timestamp 1621261055
transform 1 0 37920 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_391
timestamp 1621261055
transform 1 0 38688 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_399
timestamp 1621261055
transform 1 0 39456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_382
timestamp 1621261055
transform 1 0 37824 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_31_384
timestamp 1621261055
transform 1 0 38016 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_386
timestamp 1621261055
transform 1 0 38208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_394
timestamp 1621261055
transform 1 0 38976 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_496
timestamp 1621261055
transform 1 0 40800 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_407
timestamp 1621261055
transform 1 0 40224 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_411
timestamp 1621261055
transform 1 0 40608 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_414
timestamp 1621261055
transform 1 0 40896 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_402
timestamp 1621261055
transform 1 0 39744 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_410
timestamp 1621261055
transform 1 0 40512 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_418
timestamp 1621261055
transform 1 0 41280 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_426
timestamp 1621261055
transform 1 0 42048 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_422
timestamp 1621261055
transform 1 0 41664 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_436
timestamp 1621261055
transform 1 0 43008 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_31_432
timestamp 1621261055
transform 1 0 42624 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_430
timestamp 1621261055
transform 1 0 42432 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_435
timestamp 1621261055
transform 1 0 42912 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_430
timestamp 1621261055
transform 1 0 42432 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _186_
timestamp 1621261055
transform 1 0 42720 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _061_
timestamp 1621261055
transform 1 0 42624 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_441
timestamp 1621261055
transform 1 0 43488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_507
timestamp 1621261055
transform 1 0 43392 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_443
timestamp 1621261055
transform 1 0 43680 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_451
timestamp 1621261055
transform 1 0 44448 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_459
timestamp 1621261055
transform 1 0 45216 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_449
timestamp 1621261055
transform 1 0 44256 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_457
timestamp 1621261055
transform 1 0 45024 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_497
timestamp 1621261055
transform 1 0 46080 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_30_467
timestamp 1621261055
transform 1 0 45984 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_469
timestamp 1621261055
transform 1 0 46176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_477
timestamp 1621261055
transform 1 0 46944 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_465
timestamp 1621261055
transform 1 0 45792 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_473
timestamp 1621261055
transform 1 0 46560 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_481
timestamp 1621261055
transform 1 0 47328 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_508
timestamp 1621261055
transform 1 0 48672 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_485
timestamp 1621261055
transform 1 0 47712 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_493
timestamp 1621261055
transform 1 0 48480 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_501
timestamp 1621261055
transform 1 0 49248 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_489
timestamp 1621261055
transform 1 0 48096 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_493
timestamp 1621261055
transform 1 0 48480 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_496
timestamp 1621261055
transform 1 0 48768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_504
timestamp 1621261055
transform 1 0 49536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_498
timestamp 1621261055
transform 1 0 51360 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_509
timestamp 1621261055
transform 1 0 50016 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_517
timestamp 1621261055
transform 1 0 50784 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_521
timestamp 1621261055
transform 1 0 51168 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_524
timestamp 1621261055
transform 1 0 51456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_512
timestamp 1621261055
transform 1 0 50304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_520
timestamp 1621261055
transform 1 0 51072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_532
timestamp 1621261055
transform 1 0 52224 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_540
timestamp 1621261055
transform 1 0 52992 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_528
timestamp 1621261055
transform 1 0 51840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_536
timestamp 1621261055
transform 1 0 52608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_544
timestamp 1621261055
transform 1 0 53376 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_509
timestamp 1621261055
transform 1 0 53952 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_548
timestamp 1621261055
transform 1 0 53760 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_556
timestamp 1621261055
transform 1 0 54528 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_564
timestamp 1621261055
transform 1 0 55296 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_548
timestamp 1621261055
transform 1 0 53760 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_551
timestamp 1621261055
transform 1 0 54048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_559
timestamp 1621261055
transform 1 0 54816 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_567
timestamp 1621261055
transform 1 0 55584 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_499
timestamp 1621261055
transform 1 0 56640 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_572
timestamp 1621261055
transform 1 0 56064 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_576
timestamp 1621261055
transform 1 0 56448 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_579
timestamp 1621261055
transform 1 0 56736 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_587
timestamp 1621261055
transform 1 0 57504 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_575
timestamp 1621261055
transform 1 0 56352 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_583
timestamp 1621261055
transform 1 0 57120 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_61
timestamp 1621261055
transform -1 0 58848 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_63
timestamp 1621261055
transform -1 0 58848 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_595
timestamp 1621261055
transform 1 0 58272 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_591
timestamp 1621261055
transform 1 0 57888 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_595
timestamp 1621261055
transform 1 0 58272 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_64
timestamp 1621261055
transform 1 0 1152 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_32_4
timestamp 1621261055
transform 1 0 1536 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_12
timestamp 1621261055
transform 1 0 2304 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_20
timestamp 1621261055
transform 1 0 3072 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_510
timestamp 1621261055
transform 1 0 3840 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_29
timestamp 1621261055
transform 1 0 3936 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_37
timestamp 1621261055
transform 1 0 4704 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_45
timestamp 1621261055
transform 1 0 5472 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_53
timestamp 1621261055
transform 1 0 6240 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_61
timestamp 1621261055
transform 1 0 7008 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_511
timestamp 1621261055
transform 1 0 9120 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_69
timestamp 1621261055
transform 1 0 7776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_77
timestamp 1621261055
transform 1 0 8544 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_81
timestamp 1621261055
transform 1 0 8928 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_84
timestamp 1621261055
transform 1 0 9216 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_92
timestamp 1621261055
transform 1 0 9984 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_100
timestamp 1621261055
transform 1 0 10752 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_104
timestamp 1621261055
transform 1 0 11136 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _178_
timestamp 1621261055
transform 1 0 11424 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_32_106
timestamp 1621261055
transform 1 0 11328 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_110
timestamp 1621261055
transform 1 0 11712 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_118
timestamp 1621261055
transform 1 0 12480 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_126
timestamp 1621261055
transform 1 0 13248 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_512
timestamp 1621261055
transform 1 0 14400 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_134
timestamp 1621261055
transform 1 0 14016 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_32_139
timestamp 1621261055
transform 1 0 14496 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_147
timestamp 1621261055
transform 1 0 15264 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_155
timestamp 1621261055
transform 1 0 16032 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_163
timestamp 1621261055
transform 1 0 16800 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_171
timestamp 1621261055
transform 1 0 17568 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_179
timestamp 1621261055
transform 1 0 18336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_187
timestamp 1621261055
transform 1 0 19104 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_513
timestamp 1621261055
transform 1 0 19680 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_191
timestamp 1621261055
transform 1 0 19488 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_194
timestamp 1621261055
transform 1 0 19776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_202
timestamp 1621261055
transform 1 0 20544 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_210
timestamp 1621261055
transform 1 0 21312 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _099_
timestamp 1621261055
transform 1 0 22656 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_32_218
timestamp 1621261055
transform 1 0 22080 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_222
timestamp 1621261055
transform 1 0 22464 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_227
timestamp 1621261055
transform 1 0 22944 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_514
timestamp 1621261055
transform 1 0 24960 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_235
timestamp 1621261055
transform 1 0 23712 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_243
timestamp 1621261055
transform 1 0 24480 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_32_247
timestamp 1621261055
transform 1 0 24864 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_249
timestamp 1621261055
transform 1 0 25056 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_257
timestamp 1621261055
transform 1 0 25824 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_265
timestamp 1621261055
transform 1 0 26592 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_273
timestamp 1621261055
transform 1 0 27360 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_281
timestamp 1621261055
transform 1 0 28128 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_289
timestamp 1621261055
transform 1 0 28896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_515
timestamp 1621261055
transform 1 0 30240 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_297
timestamp 1621261055
transform 1 0 29664 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_301
timestamp 1621261055
transform 1 0 30048 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_304
timestamp 1621261055
transform 1 0 30336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_312
timestamp 1621261055
transform 1 0 31104 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_320
timestamp 1621261055
transform 1 0 31872 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_328
timestamp 1621261055
transform 1 0 32640 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_336
timestamp 1621261055
transform 1 0 33408 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_344
timestamp 1621261055
transform 1 0 34176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_352
timestamp 1621261055
transform 1 0 34944 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_356
timestamp 1621261055
transform 1 0 35328 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_516
timestamp 1621261055
transform 1 0 35520 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_359
timestamp 1621261055
transform 1 0 35616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_367
timestamp 1621261055
transform 1 0 36384 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_375
timestamp 1621261055
transform 1 0 37152 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_383
timestamp 1621261055
transform 1 0 37920 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_391
timestamp 1621261055
transform 1 0 38688 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_399
timestamp 1621261055
transform 1 0 39456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_517
timestamp 1621261055
transform 1 0 40800 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_407
timestamp 1621261055
transform 1 0 40224 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_411
timestamp 1621261055
transform 1 0 40608 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_414
timestamp 1621261055
transform 1 0 40896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_422
timestamp 1621261055
transform 1 0 41664 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_430
timestamp 1621261055
transform 1 0 42432 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_438
timestamp 1621261055
transform 1 0 43200 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_446
timestamp 1621261055
transform 1 0 43968 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_454
timestamp 1621261055
transform 1 0 44736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_462
timestamp 1621261055
transform 1 0 45504 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_518
timestamp 1621261055
transform 1 0 46080 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_466
timestamp 1621261055
transform 1 0 45888 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_469
timestamp 1621261055
transform 1 0 46176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_477
timestamp 1621261055
transform 1 0 46944 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_485
timestamp 1621261055
transform 1 0 47712 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_493
timestamp 1621261055
transform 1 0 48480 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_501
timestamp 1621261055
transform 1 0 49248 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_519
timestamp 1621261055
transform 1 0 51360 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_509
timestamp 1621261055
transform 1 0 50016 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_517
timestamp 1621261055
transform 1 0 50784 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_521
timestamp 1621261055
transform 1 0 51168 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_524
timestamp 1621261055
transform 1 0 51456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_532
timestamp 1621261055
transform 1 0 52224 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_540
timestamp 1621261055
transform 1 0 52992 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_548
timestamp 1621261055
transform 1 0 53760 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_556
timestamp 1621261055
transform 1 0 54528 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_564
timestamp 1621261055
transform 1 0 55296 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_520
timestamp 1621261055
transform 1 0 56640 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_572
timestamp 1621261055
transform 1 0 56064 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_576
timestamp 1621261055
transform 1 0 56448 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_579
timestamp 1621261055
transform 1 0 56736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_587
timestamp 1621261055
transform 1 0 57504 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_65
timestamp 1621261055
transform -1 0 58848 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_595
timestamp 1621261055
transform 1 0 58272 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_66
timestamp 1621261055
transform 1 0 1152 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_4
timestamp 1621261055
transform 1 0 1536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_12
timestamp 1621261055
transform 1 0 2304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_20
timestamp 1621261055
transform 1 0 3072 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_28
timestamp 1621261055
transform 1 0 3840 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_36
timestamp 1621261055
transform 1 0 4608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_521
timestamp 1621261055
transform 1 0 6432 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_44
timestamp 1621261055
transform 1 0 5376 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_52
timestamp 1621261055
transform 1 0 6144 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_54
timestamp 1621261055
transform 1 0 6336 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_56
timestamp 1621261055
transform 1 0 6528 0 1 24642
box -38 -49 806 715
use OAI22X1  OAI22X1
timestamp 1624074425
transform 1 0 7680 0 1 24642
box 0 -48 1440 714
use sky130_fd_sc_ls__decap_4  FILLER_33_64
timestamp 1621261055
transform 1 0 7296 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_83
timestamp 1621261055
transform 1 0 9120 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_91
timestamp 1621261055
transform 1 0 9888 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_99
timestamp 1621261055
transform 1 0 10656 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_522
timestamp 1621261055
transform 1 0 11712 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_107
timestamp 1621261055
transform 1 0 11424 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_109
timestamp 1621261055
transform 1 0 11616 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_111
timestamp 1621261055
transform 1 0 11808 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_119
timestamp 1621261055
transform 1 0 12576 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _145_
timestamp 1621261055
transform 1 0 14400 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_33_127
timestamp 1621261055
transform 1 0 13344 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_135
timestamp 1621261055
transform 1 0 14112 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_137
timestamp 1621261055
transform 1 0 14304 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_141
timestamp 1621261055
transform 1 0 14688 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_523
timestamp 1621261055
transform 1 0 16992 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_149
timestamp 1621261055
transform 1 0 15456 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_157
timestamp 1621261055
transform 1 0 16224 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_166
timestamp 1621261055
transform 1 0 17088 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_174
timestamp 1621261055
transform 1 0 17856 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_182
timestamp 1621261055
transform 1 0 18624 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_190
timestamp 1621261055
transform 1 0 19392 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_198
timestamp 1621261055
transform 1 0 20160 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_206
timestamp 1621261055
transform 1 0 20928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_524
timestamp 1621261055
transform 1 0 22272 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_214
timestamp 1621261055
transform 1 0 21696 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_218
timestamp 1621261055
transform 1 0 22080 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_221
timestamp 1621261055
transform 1 0 22368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_229
timestamp 1621261055
transform 1 0 23136 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_237
timestamp 1621261055
transform 1 0 23904 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_245
timestamp 1621261055
transform 1 0 24672 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_253
timestamp 1621261055
transform 1 0 25440 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_261
timestamp 1621261055
transform 1 0 26208 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_269
timestamp 1621261055
transform 1 0 26976 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_273
timestamp 1621261055
transform 1 0 27360 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_525
timestamp 1621261055
transform 1 0 27552 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_276
timestamp 1621261055
transform 1 0 27648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_284
timestamp 1621261055
transform 1 0 28416 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_292
timestamp 1621261055
transform 1 0 29184 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_300
timestamp 1621261055
transform 1 0 29952 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_308
timestamp 1621261055
transform 1 0 30720 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_526
timestamp 1621261055
transform 1 0 32832 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_316
timestamp 1621261055
transform 1 0 31488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_324
timestamp 1621261055
transform 1 0 32256 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_328
timestamp 1621261055
transform 1 0 32640 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_331
timestamp 1621261055
transform 1 0 32928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_339
timestamp 1621261055
transform 1 0 33696 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_347
timestamp 1621261055
transform 1 0 34464 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_355
timestamp 1621261055
transform 1 0 35232 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_363
timestamp 1621261055
transform 1 0 36000 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_371
timestamp 1621261055
transform 1 0 36768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_527
timestamp 1621261055
transform 1 0 38112 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_379
timestamp 1621261055
transform 1 0 37536 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_383
timestamp 1621261055
transform 1 0 37920 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_386
timestamp 1621261055
transform 1 0 38208 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_394
timestamp 1621261055
transform 1 0 38976 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_402
timestamp 1621261055
transform 1 0 39744 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_410
timestamp 1621261055
transform 1 0 40512 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_418
timestamp 1621261055
transform 1 0 41280 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_528
timestamp 1621261055
transform 1 0 43392 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_426
timestamp 1621261055
transform 1 0 42048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_434
timestamp 1621261055
transform 1 0 42816 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_438
timestamp 1621261055
transform 1 0 43200 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_441
timestamp 1621261055
transform 1 0 43488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_449
timestamp 1621261055
transform 1 0 44256 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_457
timestamp 1621261055
transform 1 0 45024 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_465
timestamp 1621261055
transform 1 0 45792 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_473
timestamp 1621261055
transform 1 0 46560 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_481
timestamp 1621261055
transform 1 0 47328 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_529
timestamp 1621261055
transform 1 0 48672 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_489
timestamp 1621261055
transform 1 0 48096 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_493
timestamp 1621261055
transform 1 0 48480 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_496
timestamp 1621261055
transform 1 0 48768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_33_504
timestamp 1621261055
transform 1 0 49536 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _123_
timestamp 1621261055
transform 1 0 49632 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_33_508
timestamp 1621261055
transform 1 0 49920 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_516
timestamp 1621261055
transform 1 0 50688 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_524
timestamp 1621261055
transform 1 0 51456 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _131_
timestamp 1621261055
transform 1 0 52320 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_33_532
timestamp 1621261055
transform 1 0 52224 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_536
timestamp 1621261055
transform 1 0 52608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_544
timestamp 1621261055
transform 1 0 53376 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_530
timestamp 1621261055
transform 1 0 53952 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_548
timestamp 1621261055
transform 1 0 53760 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_551
timestamp 1621261055
transform 1 0 54048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_559
timestamp 1621261055
transform 1 0 54816 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_567
timestamp 1621261055
transform 1 0 55584 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_575
timestamp 1621261055
transform 1 0 56352 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_583
timestamp 1621261055
transform 1 0 57120 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_67
timestamp 1621261055
transform -1 0 58848 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_33_591
timestamp 1621261055
transform 1 0 57888 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_595
timestamp 1621261055
transform 1 0 58272 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_68
timestamp 1621261055
transform 1 0 1152 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_4
timestamp 1621261055
transform 1 0 1536 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_12
timestamp 1621261055
transform 1 0 2304 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_20
timestamp 1621261055
transform 1 0 3072 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _194_
timestamp 1621261055
transform 1 0 4320 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_531
timestamp 1621261055
transform 1 0 3840 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_29
timestamp 1621261055
transform 1 0 3936 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_36
timestamp 1621261055
transform 1 0 4608 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _217_
timestamp 1621261055
transform 1 0 7104 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_37
timestamp 1621261055
transform 1 0 6912 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_44
timestamp 1621261055
transform 1 0 5376 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_52
timestamp 1621261055
transform 1 0 6144 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_532
timestamp 1621261055
transform 1 0 9120 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_65
timestamp 1621261055
transform 1 0 7392 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_73
timestamp 1621261055
transform 1 0 8160 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_81
timestamp 1621261055
transform 1 0 8928 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_84
timestamp 1621261055
transform 1 0 9216 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_92
timestamp 1621261055
transform 1 0 9984 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_100
timestamp 1621261055
transform 1 0 10752 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_108
timestamp 1621261055
transform 1 0 11520 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_116
timestamp 1621261055
transform 1 0 12288 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_124
timestamp 1621261055
transform 1 0 13056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_533
timestamp 1621261055
transform 1 0 14400 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_132
timestamp 1621261055
transform 1 0 13824 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_136
timestamp 1621261055
transform 1 0 14208 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_139
timestamp 1621261055
transform 1 0 14496 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_147
timestamp 1621261055
transform 1 0 15264 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_155
timestamp 1621261055
transform 1 0 16032 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_163
timestamp 1621261055
transform 1 0 16800 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_171
timestamp 1621261055
transform 1 0 17568 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_179
timestamp 1621261055
transform 1 0 18336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_187
timestamp 1621261055
transform 1 0 19104 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _050_
timestamp 1621261055
transform 1 0 21216 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_534
timestamp 1621261055
transform 1 0 19680 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_63
timestamp 1621261055
transform 1 0 21024 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_191
timestamp 1621261055
transform 1 0 19488 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_194
timestamp 1621261055
transform 1 0 19776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_202
timestamp 1621261055
transform 1 0 20544 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_34_206
timestamp 1621261055
transform 1 0 20928 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_212
timestamp 1621261055
transform 1 0 21504 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_220
timestamp 1621261055
transform 1 0 22272 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_228
timestamp 1621261055
transform 1 0 23040 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_535
timestamp 1621261055
transform 1 0 24960 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_236
timestamp 1621261055
transform 1 0 23808 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_244
timestamp 1621261055
transform 1 0 24576 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_249
timestamp 1621261055
transform 1 0 25056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_257
timestamp 1621261055
transform 1 0 25824 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_265
timestamp 1621261055
transform 1 0 26592 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_273
timestamp 1621261055
transform 1 0 27360 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_281
timestamp 1621261055
transform 1 0 28128 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_289
timestamp 1621261055
transform 1 0 28896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_536
timestamp 1621261055
transform 1 0 30240 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_297
timestamp 1621261055
transform 1 0 29664 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_301
timestamp 1621261055
transform 1 0 30048 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_304
timestamp 1621261055
transform 1 0 30336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_312
timestamp 1621261055
transform 1 0 31104 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_320
timestamp 1621261055
transform 1 0 31872 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_328
timestamp 1621261055
transform 1 0 32640 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_336
timestamp 1621261055
transform 1 0 33408 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_344
timestamp 1621261055
transform 1 0 34176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_352
timestamp 1621261055
transform 1 0 34944 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_356
timestamp 1621261055
transform 1 0 35328 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_537
timestamp 1621261055
transform 1 0 35520 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_359
timestamp 1621261055
transform 1 0 35616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_367
timestamp 1621261055
transform 1 0 36384 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_375
timestamp 1621261055
transform 1 0 37152 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_383
timestamp 1621261055
transform 1 0 37920 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_391
timestamp 1621261055
transform 1 0 38688 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_399
timestamp 1621261055
transform 1 0 39456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_538
timestamp 1621261055
transform 1 0 40800 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_407
timestamp 1621261055
transform 1 0 40224 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_411
timestamp 1621261055
transform 1 0 40608 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_414
timestamp 1621261055
transform 1 0 40896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_422
timestamp 1621261055
transform 1 0 41664 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_430
timestamp 1621261055
transform 1 0 42432 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_438
timestamp 1621261055
transform 1 0 43200 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_446
timestamp 1621261055
transform 1 0 43968 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_454
timestamp 1621261055
transform 1 0 44736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_462
timestamp 1621261055
transform 1 0 45504 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_539
timestamp 1621261055
transform 1 0 46080 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_466
timestamp 1621261055
transform 1 0 45888 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_469
timestamp 1621261055
transform 1 0 46176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_477
timestamp 1621261055
transform 1 0 46944 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_485
timestamp 1621261055
transform 1 0 47712 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_493
timestamp 1621261055
transform 1 0 48480 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_501
timestamp 1621261055
transform 1 0 49248 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_540
timestamp 1621261055
transform 1 0 51360 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_509
timestamp 1621261055
transform 1 0 50016 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_517
timestamp 1621261055
transform 1 0 50784 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_521
timestamp 1621261055
transform 1 0 51168 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_524
timestamp 1621261055
transform 1 0 51456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_532
timestamp 1621261055
transform 1 0 52224 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_540
timestamp 1621261055
transform 1 0 52992 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _055_
timestamp 1621261055
transform -1 0 55776 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_75
timestamp 1621261055
transform -1 0 55488 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_548
timestamp 1621261055
transform 1 0 53760 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_556
timestamp 1621261055
transform 1 0 54528 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_541
timestamp 1621261055
transform 1 0 56640 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_569
timestamp 1621261055
transform 1 0 55776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_34_577
timestamp 1621261055
transform 1 0 56544 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_579
timestamp 1621261055
transform 1 0 56736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_587
timestamp 1621261055
transform 1 0 57504 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_69
timestamp 1621261055
transform -1 0 58848 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_595
timestamp 1621261055
transform 1 0 58272 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_70
timestamp 1621261055
transform 1 0 1152 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_4
timestamp 1621261055
transform 1 0 1536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_12
timestamp 1621261055
transform 1 0 2304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_20
timestamp 1621261055
transform 1 0 3072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_28
timestamp 1621261055
transform 1 0 3840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_36
timestamp 1621261055
transform 1 0 4608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_542
timestamp 1621261055
transform 1 0 6432 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_44
timestamp 1621261055
transform 1 0 5376 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_52
timestamp 1621261055
transform 1 0 6144 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_35_54
timestamp 1621261055
transform 1 0 6336 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_56
timestamp 1621261055
transform 1 0 6528 0 1 25974
box -38 -49 806 715
use OR2X1  OR2X1
timestamp 1624074425
transform 1 0 7680 0 1 25974
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_4  FILLER_35_64
timestamp 1621261055
transform 1 0 7296 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_80
timestamp 1621261055
transform 1 0 8832 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_88
timestamp 1621261055
transform 1 0 9600 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_96
timestamp 1621261055
transform 1 0 10368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_104
timestamp 1621261055
transform 1 0 11136 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_543
timestamp 1621261055
transform 1 0 11712 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_108
timestamp 1621261055
transform 1 0 11520 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_111
timestamp 1621261055
transform 1 0 11808 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_119
timestamp 1621261055
transform 1 0 12576 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_127
timestamp 1621261055
transform 1 0 13344 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_135
timestamp 1621261055
transform 1 0 14112 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_143
timestamp 1621261055
transform 1 0 14880 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_544
timestamp 1621261055
transform 1 0 16992 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_151
timestamp 1621261055
transform 1 0 15648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_159
timestamp 1621261055
transform 1 0 16416 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_163
timestamp 1621261055
transform 1 0 16800 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_166
timestamp 1621261055
transform 1 0 17088 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_174
timestamp 1621261055
transform 1 0 17856 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_182
timestamp 1621261055
transform 1 0 18624 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_190
timestamp 1621261055
transform 1 0 19392 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_198
timestamp 1621261055
transform 1 0 20160 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_206
timestamp 1621261055
transform 1 0 20928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_545
timestamp 1621261055
transform 1 0 22272 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_214
timestamp 1621261055
transform 1 0 21696 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_218
timestamp 1621261055
transform 1 0 22080 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_221
timestamp 1621261055
transform 1 0 22368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_229
timestamp 1621261055
transform 1 0 23136 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _190_
timestamp 1621261055
transform 1 0 24000 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_35_237
timestamp 1621261055
transform 1 0 23904 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_241
timestamp 1621261055
transform 1 0 24288 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_249
timestamp 1621261055
transform 1 0 25056 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_257
timestamp 1621261055
transform 1 0 25824 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_265
timestamp 1621261055
transform 1 0 26592 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_273
timestamp 1621261055
transform 1 0 27360 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_546
timestamp 1621261055
transform 1 0 27552 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_276
timestamp 1621261055
transform 1 0 27648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_284
timestamp 1621261055
transform 1 0 28416 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_292
timestamp 1621261055
transform 1 0 29184 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_300
timestamp 1621261055
transform 1 0 29952 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_308
timestamp 1621261055
transform 1 0 30720 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_547
timestamp 1621261055
transform 1 0 32832 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_316
timestamp 1621261055
transform 1 0 31488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_324
timestamp 1621261055
transform 1 0 32256 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_328
timestamp 1621261055
transform 1 0 32640 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_331
timestamp 1621261055
transform 1 0 32928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_339
timestamp 1621261055
transform 1 0 33696 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_347
timestamp 1621261055
transform 1 0 34464 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_355
timestamp 1621261055
transform 1 0 35232 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_363
timestamp 1621261055
transform 1 0 36000 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_371
timestamp 1621261055
transform 1 0 36768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _116_
timestamp 1621261055
transform 1 0 38784 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_548
timestamp 1621261055
transform 1 0 38112 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_379
timestamp 1621261055
transform 1 0 37536 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_383
timestamp 1621261055
transform 1 0 37920 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_35_386
timestamp 1621261055
transform 1 0 38208 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_390
timestamp 1621261055
transform 1 0 38592 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_395
timestamp 1621261055
transform 1 0 39072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_403
timestamp 1621261055
transform 1 0 39840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_411
timestamp 1621261055
transform 1 0 40608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_419
timestamp 1621261055
transform 1 0 41376 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_549
timestamp 1621261055
transform 1 0 43392 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_427
timestamp 1621261055
transform 1 0 42144 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_435
timestamp 1621261055
transform 1 0 42912 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_35_439
timestamp 1621261055
transform 1 0 43296 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_441
timestamp 1621261055
transform 1 0 43488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_449
timestamp 1621261055
transform 1 0 44256 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_457
timestamp 1621261055
transform 1 0 45024 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_465
timestamp 1621261055
transform 1 0 45792 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_473
timestamp 1621261055
transform 1 0 46560 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_481
timestamp 1621261055
transform 1 0 47328 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_550
timestamp 1621261055
transform 1 0 48672 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_489
timestamp 1621261055
transform 1 0 48096 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_493
timestamp 1621261055
transform 1 0 48480 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_496
timestamp 1621261055
transform 1 0 48768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_504
timestamp 1621261055
transform 1 0 49536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_512
timestamp 1621261055
transform 1 0 50304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_520
timestamp 1621261055
transform 1 0 51072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_528
timestamp 1621261055
transform 1 0 51840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_536
timestamp 1621261055
transform 1 0 52608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_544
timestamp 1621261055
transform 1 0 53376 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_551
timestamp 1621261055
transform 1 0 53952 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_548
timestamp 1621261055
transform 1 0 53760 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_551
timestamp 1621261055
transform 1 0 54048 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_559
timestamp 1621261055
transform 1 0 54816 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_567
timestamp 1621261055
transform 1 0 55584 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _066_
timestamp 1621261055
transform 1 0 57120 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_35_575
timestamp 1621261055
transform 1 0 56352 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_586
timestamp 1621261055
transform 1 0 57408 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_71
timestamp 1621261055
transform -1 0 58848 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_594
timestamp 1621261055
transform 1 0 58176 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_35_596
timestamp 1621261055
transform 1 0 58368 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_72
timestamp 1621261055
transform 1 0 1152 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_4
timestamp 1621261055
transform 1 0 1536 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_12
timestamp 1621261055
transform 1 0 2304 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_20
timestamp 1621261055
transform 1 0 3072 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_552
timestamp 1621261055
transform 1 0 3840 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_29
timestamp 1621261055
transform 1 0 3936 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_37
timestamp 1621261055
transform 1 0 4704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_45
timestamp 1621261055
transform 1 0 5472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_53
timestamp 1621261055
transform 1 0 6240 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_61
timestamp 1621261055
transform 1 0 7008 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_553
timestamp 1621261055
transform 1 0 9120 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_69
timestamp 1621261055
transform 1 0 7776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_77
timestamp 1621261055
transform 1 0 8544 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_81
timestamp 1621261055
transform 1 0 8928 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_84
timestamp 1621261055
transform 1 0 9216 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_92
timestamp 1621261055
transform 1 0 9984 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_100
timestamp 1621261055
transform 1 0 10752 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_108
timestamp 1621261055
transform 1 0 11520 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_116
timestamp 1621261055
transform 1 0 12288 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_124
timestamp 1621261055
transform 1 0 13056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _002_
timestamp 1621261055
transform -1 0 15168 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_554
timestamp 1621261055
transform 1 0 14400 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_6
timestamp 1621261055
transform -1 0 14880 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_36_132
timestamp 1621261055
transform 1 0 13824 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_136
timestamp 1621261055
transform 1 0 14208 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_139
timestamp 1621261055
transform 1 0 14496 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_146
timestamp 1621261055
transform 1 0 15168 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_154
timestamp 1621261055
transform 1 0 15936 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_162
timestamp 1621261055
transform 1 0 16704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_170
timestamp 1621261055
transform 1 0 17472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_178
timestamp 1621261055
transform 1 0 18240 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_186
timestamp 1621261055
transform 1 0 19008 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_555
timestamp 1621261055
transform 1 0 19680 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_190
timestamp 1621261055
transform 1 0 19392 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_36_192
timestamp 1621261055
transform 1 0 19584 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_194
timestamp 1621261055
transform 1 0 19776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_202
timestamp 1621261055
transform 1 0 20544 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_210
timestamp 1621261055
transform 1 0 21312 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_218
timestamp 1621261055
transform 1 0 22080 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_226
timestamp 1621261055
transform 1 0 22848 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_556
timestamp 1621261055
transform 1 0 24960 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_234
timestamp 1621261055
transform 1 0 23616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_242
timestamp 1621261055
transform 1 0 24384 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_246
timestamp 1621261055
transform 1 0 24768 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_249
timestamp 1621261055
transform 1 0 25056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_257
timestamp 1621261055
transform 1 0 25824 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_265
timestamp 1621261055
transform 1 0 26592 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_273
timestamp 1621261055
transform 1 0 27360 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _168_
timestamp 1621261055
transform 1 0 28416 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_281
timestamp 1621261055
transform 1 0 28128 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_36_283
timestamp 1621261055
transform 1 0 28320 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_287
timestamp 1621261055
transform 1 0 28704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_557
timestamp 1621261055
transform 1 0 30240 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_295
timestamp 1621261055
transform 1 0 29472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_304
timestamp 1621261055
transform 1 0 30336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_312
timestamp 1621261055
transform 1 0 31104 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_320
timestamp 1621261055
transform 1 0 31872 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_328
timestamp 1621261055
transform 1 0 32640 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_336
timestamp 1621261055
transform 1 0 33408 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_344
timestamp 1621261055
transform 1 0 34176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_352
timestamp 1621261055
transform 1 0 34944 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_356
timestamp 1621261055
transform 1 0 35328 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_558
timestamp 1621261055
transform 1 0 35520 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_359
timestamp 1621261055
transform 1 0 35616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_367
timestamp 1621261055
transform 1 0 36384 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_375
timestamp 1621261055
transform 1 0 37152 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_383
timestamp 1621261055
transform 1 0 37920 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_391
timestamp 1621261055
transform 1 0 38688 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_399
timestamp 1621261055
transform 1 0 39456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_559
timestamp 1621261055
transform 1 0 40800 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_407
timestamp 1621261055
transform 1 0 40224 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_411
timestamp 1621261055
transform 1 0 40608 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_414
timestamp 1621261055
transform 1 0 40896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_422
timestamp 1621261055
transform 1 0 41664 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_430
timestamp 1621261055
transform 1 0 42432 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_438
timestamp 1621261055
transform 1 0 43200 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_446
timestamp 1621261055
transform 1 0 43968 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_454
timestamp 1621261055
transform 1 0 44736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_462
timestamp 1621261055
transform 1 0 45504 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _038_
timestamp 1621261055
transform -1 0 47712 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_560
timestamp 1621261055
transform 1 0 46080 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_87
timestamp 1621261055
transform -1 0 47424 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_466
timestamp 1621261055
transform 1 0 45888 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_469
timestamp 1621261055
transform 1 0 46176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_477
timestamp 1621261055
transform 1 0 46944 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_36_479
timestamp 1621261055
transform 1 0 47136 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_485
timestamp 1621261055
transform 1 0 47712 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_493
timestamp 1621261055
transform 1 0 48480 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_501
timestamp 1621261055
transform 1 0 49248 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_561
timestamp 1621261055
transform 1 0 51360 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_509
timestamp 1621261055
transform 1 0 50016 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_517
timestamp 1621261055
transform 1 0 50784 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_521
timestamp 1621261055
transform 1 0 51168 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_524
timestamp 1621261055
transform 1 0 51456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_532
timestamp 1621261055
transform 1 0 52224 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_540
timestamp 1621261055
transform 1 0 52992 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_548
timestamp 1621261055
transform 1 0 53760 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_556
timestamp 1621261055
transform 1 0 54528 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_564
timestamp 1621261055
transform 1 0 55296 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_562
timestamp 1621261055
transform 1 0 56640 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_572
timestamp 1621261055
transform 1 0 56064 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_576
timestamp 1621261055
transform 1 0 56448 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_579
timestamp 1621261055
transform 1 0 56736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_587
timestamp 1621261055
transform 1 0 57504 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_73
timestamp 1621261055
transform -1 0 58848 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_595
timestamp 1621261055
transform 1 0 58272 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_74
timestamp 1621261055
transform 1 0 1152 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_4
timestamp 1621261055
transform 1 0 1536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_12
timestamp 1621261055
transform 1 0 2304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_20
timestamp 1621261055
transform 1 0 3072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_28
timestamp 1621261055
transform 1 0 3840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_36
timestamp 1621261055
transform 1 0 4608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_563
timestamp 1621261055
transform 1 0 6432 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_44
timestamp 1621261055
transform 1 0 5376 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_52
timestamp 1621261055
transform 1 0 6144 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_54
timestamp 1621261055
transform 1 0 6336 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_56
timestamp 1621261055
transform 1 0 6528 0 1 27306
box -38 -49 806 715
use OR2X2  OR2X2
timestamp 1624074425
transform 1 0 7680 0 1 27306
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_4  FILLER_37_64
timestamp 1621261055
transform 1 0 7296 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_80
timestamp 1621261055
transform 1 0 8832 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_88
timestamp 1621261055
transform 1 0 9600 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_96
timestamp 1621261055
transform 1 0 10368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_104
timestamp 1621261055
transform 1 0 11136 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_564
timestamp 1621261055
transform 1 0 11712 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_108
timestamp 1621261055
transform 1 0 11520 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_111
timestamp 1621261055
transform 1 0 11808 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_119
timestamp 1621261055
transform 1 0 12576 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _198_
timestamp 1621261055
transform 1 0 14112 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_37_127
timestamp 1621261055
transform 1 0 13344 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_138
timestamp 1621261055
transform 1 0 14400 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_146
timestamp 1621261055
transform 1 0 15168 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_565
timestamp 1621261055
transform 1 0 16992 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_154
timestamp 1621261055
transform 1 0 15936 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_162
timestamp 1621261055
transform 1 0 16704 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_164
timestamp 1621261055
transform 1 0 16896 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_166
timestamp 1621261055
transform 1 0 17088 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_174
timestamp 1621261055
transform 1 0 17856 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_182
timestamp 1621261055
transform 1 0 18624 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_190
timestamp 1621261055
transform 1 0 19392 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_198
timestamp 1621261055
transform 1 0 20160 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_206
timestamp 1621261055
transform 1 0 20928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_566
timestamp 1621261055
transform 1 0 22272 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_214
timestamp 1621261055
transform 1 0 21696 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_218
timestamp 1621261055
transform 1 0 22080 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_221
timestamp 1621261055
transform 1 0 22368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_229
timestamp 1621261055
transform 1 0 23136 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_237
timestamp 1621261055
transform 1 0 23904 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_245
timestamp 1621261055
transform 1 0 24672 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_253
timestamp 1621261055
transform 1 0 25440 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_261
timestamp 1621261055
transform 1 0 26208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_269
timestamp 1621261055
transform 1 0 26976 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_273
timestamp 1621261055
transform 1 0 27360 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_567
timestamp 1621261055
transform 1 0 27552 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_276
timestamp 1621261055
transform 1 0 27648 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_284
timestamp 1621261055
transform 1 0 28416 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_292
timestamp 1621261055
transform 1 0 29184 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_300
timestamp 1621261055
transform 1 0 29952 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_308
timestamp 1621261055
transform 1 0 30720 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_568
timestamp 1621261055
transform 1 0 32832 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_316
timestamp 1621261055
transform 1 0 31488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_324
timestamp 1621261055
transform 1 0 32256 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_328
timestamp 1621261055
transform 1 0 32640 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_331
timestamp 1621261055
transform 1 0 32928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_339
timestamp 1621261055
transform 1 0 33696 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_347
timestamp 1621261055
transform 1 0 34464 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_355
timestamp 1621261055
transform 1 0 35232 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_363
timestamp 1621261055
transform 1 0 36000 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_371
timestamp 1621261055
transform 1 0 36768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_569
timestamp 1621261055
transform 1 0 38112 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_379
timestamp 1621261055
transform 1 0 37536 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_383
timestamp 1621261055
transform 1 0 37920 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_386
timestamp 1621261055
transform 1 0 38208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_394
timestamp 1621261055
transform 1 0 38976 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_402
timestamp 1621261055
transform 1 0 39744 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_410
timestamp 1621261055
transform 1 0 40512 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_418
timestamp 1621261055
transform 1 0 41280 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_570
timestamp 1621261055
transform 1 0 43392 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_426
timestamp 1621261055
transform 1 0 42048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_434
timestamp 1621261055
transform 1 0 42816 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_438
timestamp 1621261055
transform 1 0 43200 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_441
timestamp 1621261055
transform 1 0 43488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_449
timestamp 1621261055
transform 1 0 44256 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_457
timestamp 1621261055
transform 1 0 45024 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_465
timestamp 1621261055
transform 1 0 45792 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_473
timestamp 1621261055
transform 1 0 46560 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_481
timestamp 1621261055
transform 1 0 47328 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_571
timestamp 1621261055
transform 1 0 48672 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_489
timestamp 1621261055
transform 1 0 48096 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_493
timestamp 1621261055
transform 1 0 48480 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_496
timestamp 1621261055
transform 1 0 48768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_504
timestamp 1621261055
transform 1 0 49536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_512
timestamp 1621261055
transform 1 0 50304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_520
timestamp 1621261055
transform 1 0 51072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_528
timestamp 1621261055
transform 1 0 51840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_536
timestamp 1621261055
transform 1 0 52608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_544
timestamp 1621261055
transform 1 0 53376 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _046_
timestamp 1621261055
transform -1 0 55680 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_572
timestamp 1621261055
transform 1 0 53952 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_45
timestamp 1621261055
transform -1 0 55392 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_548
timestamp 1621261055
transform 1 0 53760 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_551
timestamp 1621261055
transform 1 0 54048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_559
timestamp 1621261055
transform 1 0 54816 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_568
timestamp 1621261055
transform 1 0 55680 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_576
timestamp 1621261055
transform 1 0 56448 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_584
timestamp 1621261055
transform 1 0 57216 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_75
timestamp 1621261055
transform -1 0 58848 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_37_592
timestamp 1621261055
transform 1 0 57984 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_37_596
timestamp 1621261055
transform 1 0 58368 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_76
timestamp 1621261055
transform 1 0 1152 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_78
timestamp 1621261055
transform 1 0 1152 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_4
timestamp 1621261055
transform 1 0 1536 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_12
timestamp 1621261055
transform 1 0 2304 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_20
timestamp 1621261055
transform 1 0 3072 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_4
timestamp 1621261055
transform 1 0 1536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_12
timestamp 1621261055
transform 1 0 2304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_20
timestamp 1621261055
transform 1 0 3072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_573
timestamp 1621261055
transform 1 0 3840 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_29
timestamp 1621261055
transform 1 0 3936 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_37
timestamp 1621261055
transform 1 0 4704 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_28
timestamp 1621261055
transform 1 0 3840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_36
timestamp 1621261055
transform 1 0 4608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_584
timestamp 1621261055
transform 1 0 6432 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_45
timestamp 1621261055
transform 1 0 5472 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_53
timestamp 1621261055
transform 1 0 6240 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_61
timestamp 1621261055
transform 1 0 7008 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_44
timestamp 1621261055
transform 1 0 5376 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_52
timestamp 1621261055
transform 1 0 6144 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_39_54
timestamp 1621261055
transform 1 0 6336 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_56
timestamp 1621261055
transform 1 0 6528 0 1 28638
box -38 -49 806 715
use XOR2X1  XOR2X1
timestamp 1624074425
transform 1 0 7680 0 1 28638
box 0 -48 2016 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_574
timestamp 1621261055
transform 1 0 9120 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_69
timestamp 1621261055
transform 1 0 7776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_77
timestamp 1621261055
transform 1 0 8544 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_81
timestamp 1621261055
transform 1 0 8928 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_84
timestamp 1621261055
transform 1 0 9216 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_64
timestamp 1621261055
transform 1 0 7296 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_92
timestamp 1621261055
transform 1 0 9984 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_100
timestamp 1621261055
transform 1 0 10752 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_89
timestamp 1621261055
transform 1 0 9696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_97
timestamp 1621261055
transform 1 0 10464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_105
timestamp 1621261055
transform 1 0 11232 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_585
timestamp 1621261055
transform 1 0 11712 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_108
timestamp 1621261055
transform 1 0 11520 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_116
timestamp 1621261055
transform 1 0 12288 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_124
timestamp 1621261055
transform 1 0 13056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_109
timestamp 1621261055
transform 1 0 11616 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_111
timestamp 1621261055
transform 1 0 11808 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_119
timestamp 1621261055
transform 1 0 12576 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_127
timestamp 1621261055
transform 1 0 13344 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_132
timestamp 1621261055
transform 1 0 13824 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_39_141
timestamp 1621261055
transform 1 0 14688 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_39_135
timestamp 1621261055
transform 1 0 14112 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_139
timestamp 1621261055
transform 1 0 14496 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_136
timestamp 1621261055
transform 1 0 14208 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_0
timestamp 1621261055
transform 1 0 14208 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_575
timestamp 1621261055
transform 1 0 14400 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _016_
timestamp 1621261055
transform 1 0 14400 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_38_147
timestamp 1621261055
transform 1 0 15264 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _161_
timestamp 1621261055
transform 1 0 15072 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_586
timestamp 1621261055
transform 1 0 16992 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_155
timestamp 1621261055
transform 1 0 16032 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_163
timestamp 1621261055
transform 1 0 16800 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_148
timestamp 1621261055
transform 1 0 15360 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_156
timestamp 1621261055
transform 1 0 16128 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_164
timestamp 1621261055
transform 1 0 16896 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_166
timestamp 1621261055
transform 1 0 17088 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_171
timestamp 1621261055
transform 1 0 17568 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_179
timestamp 1621261055
transform 1 0 18336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_187
timestamp 1621261055
transform 1 0 19104 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_174
timestamp 1621261055
transform 1 0 17856 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_182
timestamp 1621261055
transform 1 0 18624 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _092_
timestamp 1621261055
transform 1 0 20160 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_576
timestamp 1621261055
transform 1 0 19680 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_191
timestamp 1621261055
transform 1 0 19488 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_194
timestamp 1621261055
transform 1 0 19776 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_201
timestamp 1621261055
transform 1 0 20448 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_209
timestamp 1621261055
transform 1 0 21216 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_190
timestamp 1621261055
transform 1 0 19392 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_198
timestamp 1621261055
transform 1 0 20160 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_206
timestamp 1621261055
transform 1 0 20928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_587
timestamp 1621261055
transform 1 0 22272 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_217
timestamp 1621261055
transform 1 0 21984 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_225
timestamp 1621261055
transform 1 0 22752 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_214
timestamp 1621261055
transform 1 0 21696 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_218
timestamp 1621261055
transform 1 0 22080 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_221
timestamp 1621261055
transform 1 0 22368 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_229
timestamp 1621261055
transform 1 0 23136 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_577
timestamp 1621261055
transform 1 0 24960 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_233
timestamp 1621261055
transform 1 0 23520 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_241
timestamp 1621261055
transform 1 0 24288 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_245
timestamp 1621261055
transform 1 0 24672 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_38_247
timestamp 1621261055
transform 1 0 24864 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_249
timestamp 1621261055
transform 1 0 25056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_237
timestamp 1621261055
transform 1 0 23904 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_245
timestamp 1621261055
transform 1 0 24672 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_257
timestamp 1621261055
transform 1 0 25824 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_265
timestamp 1621261055
transform 1 0 26592 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_273
timestamp 1621261055
transform 1 0 27360 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_253
timestamp 1621261055
transform 1 0 25440 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_261
timestamp 1621261055
transform 1 0 26208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_269
timestamp 1621261055
transform 1 0 26976 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_273
timestamp 1621261055
transform 1 0 27360 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_588
timestamp 1621261055
transform 1 0 27552 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_281
timestamp 1621261055
transform 1 0 28128 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_289
timestamp 1621261055
transform 1 0 28896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_276
timestamp 1621261055
transform 1 0 27648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_284
timestamp 1621261055
transform 1 0 28416 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_292
timestamp 1621261055
transform 1 0 29184 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_578
timestamp 1621261055
transform 1 0 30240 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_297
timestamp 1621261055
transform 1 0 29664 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_301
timestamp 1621261055
transform 1 0 30048 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_304
timestamp 1621261055
transform 1 0 30336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_312
timestamp 1621261055
transform 1 0 31104 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_300
timestamp 1621261055
transform 1 0 29952 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_308
timestamp 1621261055
transform 1 0 30720 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_589
timestamp 1621261055
transform 1 0 32832 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_320
timestamp 1621261055
transform 1 0 31872 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_328
timestamp 1621261055
transform 1 0 32640 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_336
timestamp 1621261055
transform 1 0 33408 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_316
timestamp 1621261055
transform 1 0 31488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_324
timestamp 1621261055
transform 1 0 32256 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_328
timestamp 1621261055
transform 1 0 32640 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_331
timestamp 1621261055
transform 1 0 32928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_344
timestamp 1621261055
transform 1 0 34176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_352
timestamp 1621261055
transform 1 0 34944 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_356
timestamp 1621261055
transform 1 0 35328 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_339
timestamp 1621261055
transform 1 0 33696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_347
timestamp 1621261055
transform 1 0 34464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_355
timestamp 1621261055
transform 1 0 35232 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_579
timestamp 1621261055
transform 1 0 35520 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_359
timestamp 1621261055
transform 1 0 35616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_367
timestamp 1621261055
transform 1 0 36384 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_375
timestamp 1621261055
transform 1 0 37152 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_363
timestamp 1621261055
transform 1 0 36000 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_371
timestamp 1621261055
transform 1 0 36768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_386
timestamp 1621261055
transform 1 0 38208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_383
timestamp 1621261055
transform 1 0 37920 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_379
timestamp 1621261055
transform 1 0 37536 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_383
timestamp 1621261055
transform 1 0 37920 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_55
timestamp 1621261055
transform -1 0 38304 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_590
timestamp 1621261055
transform 1 0 38112 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_394
timestamp 1621261055
transform 1 0 38976 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_390
timestamp 1621261055
transform 1 0 38592 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _036_
timestamp 1621261055
transform -1 0 38592 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_38_398
timestamp 1621261055
transform 1 0 39360 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_402
timestamp 1621261055
transform 1 0 39744 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_406
timestamp 1621261055
transform 1 0 40128 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_410
timestamp 1621261055
transform 1 0 40512 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_414
timestamp 1621261055
transform 1 0 40896 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_38_412
timestamp 1621261055
transform 1 0 40704 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_410
timestamp 1621261055
transform 1 0 40512 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_580
timestamp 1621261055
transform 1 0 40800 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_418
timestamp 1621261055
transform 1 0 41280 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_38_420
timestamp 1621261055
transform 1 0 41472 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_418
timestamp 1621261055
transform 1 0 41280 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _087_
timestamp 1621261055
transform 1 0 41568 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_591
timestamp 1621261055
transform 1 0 43392 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_424
timestamp 1621261055
transform 1 0 41856 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_432
timestamp 1621261055
transform 1 0 42624 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_440
timestamp 1621261055
transform 1 0 43392 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_426
timestamp 1621261055
transform 1 0 42048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_434
timestamp 1621261055
transform 1 0 42816 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_438
timestamp 1621261055
transform 1 0 43200 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_441
timestamp 1621261055
transform 1 0 43488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _154_
timestamp 1621261055
transform 1 0 44544 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_38_448
timestamp 1621261055
transform 1 0 44160 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_456
timestamp 1621261055
transform 1 0 44928 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_449
timestamp 1621261055
transform 1 0 44256 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_39_451
timestamp 1621261055
transform 1 0 44448 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_455
timestamp 1621261055
transform 1 0 44832 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _125_
timestamp 1621261055
transform 1 0 46656 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_581
timestamp 1621261055
transform 1 0 46080 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_464
timestamp 1621261055
transform 1 0 45696 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_469
timestamp 1621261055
transform 1 0 46176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_477
timestamp 1621261055
transform 1 0 46944 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_463
timestamp 1621261055
transform 1 0 45600 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_471
timestamp 1621261055
transform 1 0 46368 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_39_473
timestamp 1621261055
transform 1 0 46560 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_477
timestamp 1621261055
transform 1 0 46944 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_592
timestamp 1621261055
transform 1 0 48672 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_485
timestamp 1621261055
transform 1 0 47712 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_493
timestamp 1621261055
transform 1 0 48480 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_501
timestamp 1621261055
transform 1 0 49248 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_485
timestamp 1621261055
transform 1 0 47712 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_493
timestamp 1621261055
transform 1 0 48480 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_496
timestamp 1621261055
transform 1 0 48768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_504
timestamp 1621261055
transform 1 0 49536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_582
timestamp 1621261055
transform 1 0 51360 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_509
timestamp 1621261055
transform 1 0 50016 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_517
timestamp 1621261055
transform 1 0 50784 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_521
timestamp 1621261055
transform 1 0 51168 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_524
timestamp 1621261055
transform 1 0 51456 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_512
timestamp 1621261055
transform 1 0 50304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_520
timestamp 1621261055
transform 1 0 51072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_532
timestamp 1621261055
transform 1 0 52224 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_540
timestamp 1621261055
transform 1 0 52992 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_528
timestamp 1621261055
transform 1 0 51840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_536
timestamp 1621261055
transform 1 0 52608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_544
timestamp 1621261055
transform 1 0 53376 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_593
timestamp 1621261055
transform 1 0 53952 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_548
timestamp 1621261055
transform 1 0 53760 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_556
timestamp 1621261055
transform 1 0 54528 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_564
timestamp 1621261055
transform 1 0 55296 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_548
timestamp 1621261055
transform 1 0 53760 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_551
timestamp 1621261055
transform 1 0 54048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_559
timestamp 1621261055
transform 1 0 54816 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_567
timestamp 1621261055
transform 1 0 55584 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _037_
timestamp 1621261055
transform -1 0 56160 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_583
timestamp 1621261055
transform 1 0 56640 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_85
timestamp 1621261055
transform -1 0 55872 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_572
timestamp 1621261055
transform 1 0 56064 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_576
timestamp 1621261055
transform 1 0 56448 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_579
timestamp 1621261055
transform 1 0 56736 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_587
timestamp 1621261055
transform 1 0 57504 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_573
timestamp 1621261055
transform 1 0 56160 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_581
timestamp 1621261055
transform 1 0 56928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_77
timestamp 1621261055
transform -1 0 58848 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_79
timestamp 1621261055
transform -1 0 58848 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_595
timestamp 1621261055
transform 1 0 58272 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_589
timestamp 1621261055
transform 1 0 57696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_80
timestamp 1621261055
transform 1 0 1152 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_40_4
timestamp 1621261055
transform 1 0 1536 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_12
timestamp 1621261055
transform 1 0 2304 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_20
timestamp 1621261055
transform 1 0 3072 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_594
timestamp 1621261055
transform 1 0 3840 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_29
timestamp 1621261055
transform 1 0 3936 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_37
timestamp 1621261055
transform 1 0 4704 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_45
timestamp 1621261055
transform 1 0 5472 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_53
timestamp 1621261055
transform 1 0 6240 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_61
timestamp 1621261055
transform 1 0 7008 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_595
timestamp 1621261055
transform 1 0 9120 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_69
timestamp 1621261055
transform 1 0 7776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_77
timestamp 1621261055
transform 1 0 8544 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_81
timestamp 1621261055
transform 1 0 8928 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_84
timestamp 1621261055
transform 1 0 9216 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_92
timestamp 1621261055
transform 1 0 9984 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_100
timestamp 1621261055
transform 1 0 10752 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_108
timestamp 1621261055
transform 1 0 11520 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_116
timestamp 1621261055
transform 1 0 12288 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_124
timestamp 1621261055
transform 1 0 13056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_596
timestamp 1621261055
transform 1 0 14400 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_132
timestamp 1621261055
transform 1 0 13824 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_136
timestamp 1621261055
transform 1 0 14208 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_139
timestamp 1621261055
transform 1 0 14496 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_147
timestamp 1621261055
transform 1 0 15264 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_155
timestamp 1621261055
transform 1 0 16032 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_163
timestamp 1621261055
transform 1 0 16800 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _132_
timestamp 1621261055
transform 1 0 19008 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _173_
timestamp 1621261055
transform 1 0 17568 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_40_174
timestamp 1621261055
transform 1 0 17856 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_182
timestamp 1621261055
transform 1 0 18624 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_40_189
timestamp 1621261055
transform 1 0 19296 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_597
timestamp 1621261055
transform 1 0 19680 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_194
timestamp 1621261055
transform 1 0 19776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_202
timestamp 1621261055
transform 1 0 20544 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_210
timestamp 1621261055
transform 1 0 21312 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_218
timestamp 1621261055
transform 1 0 22080 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_226
timestamp 1621261055
transform 1 0 22848 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_598
timestamp 1621261055
transform 1 0 24960 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_234
timestamp 1621261055
transform 1 0 23616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_242
timestamp 1621261055
transform 1 0 24384 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_246
timestamp 1621261055
transform 1 0 24768 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_249
timestamp 1621261055
transform 1 0 25056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_257
timestamp 1621261055
transform 1 0 25824 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_265
timestamp 1621261055
transform 1 0 26592 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_273
timestamp 1621261055
transform 1 0 27360 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_281
timestamp 1621261055
transform 1 0 28128 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_289
timestamp 1621261055
transform 1 0 28896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_599
timestamp 1621261055
transform 1 0 30240 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_297
timestamp 1621261055
transform 1 0 29664 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_301
timestamp 1621261055
transform 1 0 30048 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_304
timestamp 1621261055
transform 1 0 30336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_312
timestamp 1621261055
transform 1 0 31104 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_320
timestamp 1621261055
transform 1 0 31872 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_328
timestamp 1621261055
transform 1 0 32640 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_336
timestamp 1621261055
transform 1 0 33408 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_344
timestamp 1621261055
transform 1 0 34176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_352
timestamp 1621261055
transform 1 0 34944 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_356
timestamp 1621261055
transform 1 0 35328 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_600
timestamp 1621261055
transform 1 0 35520 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_359
timestamp 1621261055
transform 1 0 35616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_367
timestamp 1621261055
transform 1 0 36384 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_375
timestamp 1621261055
transform 1 0 37152 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_383
timestamp 1621261055
transform 1 0 37920 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_391
timestamp 1621261055
transform 1 0 38688 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_399
timestamp 1621261055
transform 1 0 39456 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _200_
timestamp 1621261055
transform 1 0 40128 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_601
timestamp 1621261055
transform 1 0 40800 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_403
timestamp 1621261055
transform 1 0 39840 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_40_405
timestamp 1621261055
transform 1 0 40032 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_409
timestamp 1621261055
transform 1 0 40416 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_40_414
timestamp 1621261055
transform 1 0 40896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_422
timestamp 1621261055
transform 1 0 41664 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_430
timestamp 1621261055
transform 1 0 42432 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_438
timestamp 1621261055
transform 1 0 43200 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_446
timestamp 1621261055
transform 1 0 43968 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_454
timestamp 1621261055
transform 1 0 44736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_462
timestamp 1621261055
transform 1 0 45504 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_602
timestamp 1621261055
transform 1 0 46080 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_466
timestamp 1621261055
transform 1 0 45888 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_469
timestamp 1621261055
transform 1 0 46176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_477
timestamp 1621261055
transform 1 0 46944 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_485
timestamp 1621261055
transform 1 0 47712 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_493
timestamp 1621261055
transform 1 0 48480 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_501
timestamp 1621261055
transform 1 0 49248 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _121_
timestamp 1621261055
transform 1 0 49824 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_603
timestamp 1621261055
transform 1 0 51360 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_505
timestamp 1621261055
transform 1 0 49632 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_510
timestamp 1621261055
transform 1 0 50112 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_518
timestamp 1621261055
transform 1 0 50880 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_40_522
timestamp 1621261055
transform 1 0 51264 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_524
timestamp 1621261055
transform 1 0 51456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _021_
timestamp 1621261055
transform 1 0 52416 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _078_
timestamp 1621261055
transform 1 0 53472 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_35
timestamp 1621261055
transform 1 0 52224 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_537
timestamp 1621261055
transform 1 0 52704 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _165_
timestamp 1621261055
transform 1 0 54336 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _172_
timestamp 1621261055
transform 1 0 55488 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_40_548
timestamp 1621261055
transform 1 0 53760 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_552
timestamp 1621261055
transform 1 0 54144 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_557
timestamp 1621261055
transform 1 0 54624 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_40_565
timestamp 1621261055
transform 1 0 55392 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_604
timestamp 1621261055
transform 1 0 56640 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_569
timestamp 1621261055
transform 1 0 55776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_40_577
timestamp 1621261055
transform 1 0 56544 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_579
timestamp 1621261055
transform 1 0 56736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_587
timestamp 1621261055
transform 1 0 57504 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_81
timestamp 1621261055
transform -1 0 58848 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_595
timestamp 1621261055
transform 1 0 58272 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_82
timestamp 1621261055
transform 1 0 1152 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_41_4
timestamp 1621261055
transform 1 0 1536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_12
timestamp 1621261055
transform 1 0 2304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_20
timestamp 1621261055
transform 1 0 3072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_28
timestamp 1621261055
transform 1 0 3840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_36
timestamp 1621261055
transform 1 0 4608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_605
timestamp 1621261055
transform 1 0 6432 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_44
timestamp 1621261055
transform 1 0 5376 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_52
timestamp 1621261055
transform 1 0 6144 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_41_54
timestamp 1621261055
transform 1 0 6336 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_56
timestamp 1621261055
transform 1 0 6528 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_64
timestamp 1621261055
transform 1 0 7296 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_72
timestamp 1621261055
transform 1 0 8064 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_80
timestamp 1621261055
transform 1 0 8832 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_88
timestamp 1621261055
transform 1 0 9600 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_96
timestamp 1621261055
transform 1 0 10368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_104
timestamp 1621261055
transform 1 0 11136 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_606
timestamp 1621261055
transform 1 0 11712 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_108
timestamp 1621261055
transform 1 0 11520 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_111
timestamp 1621261055
transform 1 0 11808 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_119
timestamp 1621261055
transform 1 0 12576 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_127
timestamp 1621261055
transform 1 0 13344 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_135
timestamp 1621261055
transform 1 0 14112 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_143
timestamp 1621261055
transform 1 0 14880 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_607
timestamp 1621261055
transform 1 0 16992 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_151
timestamp 1621261055
transform 1 0 15648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_159
timestamp 1621261055
transform 1 0 16416 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_163
timestamp 1621261055
transform 1 0 16800 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_166
timestamp 1621261055
transform 1 0 17088 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_174
timestamp 1621261055
transform 1 0 17856 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_182
timestamp 1621261055
transform 1 0 18624 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_190
timestamp 1621261055
transform 1 0 19392 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_198
timestamp 1621261055
transform 1 0 20160 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_206
timestamp 1621261055
transform 1 0 20928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_608
timestamp 1621261055
transform 1 0 22272 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_214
timestamp 1621261055
transform 1 0 21696 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_218
timestamp 1621261055
transform 1 0 22080 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_221
timestamp 1621261055
transform 1 0 22368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_229
timestamp 1621261055
transform 1 0 23136 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_237
timestamp 1621261055
transform 1 0 23904 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_245
timestamp 1621261055
transform 1 0 24672 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_253
timestamp 1621261055
transform 1 0 25440 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_261
timestamp 1621261055
transform 1 0 26208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_269
timestamp 1621261055
transform 1 0 26976 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_273
timestamp 1621261055
transform 1 0 27360 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_609
timestamp 1621261055
transform 1 0 27552 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_276
timestamp 1621261055
transform 1 0 27648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_284
timestamp 1621261055
transform 1 0 28416 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_292
timestamp 1621261055
transform 1 0 29184 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _211_
timestamp 1621261055
transform 1 0 29760 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_296
timestamp 1621261055
transform 1 0 29568 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_301
timestamp 1621261055
transform 1 0 30048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_309
timestamp 1621261055
transform 1 0 30816 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _086_
timestamp 1621261055
transform 1 0 31584 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_610
timestamp 1621261055
transform 1 0 32832 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_320
timestamp 1621261055
transform 1 0 31872 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_328
timestamp 1621261055
transform 1 0 32640 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_331
timestamp 1621261055
transform 1 0 32928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_339
timestamp 1621261055
transform 1 0 33696 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_347
timestamp 1621261055
transform 1 0 34464 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_355
timestamp 1621261055
transform 1 0 35232 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_363
timestamp 1621261055
transform 1 0 36000 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_371
timestamp 1621261055
transform 1 0 36768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_611
timestamp 1621261055
transform 1 0 38112 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_379
timestamp 1621261055
transform 1 0 37536 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_383
timestamp 1621261055
transform 1 0 37920 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_386
timestamp 1621261055
transform 1 0 38208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_394
timestamp 1621261055
transform 1 0 38976 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_402
timestamp 1621261055
transform 1 0 39744 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_410
timestamp 1621261055
transform 1 0 40512 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_418
timestamp 1621261055
transform 1 0 41280 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_612
timestamp 1621261055
transform 1 0 43392 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_426
timestamp 1621261055
transform 1 0 42048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_434
timestamp 1621261055
transform 1 0 42816 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_438
timestamp 1621261055
transform 1 0 43200 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_441
timestamp 1621261055
transform 1 0 43488 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_449
timestamp 1621261055
transform 1 0 44256 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_457
timestamp 1621261055
transform 1 0 45024 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_465
timestamp 1621261055
transform 1 0 45792 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_473
timestamp 1621261055
transform 1 0 46560 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_481
timestamp 1621261055
transform 1 0 47328 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_613
timestamp 1621261055
transform 1 0 48672 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_489
timestamp 1621261055
transform 1 0 48096 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_493
timestamp 1621261055
transform 1 0 48480 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_496
timestamp 1621261055
transform 1 0 48768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_504
timestamp 1621261055
transform 1 0 49536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_512
timestamp 1621261055
transform 1 0 50304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_520
timestamp 1621261055
transform 1 0 51072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_528
timestamp 1621261055
transform 1 0 51840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_536
timestamp 1621261055
transform 1 0 52608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_544
timestamp 1621261055
transform 1 0 53376 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_614
timestamp 1621261055
transform 1 0 53952 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_548
timestamp 1621261055
transform 1 0 53760 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_551
timestamp 1621261055
transform 1 0 54048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_559
timestamp 1621261055
transform 1 0 54816 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_567
timestamp 1621261055
transform 1 0 55584 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_575
timestamp 1621261055
transform 1 0 56352 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_583
timestamp 1621261055
transform 1 0 57120 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_83
timestamp 1621261055
transform -1 0 58848 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_41_591
timestamp 1621261055
transform 1 0 57888 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_595
timestamp 1621261055
transform 1 0 58272 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_84
timestamp 1621261055
transform 1 0 1152 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_42_4
timestamp 1621261055
transform 1 0 1536 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_12
timestamp 1621261055
transform 1 0 2304 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_20
timestamp 1621261055
transform 1 0 3072 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_615
timestamp 1621261055
transform 1 0 3840 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_29
timestamp 1621261055
transform 1 0 3936 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_37
timestamp 1621261055
transform 1 0 4704 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_45
timestamp 1621261055
transform 1 0 5472 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_53
timestamp 1621261055
transform 1 0 6240 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_61
timestamp 1621261055
transform 1 0 7008 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_616
timestamp 1621261055
transform 1 0 9120 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_69
timestamp 1621261055
transform 1 0 7776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_77
timestamp 1621261055
transform 1 0 8544 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_81
timestamp 1621261055
transform 1 0 8928 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_84
timestamp 1621261055
transform 1 0 9216 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_92
timestamp 1621261055
transform 1 0 9984 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_100
timestamp 1621261055
transform 1 0 10752 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_108
timestamp 1621261055
transform 1 0 11520 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_116
timestamp 1621261055
transform 1 0 12288 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_124
timestamp 1621261055
transform 1 0 13056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_617
timestamp 1621261055
transform 1 0 14400 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_132
timestamp 1621261055
transform 1 0 13824 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_136
timestamp 1621261055
transform 1 0 14208 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_139
timestamp 1621261055
transform 1 0 14496 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_147
timestamp 1621261055
transform 1 0 15264 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _053_
timestamp 1621261055
transform 1 0 16704 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_42_155
timestamp 1621261055
transform 1 0 16032 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_159
timestamp 1621261055
transform 1 0 16416 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_42_161
timestamp 1621261055
transform 1 0 16608 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_165
timestamp 1621261055
transform 1 0 16992 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _135_
timestamp 1621261055
transform 1 0 17376 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_172
timestamp 1621261055
transform 1 0 17664 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_180
timestamp 1621261055
transform 1 0 18432 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_188
timestamp 1621261055
transform 1 0 19200 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_618
timestamp 1621261055
transform 1 0 19680 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_42_192
timestamp 1621261055
transform 1 0 19584 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_194
timestamp 1621261055
transform 1 0 19776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_202
timestamp 1621261055
transform 1 0 20544 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_210
timestamp 1621261055
transform 1 0 21312 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_218
timestamp 1621261055
transform 1 0 22080 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_226
timestamp 1621261055
transform 1 0 22848 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_619
timestamp 1621261055
transform 1 0 24960 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_234
timestamp 1621261055
transform 1 0 23616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_242
timestamp 1621261055
transform 1 0 24384 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_246
timestamp 1621261055
transform 1 0 24768 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_249
timestamp 1621261055
transform 1 0 25056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_257
timestamp 1621261055
transform 1 0 25824 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_265
timestamp 1621261055
transform 1 0 26592 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_273
timestamp 1621261055
transform 1 0 27360 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_281
timestamp 1621261055
transform 1 0 28128 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_289
timestamp 1621261055
transform 1 0 28896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_620
timestamp 1621261055
transform 1 0 30240 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_297
timestamp 1621261055
transform 1 0 29664 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_301
timestamp 1621261055
transform 1 0 30048 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_304
timestamp 1621261055
transform 1 0 30336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_312
timestamp 1621261055
transform 1 0 31104 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_320
timestamp 1621261055
transform 1 0 31872 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_328
timestamp 1621261055
transform 1 0 32640 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_336
timestamp 1621261055
transform 1 0 33408 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_344
timestamp 1621261055
transform 1 0 34176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_352
timestamp 1621261055
transform 1 0 34944 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_356
timestamp 1621261055
transform 1 0 35328 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_621
timestamp 1621261055
transform 1 0 35520 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_359
timestamp 1621261055
transform 1 0 35616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_367
timestamp 1621261055
transform 1 0 36384 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_375
timestamp 1621261055
transform 1 0 37152 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_383
timestamp 1621261055
transform 1 0 37920 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_391
timestamp 1621261055
transform 1 0 38688 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_399
timestamp 1621261055
transform 1 0 39456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_622
timestamp 1621261055
transform 1 0 40800 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_407
timestamp 1621261055
transform 1 0 40224 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_411
timestamp 1621261055
transform 1 0 40608 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_414
timestamp 1621261055
transform 1 0 40896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_422
timestamp 1621261055
transform 1 0 41664 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_430
timestamp 1621261055
transform 1 0 42432 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_438
timestamp 1621261055
transform 1 0 43200 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_446
timestamp 1621261055
transform 1 0 43968 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_454
timestamp 1621261055
transform 1 0 44736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_462
timestamp 1621261055
transform 1 0 45504 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_623
timestamp 1621261055
transform 1 0 46080 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_466
timestamp 1621261055
transform 1 0 45888 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_469
timestamp 1621261055
transform 1 0 46176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_477
timestamp 1621261055
transform 1 0 46944 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_485
timestamp 1621261055
transform 1 0 47712 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_493
timestamp 1621261055
transform 1 0 48480 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_501
timestamp 1621261055
transform 1 0 49248 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_624
timestamp 1621261055
transform 1 0 51360 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_509
timestamp 1621261055
transform 1 0 50016 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_517
timestamp 1621261055
transform 1 0 50784 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_521
timestamp 1621261055
transform 1 0 51168 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_524
timestamp 1621261055
transform 1 0 51456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_532
timestamp 1621261055
transform 1 0 52224 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_540
timestamp 1621261055
transform 1 0 52992 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_548
timestamp 1621261055
transform 1 0 53760 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_556
timestamp 1621261055
transform 1 0 54528 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_564
timestamp 1621261055
transform 1 0 55296 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_625
timestamp 1621261055
transform 1 0 56640 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_572
timestamp 1621261055
transform 1 0 56064 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_576
timestamp 1621261055
transform 1 0 56448 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_579
timestamp 1621261055
transform 1 0 56736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_587
timestamp 1621261055
transform 1 0 57504 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_85
timestamp 1621261055
transform -1 0 58848 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_595
timestamp 1621261055
transform 1 0 58272 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_86
timestamp 1621261055
transform 1 0 1152 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_43_4
timestamp 1621261055
transform 1 0 1536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_12
timestamp 1621261055
transform 1 0 2304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_20
timestamp 1621261055
transform 1 0 3072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_28
timestamp 1621261055
transform 1 0 3840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_36
timestamp 1621261055
transform 1 0 4608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_626
timestamp 1621261055
transform 1 0 6432 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_44
timestamp 1621261055
transform 1 0 5376 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_52
timestamp 1621261055
transform 1 0 6144 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_43_54
timestamp 1621261055
transform 1 0 6336 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_56
timestamp 1621261055
transform 1 0 6528 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_64
timestamp 1621261055
transform 1 0 7296 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_72
timestamp 1621261055
transform 1 0 8064 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_80
timestamp 1621261055
transform 1 0 8832 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_88
timestamp 1621261055
transform 1 0 9600 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_96
timestamp 1621261055
transform 1 0 10368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_104
timestamp 1621261055
transform 1 0 11136 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_627
timestamp 1621261055
transform 1 0 11712 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_108
timestamp 1621261055
transform 1 0 11520 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_111
timestamp 1621261055
transform 1 0 11808 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_119
timestamp 1621261055
transform 1 0 12576 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_127
timestamp 1621261055
transform 1 0 13344 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_135
timestamp 1621261055
transform 1 0 14112 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_143
timestamp 1621261055
transform 1 0 14880 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_628
timestamp 1621261055
transform 1 0 16992 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_151
timestamp 1621261055
transform 1 0 15648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_159
timestamp 1621261055
transform 1 0 16416 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_163
timestamp 1621261055
transform 1 0 16800 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_166
timestamp 1621261055
transform 1 0 17088 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_174
timestamp 1621261055
transform 1 0 17856 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_182
timestamp 1621261055
transform 1 0 18624 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_190
timestamp 1621261055
transform 1 0 19392 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_198
timestamp 1621261055
transform 1 0 20160 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_206
timestamp 1621261055
transform 1 0 20928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_629
timestamp 1621261055
transform 1 0 22272 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_214
timestamp 1621261055
transform 1 0 21696 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_218
timestamp 1621261055
transform 1 0 22080 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_221
timestamp 1621261055
transform 1 0 22368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_229
timestamp 1621261055
transform 1 0 23136 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_237
timestamp 1621261055
transform 1 0 23904 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_245
timestamp 1621261055
transform 1 0 24672 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_253
timestamp 1621261055
transform 1 0 25440 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_261
timestamp 1621261055
transform 1 0 26208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_269
timestamp 1621261055
transform 1 0 26976 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_273
timestamp 1621261055
transform 1 0 27360 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_630
timestamp 1621261055
transform 1 0 27552 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_276
timestamp 1621261055
transform 1 0 27648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_284
timestamp 1621261055
transform 1 0 28416 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_292
timestamp 1621261055
transform 1 0 29184 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_300
timestamp 1621261055
transform 1 0 29952 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_308
timestamp 1621261055
transform 1 0 30720 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_631
timestamp 1621261055
transform 1 0 32832 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_316
timestamp 1621261055
transform 1 0 31488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_324
timestamp 1621261055
transform 1 0 32256 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_328
timestamp 1621261055
transform 1 0 32640 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_331
timestamp 1621261055
transform 1 0 32928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_339
timestamp 1621261055
transform 1 0 33696 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_347
timestamp 1621261055
transform 1 0 34464 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_355
timestamp 1621261055
transform 1 0 35232 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_363
timestamp 1621261055
transform 1 0 36000 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_371
timestamp 1621261055
transform 1 0 36768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_632
timestamp 1621261055
transform 1 0 38112 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_379
timestamp 1621261055
transform 1 0 37536 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_383
timestamp 1621261055
transform 1 0 37920 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_386
timestamp 1621261055
transform 1 0 38208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_394
timestamp 1621261055
transform 1 0 38976 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_398
timestamp 1621261055
transform 1 0 39360 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _052_
timestamp 1621261055
transform 1 0 39648 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_43_400
timestamp 1621261055
transform 1 0 39552 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_404
timestamp 1621261055
transform 1 0 39936 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_412
timestamp 1621261055
transform 1 0 40704 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_420
timestamp 1621261055
transform 1 0 41472 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_633
timestamp 1621261055
transform 1 0 43392 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_428
timestamp 1621261055
transform 1 0 42240 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_436
timestamp 1621261055
transform 1 0 43008 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_43_441
timestamp 1621261055
transform 1 0 43488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_449
timestamp 1621261055
transform 1 0 44256 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_457
timestamp 1621261055
transform 1 0 45024 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_465
timestamp 1621261055
transform 1 0 45792 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_473
timestamp 1621261055
transform 1 0 46560 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_481
timestamp 1621261055
transform 1 0 47328 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_634
timestamp 1621261055
transform 1 0 48672 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_489
timestamp 1621261055
transform 1 0 48096 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_493
timestamp 1621261055
transform 1 0 48480 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_496
timestamp 1621261055
transform 1 0 48768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_504
timestamp 1621261055
transform 1 0 49536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_512
timestamp 1621261055
transform 1 0 50304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_520
timestamp 1621261055
transform 1 0 51072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_528
timestamp 1621261055
transform 1 0 51840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_536
timestamp 1621261055
transform 1 0 52608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_544
timestamp 1621261055
transform 1 0 53376 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_635
timestamp 1621261055
transform 1 0 53952 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_548
timestamp 1621261055
transform 1 0 53760 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_551
timestamp 1621261055
transform 1 0 54048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_559
timestamp 1621261055
transform 1 0 54816 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_567
timestamp 1621261055
transform 1 0 55584 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_575
timestamp 1621261055
transform 1 0 56352 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_583
timestamp 1621261055
transform 1 0 57120 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_587
timestamp 1621261055
transform 1 0 57504 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _146_
timestamp 1621261055
transform 1 0 57792 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_87
timestamp 1621261055
transform -1 0 58848 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_43_589
timestamp 1621261055
transform 1 0 57696 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_593
timestamp 1621261055
transform 1 0 58080 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_88
timestamp 1621261055
transform 1 0 1152 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_44_4
timestamp 1621261055
transform 1 0 1536 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_12
timestamp 1621261055
transform 1 0 2304 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_20
timestamp 1621261055
transform 1 0 3072 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_636
timestamp 1621261055
transform 1 0 3840 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_29
timestamp 1621261055
transform 1 0 3936 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_37
timestamp 1621261055
transform 1 0 4704 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_45
timestamp 1621261055
transform 1 0 5472 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_53
timestamp 1621261055
transform 1 0 6240 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_61
timestamp 1621261055
transform 1 0 7008 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_637
timestamp 1621261055
transform 1 0 9120 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_69
timestamp 1621261055
transform 1 0 7776 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_77
timestamp 1621261055
transform 1 0 8544 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_81
timestamp 1621261055
transform 1 0 8928 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_84
timestamp 1621261055
transform 1 0 9216 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_92
timestamp 1621261055
transform 1 0 9984 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_100
timestamp 1621261055
transform 1 0 10752 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_108
timestamp 1621261055
transform 1 0 11520 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_116
timestamp 1621261055
transform 1 0 12288 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_124
timestamp 1621261055
transform 1 0 13056 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _091_
timestamp 1621261055
transform 1 0 13728 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_638
timestamp 1621261055
transform 1 0 14400 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_128
timestamp 1621261055
transform 1 0 13440 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_44_130
timestamp 1621261055
transform 1 0 13632 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_134
timestamp 1621261055
transform 1 0 14016 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_44_139
timestamp 1621261055
transform 1 0 14496 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_147
timestamp 1621261055
transform 1 0 15264 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_155
timestamp 1621261055
transform 1 0 16032 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_163
timestamp 1621261055
transform 1 0 16800 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _000_
timestamp 1621261055
transform 1 0 19008 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_44_171
timestamp 1621261055
transform 1 0 17568 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_179
timestamp 1621261055
transform 1 0 18336 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_183
timestamp 1621261055
transform 1 0 18720 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_44_185
timestamp 1621261055
transform 1 0 18912 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_189
timestamp 1621261055
transform 1 0 19296 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_639
timestamp 1621261055
transform 1 0 19680 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_194
timestamp 1621261055
transform 1 0 19776 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_202
timestamp 1621261055
transform 1 0 20544 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_210
timestamp 1621261055
transform 1 0 21312 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_218
timestamp 1621261055
transform 1 0 22080 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_226
timestamp 1621261055
transform 1 0 22848 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_640
timestamp 1621261055
transform 1 0 24960 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_234
timestamp 1621261055
transform 1 0 23616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_242
timestamp 1621261055
transform 1 0 24384 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_246
timestamp 1621261055
transform 1 0 24768 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_249
timestamp 1621261055
transform 1 0 25056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_257
timestamp 1621261055
transform 1 0 25824 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_265
timestamp 1621261055
transform 1 0 26592 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_273
timestamp 1621261055
transform 1 0 27360 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_281
timestamp 1621261055
transform 1 0 28128 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_289
timestamp 1621261055
transform 1 0 28896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _134_
timestamp 1621261055
transform 1 0 30720 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_641
timestamp 1621261055
transform 1 0 30240 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_297
timestamp 1621261055
transform 1 0 29664 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_301
timestamp 1621261055
transform 1 0 30048 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_44_304
timestamp 1621261055
transform 1 0 30336 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_44_311
timestamp 1621261055
transform 1 0 31008 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_319
timestamp 1621261055
transform 1 0 31776 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_327
timestamp 1621261055
transform 1 0 32544 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_335
timestamp 1621261055
transform 1 0 33312 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _111_
timestamp 1621261055
transform 1 0 33888 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_339
timestamp 1621261055
transform 1 0 33696 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_344
timestamp 1621261055
transform 1 0 34176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_352
timestamp 1621261055
transform 1 0 34944 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_356
timestamp 1621261055
transform 1 0 35328 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_642
timestamp 1621261055
transform 1 0 35520 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_359
timestamp 1621261055
transform 1 0 35616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_367
timestamp 1621261055
transform 1 0 36384 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_375
timestamp 1621261055
transform 1 0 37152 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_383
timestamp 1621261055
transform 1 0 37920 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_391
timestamp 1621261055
transform 1 0 38688 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_399
timestamp 1621261055
transform 1 0 39456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_643
timestamp 1621261055
transform 1 0 40800 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_407
timestamp 1621261055
transform 1 0 40224 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_411
timestamp 1621261055
transform 1 0 40608 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_414
timestamp 1621261055
transform 1 0 40896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_422
timestamp 1621261055
transform 1 0 41664 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_430
timestamp 1621261055
transform 1 0 42432 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_438
timestamp 1621261055
transform 1 0 43200 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_446
timestamp 1621261055
transform 1 0 43968 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_454
timestamp 1621261055
transform 1 0 44736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_462
timestamp 1621261055
transform 1 0 45504 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_644
timestamp 1621261055
transform 1 0 46080 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_466
timestamp 1621261055
transform 1 0 45888 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_469
timestamp 1621261055
transform 1 0 46176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_477
timestamp 1621261055
transform 1 0 46944 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_485
timestamp 1621261055
transform 1 0 47712 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_493
timestamp 1621261055
transform 1 0 48480 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_501
timestamp 1621261055
transform 1 0 49248 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_645
timestamp 1621261055
transform 1 0 51360 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_509
timestamp 1621261055
transform 1 0 50016 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_517
timestamp 1621261055
transform 1 0 50784 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_521
timestamp 1621261055
transform 1 0 51168 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_524
timestamp 1621261055
transform 1 0 51456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_532
timestamp 1621261055
transform 1 0 52224 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_540
timestamp 1621261055
transform 1 0 52992 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_548
timestamp 1621261055
transform 1 0 53760 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_556
timestamp 1621261055
transform 1 0 54528 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_564
timestamp 1621261055
transform 1 0 55296 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_646
timestamp 1621261055
transform 1 0 56640 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_572
timestamp 1621261055
transform 1 0 56064 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_576
timestamp 1621261055
transform 1 0 56448 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_579
timestamp 1621261055
transform 1 0 56736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_587
timestamp 1621261055
transform 1 0 57504 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_89
timestamp 1621261055
transform -1 0 58848 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_595
timestamp 1621261055
transform 1 0 58272 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_90
timestamp 1621261055
transform 1 0 1152 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_4
timestamp 1621261055
transform 1 0 1536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_12
timestamp 1621261055
transform 1 0 2304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_20
timestamp 1621261055
transform 1 0 3072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_28
timestamp 1621261055
transform 1 0 3840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_36
timestamp 1621261055
transform 1 0 4608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_647
timestamp 1621261055
transform 1 0 6432 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_44
timestamp 1621261055
transform 1 0 5376 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_52
timestamp 1621261055
transform 1 0 6144 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_54
timestamp 1621261055
transform 1 0 6336 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_56
timestamp 1621261055
transform 1 0 6528 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_64
timestamp 1621261055
transform 1 0 7296 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_72
timestamp 1621261055
transform 1 0 8064 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_80
timestamp 1621261055
transform 1 0 8832 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_88
timestamp 1621261055
transform 1 0 9600 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_96
timestamp 1621261055
transform 1 0 10368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_104
timestamp 1621261055
transform 1 0 11136 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_648
timestamp 1621261055
transform 1 0 11712 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_108
timestamp 1621261055
transform 1 0 11520 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_111
timestamp 1621261055
transform 1 0 11808 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_119
timestamp 1621261055
transform 1 0 12576 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_127
timestamp 1621261055
transform 1 0 13344 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_135
timestamp 1621261055
transform 1 0 14112 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_143
timestamp 1621261055
transform 1 0 14880 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_649
timestamp 1621261055
transform 1 0 16992 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_151
timestamp 1621261055
transform 1 0 15648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_159
timestamp 1621261055
transform 1 0 16416 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_163
timestamp 1621261055
transform 1 0 16800 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_166
timestamp 1621261055
transform 1 0 17088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _058_
timestamp 1621261055
transform 1 0 18816 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_45_174
timestamp 1621261055
transform 1 0 17856 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_182
timestamp 1621261055
transform 1 0 18624 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_187
timestamp 1621261055
transform 1 0 19104 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_195
timestamp 1621261055
transform 1 0 19872 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_203
timestamp 1621261055
transform 1 0 20640 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_650
timestamp 1621261055
transform 1 0 22272 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_211
timestamp 1621261055
transform 1 0 21408 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_45_219
timestamp 1621261055
transform 1 0 22176 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_221
timestamp 1621261055
transform 1 0 22368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_229
timestamp 1621261055
transform 1 0 23136 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_237
timestamp 1621261055
transform 1 0 23904 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_245
timestamp 1621261055
transform 1 0 24672 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_253
timestamp 1621261055
transform 1 0 25440 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_261
timestamp 1621261055
transform 1 0 26208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_269
timestamp 1621261055
transform 1 0 26976 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_273
timestamp 1621261055
transform 1 0 27360 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _035_
timestamp 1621261055
transform 1 0 28032 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_651
timestamp 1621261055
transform 1 0 27552 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_276
timestamp 1621261055
transform 1 0 27648 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_283
timestamp 1621261055
transform 1 0 28320 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_291
timestamp 1621261055
transform 1 0 29088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_299
timestamp 1621261055
transform 1 0 29856 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_307
timestamp 1621261055
transform 1 0 30624 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_315
timestamp 1621261055
transform 1 0 31392 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_652
timestamp 1621261055
transform 1 0 32832 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_323
timestamp 1621261055
transform 1 0 32160 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_327
timestamp 1621261055
transform 1 0 32544 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_329
timestamp 1621261055
transform 1 0 32736 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_331
timestamp 1621261055
transform 1 0 32928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_339
timestamp 1621261055
transform 1 0 33696 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_347
timestamp 1621261055
transform 1 0 34464 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_355
timestamp 1621261055
transform 1 0 35232 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_363
timestamp 1621261055
transform 1 0 36000 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_371
timestamp 1621261055
transform 1 0 36768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_653
timestamp 1621261055
transform 1 0 38112 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_379
timestamp 1621261055
transform 1 0 37536 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_383
timestamp 1621261055
transform 1 0 37920 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_386
timestamp 1621261055
transform 1 0 38208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_394
timestamp 1621261055
transform 1 0 38976 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_402
timestamp 1621261055
transform 1 0 39744 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_410
timestamp 1621261055
transform 1 0 40512 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_418
timestamp 1621261055
transform 1 0 41280 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _063_
timestamp 1621261055
transform 1 0 42144 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_654
timestamp 1621261055
transform 1 0 43392 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_45_426
timestamp 1621261055
transform 1 0 42048 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_430
timestamp 1621261055
transform 1 0 42432 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_438
timestamp 1621261055
transform 1 0 43200 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_441
timestamp 1621261055
transform 1 0 43488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_449
timestamp 1621261055
transform 1 0 44256 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_457
timestamp 1621261055
transform 1 0 45024 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _040_
timestamp 1621261055
transform 1 0 47520 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_45_465
timestamp 1621261055
transform 1 0 45792 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_473
timestamp 1621261055
transform 1 0 46560 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_481
timestamp 1621261055
transform 1 0 47328 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_655
timestamp 1621261055
transform 1 0 48672 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_486
timestamp 1621261055
transform 1 0 47808 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_45_494
timestamp 1621261055
transform 1 0 48576 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_496
timestamp 1621261055
transform 1 0 48768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_504
timestamp 1621261055
transform 1 0 49536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_512
timestamp 1621261055
transform 1 0 50304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_520
timestamp 1621261055
transform 1 0 51072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_528
timestamp 1621261055
transform 1 0 51840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_536
timestamp 1621261055
transform 1 0 52608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_544
timestamp 1621261055
transform 1 0 53376 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_656
timestamp 1621261055
transform 1 0 53952 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_548
timestamp 1621261055
transform 1 0 53760 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_551
timestamp 1621261055
transform 1 0 54048 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_559
timestamp 1621261055
transform 1 0 54816 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_567
timestamp 1621261055
transform 1 0 55584 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_575
timestamp 1621261055
transform 1 0 56352 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_583
timestamp 1621261055
transform 1 0 57120 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_91
timestamp 1621261055
transform -1 0 58848 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_45_591
timestamp 1621261055
transform 1 0 57888 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_595
timestamp 1621261055
transform 1 0 58272 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_92
timestamp 1621261055
transform 1 0 1152 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_94
timestamp 1621261055
transform 1 0 1152 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_4
timestamp 1621261055
transform 1 0 1536 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_12
timestamp 1621261055
transform 1 0 2304 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_20
timestamp 1621261055
transform 1 0 3072 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_4
timestamp 1621261055
transform 1 0 1536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_12
timestamp 1621261055
transform 1 0 2304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_20
timestamp 1621261055
transform 1 0 3072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_657
timestamp 1621261055
transform 1 0 3840 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_29
timestamp 1621261055
transform 1 0 3936 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_37
timestamp 1621261055
transform 1 0 4704 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_28
timestamp 1621261055
transform 1 0 3840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_36
timestamp 1621261055
transform 1 0 4608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_668
timestamp 1621261055
transform 1 0 6432 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_45
timestamp 1621261055
transform 1 0 5472 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_53
timestamp 1621261055
transform 1 0 6240 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_61
timestamp 1621261055
transform 1 0 7008 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_44
timestamp 1621261055
transform 1 0 5376 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_52
timestamp 1621261055
transform 1 0 6144 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_47_54
timestamp 1621261055
transform 1 0 6336 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_56
timestamp 1621261055
transform 1 0 6528 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_658
timestamp 1621261055
transform 1 0 9120 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_69
timestamp 1621261055
transform 1 0 7776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_77
timestamp 1621261055
transform 1 0 8544 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_81
timestamp 1621261055
transform 1 0 8928 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_84
timestamp 1621261055
transform 1 0 9216 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_64
timestamp 1621261055
transform 1 0 7296 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_72
timestamp 1621261055
transform 1 0 8064 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_80
timestamp 1621261055
transform 1 0 8832 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_92
timestamp 1621261055
transform 1 0 9984 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_100
timestamp 1621261055
transform 1 0 10752 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_88
timestamp 1621261055
transform 1 0 9600 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_96
timestamp 1621261055
transform 1 0 10368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_104
timestamp 1621261055
transform 1 0 11136 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_669
timestamp 1621261055
transform 1 0 11712 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_108
timestamp 1621261055
transform 1 0 11520 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_116
timestamp 1621261055
transform 1 0 12288 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_124
timestamp 1621261055
transform 1 0 13056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_108
timestamp 1621261055
transform 1 0 11520 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_111
timestamp 1621261055
transform 1 0 11808 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_119
timestamp 1621261055
transform 1 0 12576 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_659
timestamp 1621261055
transform 1 0 14400 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_132
timestamp 1621261055
transform 1 0 13824 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_136
timestamp 1621261055
transform 1 0 14208 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_139
timestamp 1621261055
transform 1 0 14496 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_147
timestamp 1621261055
transform 1 0 15264 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_127
timestamp 1621261055
transform 1 0 13344 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_135
timestamp 1621261055
transform 1 0 14112 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_143
timestamp 1621261055
transform 1 0 14880 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_670
timestamp 1621261055
transform 1 0 16992 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_155
timestamp 1621261055
transform 1 0 16032 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_163
timestamp 1621261055
transform 1 0 16800 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_151
timestamp 1621261055
transform 1 0 15648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_159
timestamp 1621261055
transform 1 0 16416 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_163
timestamp 1621261055
transform 1 0 16800 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_166
timestamp 1621261055
transform 1 0 17088 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_171
timestamp 1621261055
transform 1 0 17568 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_179
timestamp 1621261055
transform 1 0 18336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_187
timestamp 1621261055
transform 1 0 19104 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_174
timestamp 1621261055
transform 1 0 17856 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_182
timestamp 1621261055
transform 1 0 18624 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_660
timestamp 1621261055
transform 1 0 19680 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_191
timestamp 1621261055
transform 1 0 19488 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_194
timestamp 1621261055
transform 1 0 19776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_202
timestamp 1621261055
transform 1 0 20544 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_210
timestamp 1621261055
transform 1 0 21312 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_190
timestamp 1621261055
transform 1 0 19392 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_198
timestamp 1621261055
transform 1 0 20160 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_206
timestamp 1621261055
transform 1 0 20928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_671
timestamp 1621261055
transform 1 0 22272 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_218
timestamp 1621261055
transform 1 0 22080 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_226
timestamp 1621261055
transform 1 0 22848 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_214
timestamp 1621261055
transform 1 0 21696 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_218
timestamp 1621261055
transform 1 0 22080 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_221
timestamp 1621261055
transform 1 0 22368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_229
timestamp 1621261055
transform 1 0 23136 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_661
timestamp 1621261055
transform 1 0 24960 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_234
timestamp 1621261055
transform 1 0 23616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_242
timestamp 1621261055
transform 1 0 24384 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_246
timestamp 1621261055
transform 1 0 24768 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_249
timestamp 1621261055
transform 1 0 25056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_237
timestamp 1621261055
transform 1 0 23904 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_245
timestamp 1621261055
transform 1 0 24672 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_257
timestamp 1621261055
transform 1 0 25824 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_265
timestamp 1621261055
transform 1 0 26592 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_273
timestamp 1621261055
transform 1 0 27360 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_253
timestamp 1621261055
transform 1 0 25440 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_261
timestamp 1621261055
transform 1 0 26208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_269
timestamp 1621261055
transform 1 0 26976 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_273
timestamp 1621261055
transform 1 0 27360 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_672
timestamp 1621261055
transform 1 0 27552 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_281
timestamp 1621261055
transform 1 0 28128 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_289
timestamp 1621261055
transform 1 0 28896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_276
timestamp 1621261055
transform 1 0 27648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_284
timestamp 1621261055
transform 1 0 28416 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_292
timestamp 1621261055
transform 1 0 29184 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_662
timestamp 1621261055
transform 1 0 30240 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_297
timestamp 1621261055
transform 1 0 29664 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_301
timestamp 1621261055
transform 1 0 30048 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_304
timestamp 1621261055
transform 1 0 30336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_312
timestamp 1621261055
transform 1 0 31104 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_300
timestamp 1621261055
transform 1 0 29952 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_308
timestamp 1621261055
transform 1 0 30720 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_673
timestamp 1621261055
transform 1 0 32832 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_320
timestamp 1621261055
transform 1 0 31872 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_328
timestamp 1621261055
transform 1 0 32640 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_336
timestamp 1621261055
transform 1 0 33408 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_316
timestamp 1621261055
transform 1 0 31488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_324
timestamp 1621261055
transform 1 0 32256 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_328
timestamp 1621261055
transform 1 0 32640 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_331
timestamp 1621261055
transform 1 0 32928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_344
timestamp 1621261055
transform 1 0 34176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_352
timestamp 1621261055
transform 1 0 34944 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_356
timestamp 1621261055
transform 1 0 35328 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_339
timestamp 1621261055
transform 1 0 33696 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_347
timestamp 1621261055
transform 1 0 34464 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_355
timestamp 1621261055
transform 1 0 35232 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_663
timestamp 1621261055
transform 1 0 35520 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_359
timestamp 1621261055
transform 1 0 35616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_367
timestamp 1621261055
transform 1 0 36384 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_375
timestamp 1621261055
transform 1 0 37152 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_363
timestamp 1621261055
transform 1 0 36000 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_371
timestamp 1621261055
transform 1 0 36768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_674
timestamp 1621261055
transform 1 0 38112 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_383
timestamp 1621261055
transform 1 0 37920 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_391
timestamp 1621261055
transform 1 0 38688 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_399
timestamp 1621261055
transform 1 0 39456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_379
timestamp 1621261055
transform 1 0 37536 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_383
timestamp 1621261055
transform 1 0 37920 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_386
timestamp 1621261055
transform 1 0 38208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_394
timestamp 1621261055
transform 1 0 38976 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_664
timestamp 1621261055
transform 1 0 40800 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_407
timestamp 1621261055
transform 1 0 40224 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_411
timestamp 1621261055
transform 1 0 40608 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_414
timestamp 1621261055
transform 1 0 40896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_402
timestamp 1621261055
transform 1 0 39744 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_410
timestamp 1621261055
transform 1 0 40512 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_418
timestamp 1621261055
transform 1 0 41280 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_675
timestamp 1621261055
transform 1 0 43392 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_422
timestamp 1621261055
transform 1 0 41664 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_430
timestamp 1621261055
transform 1 0 42432 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_438
timestamp 1621261055
transform 1 0 43200 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_426
timestamp 1621261055
transform 1 0 42048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_434
timestamp 1621261055
transform 1 0 42816 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_438
timestamp 1621261055
transform 1 0 43200 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_441
timestamp 1621261055
transform 1 0 43488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_446
timestamp 1621261055
transform 1 0 43968 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_454
timestamp 1621261055
transform 1 0 44736 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_462
timestamp 1621261055
transform 1 0 45504 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_449
timestamp 1621261055
transform 1 0 44256 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_457
timestamp 1621261055
transform 1 0 45024 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _083_
timestamp 1621261055
transform 1 0 47040 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_665
timestamp 1621261055
transform 1 0 46080 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_466
timestamp 1621261055
transform 1 0 45888 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_469
timestamp 1621261055
transform 1 0 46176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_477
timestamp 1621261055
transform 1 0 46944 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_465
timestamp 1621261055
transform 1 0 45792 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_473
timestamp 1621261055
transform 1 0 46560 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_47_477
timestamp 1621261055
transform 1 0 46944 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_481
timestamp 1621261055
transform 1 0 47328 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_676
timestamp 1621261055
transform 1 0 48672 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_485
timestamp 1621261055
transform 1 0 47712 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_493
timestamp 1621261055
transform 1 0 48480 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_501
timestamp 1621261055
transform 1 0 49248 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_489
timestamp 1621261055
transform 1 0 48096 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_493
timestamp 1621261055
transform 1 0 48480 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_496
timestamp 1621261055
transform 1 0 48768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_504
timestamp 1621261055
transform 1 0 49536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_666
timestamp 1621261055
transform 1 0 51360 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_509
timestamp 1621261055
transform 1 0 50016 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_517
timestamp 1621261055
transform 1 0 50784 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_521
timestamp 1621261055
transform 1 0 51168 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_524
timestamp 1621261055
transform 1 0 51456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_512
timestamp 1621261055
transform 1 0 50304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_520
timestamp 1621261055
transform 1 0 51072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_532
timestamp 1621261055
transform 1 0 52224 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_540
timestamp 1621261055
transform 1 0 52992 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_528
timestamp 1621261055
transform 1 0 51840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_536
timestamp 1621261055
transform 1 0 52608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_544
timestamp 1621261055
transform 1 0 53376 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_677
timestamp 1621261055
transform 1 0 53952 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_548
timestamp 1621261055
transform 1 0 53760 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_556
timestamp 1621261055
transform 1 0 54528 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_564
timestamp 1621261055
transform 1 0 55296 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_548
timestamp 1621261055
transform 1 0 53760 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_551
timestamp 1621261055
transform 1 0 54048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_559
timestamp 1621261055
transform 1 0 54816 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_567
timestamp 1621261055
transform 1 0 55584 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _090_
timestamp 1621261055
transform -1 0 57600 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_667
timestamp 1621261055
transform 1 0 56640 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_142
timestamp 1621261055
transform -1 0 57312 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_572
timestamp 1621261055
transform 1 0 56064 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_576
timestamp 1621261055
transform 1 0 56448 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_579
timestamp 1621261055
transform 1 0 56736 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_588
timestamp 1621261055
transform 1 0 57600 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_575
timestamp 1621261055
transform 1 0 56352 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_583
timestamp 1621261055
transform 1 0 57120 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_93
timestamp 1621261055
transform -1 0 58848 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_95
timestamp 1621261055
transform -1 0 58848 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_46_596
timestamp 1621261055
transform 1 0 58368 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_47_591
timestamp 1621261055
transform 1 0 57888 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_595
timestamp 1621261055
transform 1 0 58272 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_96
timestamp 1621261055
transform 1 0 1152 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_4
timestamp 1621261055
transform 1 0 1536 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_12
timestamp 1621261055
transform 1 0 2304 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_20
timestamp 1621261055
transform 1 0 3072 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_678
timestamp 1621261055
transform 1 0 3840 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_29
timestamp 1621261055
transform 1 0 3936 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_37
timestamp 1621261055
transform 1 0 4704 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_45
timestamp 1621261055
transform 1 0 5472 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_53
timestamp 1621261055
transform 1 0 6240 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_61
timestamp 1621261055
transform 1 0 7008 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_679
timestamp 1621261055
transform 1 0 9120 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_69
timestamp 1621261055
transform 1 0 7776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_77
timestamp 1621261055
transform 1 0 8544 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_81
timestamp 1621261055
transform 1 0 8928 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_84
timestamp 1621261055
transform 1 0 9216 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_92
timestamp 1621261055
transform 1 0 9984 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_100
timestamp 1621261055
transform 1 0 10752 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_108
timestamp 1621261055
transform 1 0 11520 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_116
timestamp 1621261055
transform 1 0 12288 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_124
timestamp 1621261055
transform 1 0 13056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _095_
timestamp 1621261055
transform 1 0 14880 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_680
timestamp 1621261055
transform 1 0 14400 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_148
timestamp 1621261055
transform 1 0 14688 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_132
timestamp 1621261055
transform 1 0 13824 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_136
timestamp 1621261055
transform 1 0 14208 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_139
timestamp 1621261055
transform 1 0 14496 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_146
timestamp 1621261055
transform 1 0 15168 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_154
timestamp 1621261055
transform 1 0 15936 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_162
timestamp 1621261055
transform 1 0 16704 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_170
timestamp 1621261055
transform 1 0 17472 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_178
timestamp 1621261055
transform 1 0 18240 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_186
timestamp 1621261055
transform 1 0 19008 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_681
timestamp 1621261055
transform 1 0 19680 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_190
timestamp 1621261055
transform 1 0 19392 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_192
timestamp 1621261055
transform 1 0 19584 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_194
timestamp 1621261055
transform 1 0 19776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_202
timestamp 1621261055
transform 1 0 20544 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_210
timestamp 1621261055
transform 1 0 21312 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_218
timestamp 1621261055
transform 1 0 22080 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_226
timestamp 1621261055
transform 1 0 22848 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_682
timestamp 1621261055
transform 1 0 24960 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_234
timestamp 1621261055
transform 1 0 23616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_242
timestamp 1621261055
transform 1 0 24384 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_246
timestamp 1621261055
transform 1 0 24768 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_249
timestamp 1621261055
transform 1 0 25056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_257
timestamp 1621261055
transform 1 0 25824 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_265
timestamp 1621261055
transform 1 0 26592 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_273
timestamp 1621261055
transform 1 0 27360 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_281
timestamp 1621261055
transform 1 0 28128 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_289
timestamp 1621261055
transform 1 0 28896 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_683
timestamp 1621261055
transform 1 0 30240 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_297
timestamp 1621261055
transform 1 0 29664 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_301
timestamp 1621261055
transform 1 0 30048 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_304
timestamp 1621261055
transform 1 0 30336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_312
timestamp 1621261055
transform 1 0 31104 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _199_
timestamp 1621261055
transform -1 0 33024 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_216
timestamp 1621261055
transform -1 0 32736 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_320
timestamp 1621261055
transform 1 0 31872 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_324
timestamp 1621261055
transform 1 0 32256 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_326
timestamp 1621261055
transform 1 0 32448 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_332
timestamp 1621261055
transform 1 0 33024 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_340
timestamp 1621261055
transform 1 0 33792 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_348
timestamp 1621261055
transform 1 0 34560 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_356
timestamp 1621261055
transform 1 0 35328 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_684
timestamp 1621261055
transform 1 0 35520 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_359
timestamp 1621261055
transform 1 0 35616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_367
timestamp 1621261055
transform 1 0 36384 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_375
timestamp 1621261055
transform 1 0 37152 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_383
timestamp 1621261055
transform 1 0 37920 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_391
timestamp 1621261055
transform 1 0 38688 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_399
timestamp 1621261055
transform 1 0 39456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _043_
timestamp 1621261055
transform 1 0 41280 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_685
timestamp 1621261055
transform 1 0 40800 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_407
timestamp 1621261055
transform 1 0 40224 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_411
timestamp 1621261055
transform 1 0 40608 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_414
timestamp 1621261055
transform 1 0 40896 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_421
timestamp 1621261055
transform 1 0 41568 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_429
timestamp 1621261055
transform 1 0 42336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_437
timestamp 1621261055
transform 1 0 43104 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_445
timestamp 1621261055
transform 1 0 43872 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_453
timestamp 1621261055
transform 1 0 44640 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_461
timestamp 1621261055
transform 1 0 45408 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_686
timestamp 1621261055
transform 1 0 46080 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_465
timestamp 1621261055
transform 1 0 45792 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_467
timestamp 1621261055
transform 1 0 45984 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_469
timestamp 1621261055
transform 1 0 46176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_477
timestamp 1621261055
transform 1 0 46944 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_485
timestamp 1621261055
transform 1 0 47712 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_493
timestamp 1621261055
transform 1 0 48480 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_501
timestamp 1621261055
transform 1 0 49248 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_687
timestamp 1621261055
transform 1 0 51360 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_509
timestamp 1621261055
transform 1 0 50016 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_517
timestamp 1621261055
transform 1 0 50784 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_521
timestamp 1621261055
transform 1 0 51168 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_524
timestamp 1621261055
transform 1 0 51456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_532
timestamp 1621261055
transform 1 0 52224 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_540
timestamp 1621261055
transform 1 0 52992 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_548
timestamp 1621261055
transform 1 0 53760 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_556
timestamp 1621261055
transform 1 0 54528 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_564
timestamp 1621261055
transform 1 0 55296 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_688
timestamp 1621261055
transform 1 0 56640 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_572
timestamp 1621261055
transform 1 0 56064 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_576
timestamp 1621261055
transform 1 0 56448 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_579
timestamp 1621261055
transform 1 0 56736 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_587
timestamp 1621261055
transform 1 0 57504 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_97
timestamp 1621261055
transform -1 0 58848 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_595
timestamp 1621261055
transform 1 0 58272 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_98
timestamp 1621261055
transform 1 0 1152 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_49_4
timestamp 1621261055
transform 1 0 1536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_12
timestamp 1621261055
transform 1 0 2304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_20
timestamp 1621261055
transform 1 0 3072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_28
timestamp 1621261055
transform 1 0 3840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_36
timestamp 1621261055
transform 1 0 4608 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_689
timestamp 1621261055
transform 1 0 6432 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_44
timestamp 1621261055
transform 1 0 5376 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_52
timestamp 1621261055
transform 1 0 6144 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_54
timestamp 1621261055
transform 1 0 6336 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_56
timestamp 1621261055
transform 1 0 6528 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_64
timestamp 1621261055
transform 1 0 7296 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_72
timestamp 1621261055
transform 1 0 8064 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_80
timestamp 1621261055
transform 1 0 8832 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_88
timestamp 1621261055
transform 1 0 9600 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_96
timestamp 1621261055
transform 1 0 10368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_104
timestamp 1621261055
transform 1 0 11136 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_690
timestamp 1621261055
transform 1 0 11712 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_108
timestamp 1621261055
transform 1 0 11520 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_111
timestamp 1621261055
transform 1 0 11808 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_119
timestamp 1621261055
transform 1 0 12576 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_127
timestamp 1621261055
transform 1 0 13344 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_135
timestamp 1621261055
transform 1 0 14112 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_143
timestamp 1621261055
transform 1 0 14880 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_691
timestamp 1621261055
transform 1 0 16992 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_151
timestamp 1621261055
transform 1 0 15648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_159
timestamp 1621261055
transform 1 0 16416 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_163
timestamp 1621261055
transform 1 0 16800 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_166
timestamp 1621261055
transform 1 0 17088 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_174
timestamp 1621261055
transform 1 0 17856 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_182
timestamp 1621261055
transform 1 0 18624 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_190
timestamp 1621261055
transform 1 0 19392 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_198
timestamp 1621261055
transform 1 0 20160 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_206
timestamp 1621261055
transform 1 0 20928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_692
timestamp 1621261055
transform 1 0 22272 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_214
timestamp 1621261055
transform 1 0 21696 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_218
timestamp 1621261055
transform 1 0 22080 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_221
timestamp 1621261055
transform 1 0 22368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_229
timestamp 1621261055
transform 1 0 23136 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_237
timestamp 1621261055
transform 1 0 23904 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_245
timestamp 1621261055
transform 1 0 24672 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_253
timestamp 1621261055
transform 1 0 25440 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_261
timestamp 1621261055
transform 1 0 26208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_269
timestamp 1621261055
transform 1 0 26976 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_273
timestamp 1621261055
transform 1 0 27360 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_693
timestamp 1621261055
transform 1 0 27552 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_276
timestamp 1621261055
transform 1 0 27648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_284
timestamp 1621261055
transform 1 0 28416 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_292
timestamp 1621261055
transform 1 0 29184 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_300
timestamp 1621261055
transform 1 0 29952 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_308
timestamp 1621261055
transform 1 0 30720 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _115_
timestamp 1621261055
transform 1 0 33312 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_694
timestamp 1621261055
transform 1 0 32832 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_176
timestamp 1621261055
transform 1 0 33120 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_316
timestamp 1621261055
transform 1 0 31488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_324
timestamp 1621261055
transform 1 0 32256 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_328
timestamp 1621261055
transform 1 0 32640 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_331
timestamp 1621261055
transform 1 0 32928 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_338
timestamp 1621261055
transform 1 0 33600 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_346
timestamp 1621261055
transform 1 0 34368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_354
timestamp 1621261055
transform 1 0 35136 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _100_
timestamp 1621261055
transform 1 0 35808 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_358
timestamp 1621261055
transform 1 0 35520 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_360
timestamp 1621261055
transform 1 0 35712 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_364
timestamp 1621261055
transform 1 0 36096 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_372
timestamp 1621261055
transform 1 0 36864 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_695
timestamp 1621261055
transform 1 0 38112 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_380
timestamp 1621261055
transform 1 0 37632 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_49_384
timestamp 1621261055
transform 1 0 38016 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_386
timestamp 1621261055
transform 1 0 38208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_394
timestamp 1621261055
transform 1 0 38976 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_402
timestamp 1621261055
transform 1 0 39744 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_410
timestamp 1621261055
transform 1 0 40512 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_418
timestamp 1621261055
transform 1 0 41280 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_696
timestamp 1621261055
transform 1 0 43392 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_426
timestamp 1621261055
transform 1 0 42048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_434
timestamp 1621261055
transform 1 0 42816 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_438
timestamp 1621261055
transform 1 0 43200 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_441
timestamp 1621261055
transform 1 0 43488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_449
timestamp 1621261055
transform 1 0 44256 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_457
timestamp 1621261055
transform 1 0 45024 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_465
timestamp 1621261055
transform 1 0 45792 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_473
timestamp 1621261055
transform 1 0 46560 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_481
timestamp 1621261055
transform 1 0 47328 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_697
timestamp 1621261055
transform 1 0 48672 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_489
timestamp 1621261055
transform 1 0 48096 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_493
timestamp 1621261055
transform 1 0 48480 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_496
timestamp 1621261055
transform 1 0 48768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_504
timestamp 1621261055
transform 1 0 49536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_512
timestamp 1621261055
transform 1 0 50304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_520
timestamp 1621261055
transform 1 0 51072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _216_
timestamp 1621261055
transform 1 0 51840 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_49_531
timestamp 1621261055
transform 1 0 52128 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_539
timestamp 1621261055
transform 1 0 52896 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_698
timestamp 1621261055
transform 1 0 53952 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_547
timestamp 1621261055
transform 1 0 53664 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_549
timestamp 1621261055
transform 1 0 53856 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_551
timestamp 1621261055
transform 1 0 54048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_559
timestamp 1621261055
transform 1 0 54816 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_567
timestamp 1621261055
transform 1 0 55584 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_575
timestamp 1621261055
transform 1 0 56352 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_583
timestamp 1621261055
transform 1 0 57120 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_99
timestamp 1621261055
transform -1 0 58848 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_49_591
timestamp 1621261055
transform 1 0 57888 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_595
timestamp 1621261055
transform 1 0 58272 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_100
timestamp 1621261055
transform 1 0 1152 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_4
timestamp 1621261055
transform 1 0 1536 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_12
timestamp 1621261055
transform 1 0 2304 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_20
timestamp 1621261055
transform 1 0 3072 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_699
timestamp 1621261055
transform 1 0 3840 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_29
timestamp 1621261055
transform 1 0 3936 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_37
timestamp 1621261055
transform 1 0 4704 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_45
timestamp 1621261055
transform 1 0 5472 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_53
timestamp 1621261055
transform 1 0 6240 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_61
timestamp 1621261055
transform 1 0 7008 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_700
timestamp 1621261055
transform 1 0 9120 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_69
timestamp 1621261055
transform 1 0 7776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_77
timestamp 1621261055
transform 1 0 8544 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_81
timestamp 1621261055
transform 1 0 8928 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_84
timestamp 1621261055
transform 1 0 9216 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_92
timestamp 1621261055
transform 1 0 9984 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_100
timestamp 1621261055
transform 1 0 10752 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_108
timestamp 1621261055
transform 1 0 11520 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_116
timestamp 1621261055
transform 1 0 12288 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_124
timestamp 1621261055
transform 1 0 13056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _192_
timestamp 1621261055
transform -1 0 15456 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_701
timestamp 1621261055
transform 1 0 14400 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_238
timestamp 1621261055
transform -1 0 15168 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_50_132
timestamp 1621261055
transform 1 0 13824 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_136
timestamp 1621261055
transform 1 0 14208 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_50_139
timestamp 1621261055
transform 1 0 14496 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_50_143
timestamp 1621261055
transform 1 0 14880 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_149
timestamp 1621261055
transform 1 0 15456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_157
timestamp 1621261055
transform 1 0 16224 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_165
timestamp 1621261055
transform 1 0 16992 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_173
timestamp 1621261055
transform 1 0 17760 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_181
timestamp 1621261055
transform 1 0 18528 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_189
timestamp 1621261055
transform 1 0 19296 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_702
timestamp 1621261055
transform 1 0 19680 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_194
timestamp 1621261055
transform 1 0 19776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_202
timestamp 1621261055
transform 1 0 20544 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_210
timestamp 1621261055
transform 1 0 21312 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_218
timestamp 1621261055
transform 1 0 22080 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_226
timestamp 1621261055
transform 1 0 22848 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_703
timestamp 1621261055
transform 1 0 24960 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_234
timestamp 1621261055
transform 1 0 23616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_242
timestamp 1621261055
transform 1 0 24384 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_246
timestamp 1621261055
transform 1 0 24768 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_249
timestamp 1621261055
transform 1 0 25056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_257
timestamp 1621261055
transform 1 0 25824 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_265
timestamp 1621261055
transform 1 0 26592 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_273
timestamp 1621261055
transform 1 0 27360 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_281
timestamp 1621261055
transform 1 0 28128 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_289
timestamp 1621261055
transform 1 0 28896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_704
timestamp 1621261055
transform 1 0 30240 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_297
timestamp 1621261055
transform 1 0 29664 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_301
timestamp 1621261055
transform 1 0 30048 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_304
timestamp 1621261055
transform 1 0 30336 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_312
timestamp 1621261055
transform 1 0 31104 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_320
timestamp 1621261055
transform 1 0 31872 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_328
timestamp 1621261055
transform 1 0 32640 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_336
timestamp 1621261055
transform 1 0 33408 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_344
timestamp 1621261055
transform 1 0 34176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_352
timestamp 1621261055
transform 1 0 34944 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_356
timestamp 1621261055
transform 1 0 35328 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_705
timestamp 1621261055
transform 1 0 35520 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_359
timestamp 1621261055
transform 1 0 35616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_367
timestamp 1621261055
transform 1 0 36384 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_375
timestamp 1621261055
transform 1 0 37152 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_383
timestamp 1621261055
transform 1 0 37920 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_391
timestamp 1621261055
transform 1 0 38688 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_399
timestamp 1621261055
transform 1 0 39456 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _143_
timestamp 1621261055
transform 1 0 40128 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_706
timestamp 1621261055
transform 1 0 40800 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_196
timestamp 1621261055
transform 1 0 39936 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_50_403
timestamp 1621261055
transform 1 0 39840 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_409
timestamp 1621261055
transform 1 0 40416 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_414
timestamp 1621261055
transform 1 0 40896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_422
timestamp 1621261055
transform 1 0 41664 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_430
timestamp 1621261055
transform 1 0 42432 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_438
timestamp 1621261055
transform 1 0 43200 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_446
timestamp 1621261055
transform 1 0 43968 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_454
timestamp 1621261055
transform 1 0 44736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_462
timestamp 1621261055
transform 1 0 45504 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _189_
timestamp 1621261055
transform -1 0 46848 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_707
timestamp 1621261055
transform 1 0 46080 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_236
timestamp 1621261055
transform -1 0 46560 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_466
timestamp 1621261055
transform 1 0 45888 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_469
timestamp 1621261055
transform 1 0 46176 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_476
timestamp 1621261055
transform 1 0 46848 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_484
timestamp 1621261055
transform 1 0 47616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_492
timestamp 1621261055
transform 1 0 48384 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_500
timestamp 1621261055
transform 1 0 49152 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_708
timestamp 1621261055
transform 1 0 51360 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_508
timestamp 1621261055
transform 1 0 49920 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_516
timestamp 1621261055
transform 1 0 50688 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_520
timestamp 1621261055
transform 1 0 51072 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_50_522
timestamp 1621261055
transform 1 0 51264 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_524
timestamp 1621261055
transform 1 0 51456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_532
timestamp 1621261055
transform 1 0 52224 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_540
timestamp 1621261055
transform 1 0 52992 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_548
timestamp 1621261055
transform 1 0 53760 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_556
timestamp 1621261055
transform 1 0 54528 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_564
timestamp 1621261055
transform 1 0 55296 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_709
timestamp 1621261055
transform 1 0 56640 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_572
timestamp 1621261055
transform 1 0 56064 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_576
timestamp 1621261055
transform 1 0 56448 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_579
timestamp 1621261055
transform 1 0 56736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_587
timestamp 1621261055
transform 1 0 57504 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_101
timestamp 1621261055
transform -1 0 58848 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_595
timestamp 1621261055
transform 1 0 58272 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_102
timestamp 1621261055
transform 1 0 1152 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_4
timestamp 1621261055
transform 1 0 1536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_12
timestamp 1621261055
transform 1 0 2304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_20
timestamp 1621261055
transform 1 0 3072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_28
timestamp 1621261055
transform 1 0 3840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_36
timestamp 1621261055
transform 1 0 4608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_710
timestamp 1621261055
transform 1 0 6432 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_44
timestamp 1621261055
transform 1 0 5376 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_52
timestamp 1621261055
transform 1 0 6144 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_54
timestamp 1621261055
transform 1 0 6336 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_56
timestamp 1621261055
transform 1 0 6528 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_64
timestamp 1621261055
transform 1 0 7296 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_72
timestamp 1621261055
transform 1 0 8064 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_80
timestamp 1621261055
transform 1 0 8832 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_88
timestamp 1621261055
transform 1 0 9600 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_96
timestamp 1621261055
transform 1 0 10368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_104
timestamp 1621261055
transform 1 0 11136 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_711
timestamp 1621261055
transform 1 0 11712 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_108
timestamp 1621261055
transform 1 0 11520 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_111
timestamp 1621261055
transform 1 0 11808 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_119
timestamp 1621261055
transform 1 0 12576 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_127
timestamp 1621261055
transform 1 0 13344 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_135
timestamp 1621261055
transform 1 0 14112 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_143
timestamp 1621261055
transform 1 0 14880 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_712
timestamp 1621261055
transform 1 0 16992 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_151
timestamp 1621261055
transform 1 0 15648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_159
timestamp 1621261055
transform 1 0 16416 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_163
timestamp 1621261055
transform 1 0 16800 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_166
timestamp 1621261055
transform 1 0 17088 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_174
timestamp 1621261055
transform 1 0 17856 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_182
timestamp 1621261055
transform 1 0 18624 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_190
timestamp 1621261055
transform 1 0 19392 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_198
timestamp 1621261055
transform 1 0 20160 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_206
timestamp 1621261055
transform 1 0 20928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_713
timestamp 1621261055
transform 1 0 22272 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_214
timestamp 1621261055
transform 1 0 21696 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_218
timestamp 1621261055
transform 1 0 22080 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_221
timestamp 1621261055
transform 1 0 22368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_229
timestamp 1621261055
transform 1 0 23136 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_237
timestamp 1621261055
transform 1 0 23904 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_245
timestamp 1621261055
transform 1 0 24672 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_253
timestamp 1621261055
transform 1 0 25440 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_261
timestamp 1621261055
transform 1 0 26208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_269
timestamp 1621261055
transform 1 0 26976 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_273
timestamp 1621261055
transform 1 0 27360 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_714
timestamp 1621261055
transform 1 0 27552 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_276
timestamp 1621261055
transform 1 0 27648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_284
timestamp 1621261055
transform 1 0 28416 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_292
timestamp 1621261055
transform 1 0 29184 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_300
timestamp 1621261055
transform 1 0 29952 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_308
timestamp 1621261055
transform 1 0 30720 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_715
timestamp 1621261055
transform 1 0 32832 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_316
timestamp 1621261055
transform 1 0 31488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_324
timestamp 1621261055
transform 1 0 32256 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_328
timestamp 1621261055
transform 1 0 32640 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_331
timestamp 1621261055
transform 1 0 32928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_339
timestamp 1621261055
transform 1 0 33696 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_347
timestamp 1621261055
transform 1 0 34464 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_355
timestamp 1621261055
transform 1 0 35232 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_363
timestamp 1621261055
transform 1 0 36000 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_371
timestamp 1621261055
transform 1 0 36768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_716
timestamp 1621261055
transform 1 0 38112 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_379
timestamp 1621261055
transform 1 0 37536 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_383
timestamp 1621261055
transform 1 0 37920 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_386
timestamp 1621261055
transform 1 0 38208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_394
timestamp 1621261055
transform 1 0 38976 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_402
timestamp 1621261055
transform 1 0 39744 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_410
timestamp 1621261055
transform 1 0 40512 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_418
timestamp 1621261055
transform 1 0 41280 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_717
timestamp 1621261055
transform 1 0 43392 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_426
timestamp 1621261055
transform 1 0 42048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_434
timestamp 1621261055
transform 1 0 42816 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_438
timestamp 1621261055
transform 1 0 43200 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_51_441
timestamp 1621261055
transform 1 0 43488 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _062_
timestamp 1621261055
transform -1 0 44448 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_146
timestamp 1621261055
transform -1 0 44160 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_445
timestamp 1621261055
transform 1 0 43872 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_451
timestamp 1621261055
transform 1 0 44448 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_459
timestamp 1621261055
transform 1 0 45216 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_467
timestamp 1621261055
transform 1 0 45984 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_475
timestamp 1621261055
transform 1 0 46752 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_483
timestamp 1621261055
transform 1 0 47520 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_718
timestamp 1621261055
transform 1 0 48672 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_491
timestamp 1621261055
transform 1 0 48288 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_496
timestamp 1621261055
transform 1 0 48768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_504
timestamp 1621261055
transform 1 0 49536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_512
timestamp 1621261055
transform 1 0 50304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_520
timestamp 1621261055
transform 1 0 51072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_528
timestamp 1621261055
transform 1 0 51840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_536
timestamp 1621261055
transform 1 0 52608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_544
timestamp 1621261055
transform 1 0 53376 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_719
timestamp 1621261055
transform 1 0 53952 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_548
timestamp 1621261055
transform 1 0 53760 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_551
timestamp 1621261055
transform 1 0 54048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_559
timestamp 1621261055
transform 1 0 54816 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_567
timestamp 1621261055
transform 1 0 55584 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_575
timestamp 1621261055
transform 1 0 56352 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_583
timestamp 1621261055
transform 1 0 57120 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_103
timestamp 1621261055
transform -1 0 58848 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_51_591
timestamp 1621261055
transform 1 0 57888 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_595
timestamp 1621261055
transform 1 0 58272 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_104
timestamp 1621261055
transform 1 0 1152 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_52_4
timestamp 1621261055
transform 1 0 1536 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_12
timestamp 1621261055
transform 1 0 2304 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_20
timestamp 1621261055
transform 1 0 3072 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_720
timestamp 1621261055
transform 1 0 3840 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_29
timestamp 1621261055
transform 1 0 3936 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_37
timestamp 1621261055
transform 1 0 4704 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_45
timestamp 1621261055
transform 1 0 5472 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_53
timestamp 1621261055
transform 1 0 6240 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_61
timestamp 1621261055
transform 1 0 7008 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_721
timestamp 1621261055
transform 1 0 9120 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_69
timestamp 1621261055
transform 1 0 7776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_77
timestamp 1621261055
transform 1 0 8544 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_81
timestamp 1621261055
transform 1 0 8928 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_84
timestamp 1621261055
transform 1 0 9216 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _060_
timestamp 1621261055
transform 1 0 11040 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_95
timestamp 1621261055
transform 1 0 10848 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_92
timestamp 1621261055
transform 1 0 9984 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_52_100
timestamp 1621261055
transform 1 0 10752 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_106
timestamp 1621261055
transform 1 0 11328 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_114
timestamp 1621261055
transform 1 0 12096 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_122
timestamp 1621261055
transform 1 0 12864 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_722
timestamp 1621261055
transform 1 0 14400 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_130
timestamp 1621261055
transform 1 0 13632 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_139
timestamp 1621261055
transform 1 0 14496 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_147
timestamp 1621261055
transform 1 0 15264 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_155
timestamp 1621261055
transform 1 0 16032 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_163
timestamp 1621261055
transform 1 0 16800 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_171
timestamp 1621261055
transform 1 0 17568 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_179
timestamp 1621261055
transform 1 0 18336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_187
timestamp 1621261055
transform 1 0 19104 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_723
timestamp 1621261055
transform 1 0 19680 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_191
timestamp 1621261055
transform 1 0 19488 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_194
timestamp 1621261055
transform 1 0 19776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_202
timestamp 1621261055
transform 1 0 20544 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_210
timestamp 1621261055
transform 1 0 21312 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_218
timestamp 1621261055
transform 1 0 22080 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_226
timestamp 1621261055
transform 1 0 22848 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_724
timestamp 1621261055
transform 1 0 24960 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_234
timestamp 1621261055
transform 1 0 23616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_242
timestamp 1621261055
transform 1 0 24384 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_246
timestamp 1621261055
transform 1 0 24768 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_249
timestamp 1621261055
transform 1 0 25056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_257
timestamp 1621261055
transform 1 0 25824 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_265
timestamp 1621261055
transform 1 0 26592 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_273
timestamp 1621261055
transform 1 0 27360 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_281
timestamp 1621261055
transform 1 0 28128 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_289
timestamp 1621261055
transform 1 0 28896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_725
timestamp 1621261055
transform 1 0 30240 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_297
timestamp 1621261055
transform 1 0 29664 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_301
timestamp 1621261055
transform 1 0 30048 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_304
timestamp 1621261055
transform 1 0 30336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_312
timestamp 1621261055
transform 1 0 31104 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _156_
timestamp 1621261055
transform 1 0 33024 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_99
timestamp 1621261055
transform 1 0 32832 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_320
timestamp 1621261055
transform 1 0 31872 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_328
timestamp 1621261055
transform 1 0 32640 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_335
timestamp 1621261055
transform 1 0 33312 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_343
timestamp 1621261055
transform 1 0 34080 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_351
timestamp 1621261055
transform 1 0 34848 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_355
timestamp 1621261055
transform 1 0 35232 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_357
timestamp 1621261055
transform 1 0 35424 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_726
timestamp 1621261055
transform 1 0 35520 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_359
timestamp 1621261055
transform 1 0 35616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_367
timestamp 1621261055
transform 1 0 36384 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_375
timestamp 1621261055
transform 1 0 37152 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_383
timestamp 1621261055
transform 1 0 37920 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_391
timestamp 1621261055
transform 1 0 38688 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_399
timestamp 1621261055
transform 1 0 39456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_727
timestamp 1621261055
transform 1 0 40800 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_407
timestamp 1621261055
transform 1 0 40224 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_411
timestamp 1621261055
transform 1 0 40608 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_414
timestamp 1621261055
transform 1 0 40896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_422
timestamp 1621261055
transform 1 0 41664 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_430
timestamp 1621261055
transform 1 0 42432 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_438
timestamp 1621261055
transform 1 0 43200 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_446
timestamp 1621261055
transform 1 0 43968 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_454
timestamp 1621261055
transform 1 0 44736 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_462
timestamp 1621261055
transform 1 0 45504 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_728
timestamp 1621261055
transform 1 0 46080 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_466
timestamp 1621261055
transform 1 0 45888 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_469
timestamp 1621261055
transform 1 0 46176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_477
timestamp 1621261055
transform 1 0 46944 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_485
timestamp 1621261055
transform 1 0 47712 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_493
timestamp 1621261055
transform 1 0 48480 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_501
timestamp 1621261055
transform 1 0 49248 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_729
timestamp 1621261055
transform 1 0 51360 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_509
timestamp 1621261055
transform 1 0 50016 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_517
timestamp 1621261055
transform 1 0 50784 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_521
timestamp 1621261055
transform 1 0 51168 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_524
timestamp 1621261055
transform 1 0 51456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_532
timestamp 1621261055
transform 1 0 52224 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_540
timestamp 1621261055
transform 1 0 52992 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_548
timestamp 1621261055
transform 1 0 53760 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_556
timestamp 1621261055
transform 1 0 54528 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_564
timestamp 1621261055
transform 1 0 55296 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _170_
timestamp 1621261055
transform 1 0 57120 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_730
timestamp 1621261055
transform 1 0 56640 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_572
timestamp 1621261055
transform 1 0 56064 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_576
timestamp 1621261055
transform 1 0 56448 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_52_579
timestamp 1621261055
transform 1 0 56736 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_52_586
timestamp 1621261055
transform 1 0 57408 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_105
timestamp 1621261055
transform -1 0 58848 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_594
timestamp 1621261055
transform 1 0 58176 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_596
timestamp 1621261055
transform 1 0 58368 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_106
timestamp 1621261055
transform 1 0 1152 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_4
timestamp 1621261055
transform 1 0 1536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_12
timestamp 1621261055
transform 1 0 2304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_20
timestamp 1621261055
transform 1 0 3072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_28
timestamp 1621261055
transform 1 0 3840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_36
timestamp 1621261055
transform 1 0 4608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_731
timestamp 1621261055
transform 1 0 6432 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_44
timestamp 1621261055
transform 1 0 5376 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_52
timestamp 1621261055
transform 1 0 6144 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_54
timestamp 1621261055
transform 1 0 6336 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_56
timestamp 1621261055
transform 1 0 6528 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_64
timestamp 1621261055
transform 1 0 7296 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_72
timestamp 1621261055
transform 1 0 8064 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_80
timestamp 1621261055
transform 1 0 8832 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_88
timestamp 1621261055
transform 1 0 9600 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_96
timestamp 1621261055
transform 1 0 10368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_104
timestamp 1621261055
transform 1 0 11136 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_732
timestamp 1621261055
transform 1 0 11712 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_108
timestamp 1621261055
transform 1 0 11520 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_111
timestamp 1621261055
transform 1 0 11808 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_119
timestamp 1621261055
transform 1 0 12576 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _197_
timestamp 1621261055
transform -1 0 14688 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_214
timestamp 1621261055
transform -1 0 14400 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_127
timestamp 1621261055
transform 1 0 13344 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_53_135
timestamp 1621261055
transform 1 0 14112 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_141
timestamp 1621261055
transform 1 0 14688 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_733
timestamp 1621261055
transform 1 0 16992 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_149
timestamp 1621261055
transform 1 0 15456 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_157
timestamp 1621261055
transform 1 0 16224 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_166
timestamp 1621261055
transform 1 0 17088 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _196_
timestamp 1621261055
transform -1 0 18528 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_212
timestamp 1621261055
transform -1 0 18240 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_174
timestamp 1621261055
transform 1 0 17856 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_181
timestamp 1621261055
transform 1 0 18528 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_189
timestamp 1621261055
transform 1 0 19296 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_197
timestamp 1621261055
transform 1 0 20064 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_205
timestamp 1621261055
transform 1 0 20832 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_734
timestamp 1621261055
transform 1 0 22272 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_213
timestamp 1621261055
transform 1 0 21600 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_217
timestamp 1621261055
transform 1 0 21984 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_219
timestamp 1621261055
transform 1 0 22176 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_221
timestamp 1621261055
transform 1 0 22368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_229
timestamp 1621261055
transform 1 0 23136 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _030_
timestamp 1621261055
transform 1 0 23712 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_233
timestamp 1621261055
transform 1 0 23520 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_238
timestamp 1621261055
transform 1 0 24000 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_246
timestamp 1621261055
transform 1 0 24768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_254
timestamp 1621261055
transform 1 0 25536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_262
timestamp 1621261055
transform 1 0 26304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_270
timestamp 1621261055
transform 1 0 27072 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_735
timestamp 1621261055
transform 1 0 27552 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_53_274
timestamp 1621261055
transform 1 0 27456 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_276
timestamp 1621261055
transform 1 0 27648 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_284
timestamp 1621261055
transform 1 0 28416 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_292
timestamp 1621261055
transform 1 0 29184 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _022_
timestamp 1621261055
transform 1 0 29856 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _031_
timestamp 1621261055
transform 1 0 30528 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_296
timestamp 1621261055
transform 1 0 29568 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_298
timestamp 1621261055
transform 1 0 29760 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_302
timestamp 1621261055
transform 1 0 30144 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_309
timestamp 1621261055
transform 1 0 30816 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_736
timestamp 1621261055
transform 1 0 32832 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_317
timestamp 1621261055
transform 1 0 31584 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_325
timestamp 1621261055
transform 1 0 32352 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_53_329
timestamp 1621261055
transform 1 0 32736 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_331
timestamp 1621261055
transform 1 0 32928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_339
timestamp 1621261055
transform 1 0 33696 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_347
timestamp 1621261055
transform 1 0 34464 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_355
timestamp 1621261055
transform 1 0 35232 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_363
timestamp 1621261055
transform 1 0 36000 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_371
timestamp 1621261055
transform 1 0 36768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _106_
timestamp 1621261055
transform -1 0 38976 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_737
timestamp 1621261055
transform 1 0 38112 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_168
timestamp 1621261055
transform -1 0 38688 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_53_379
timestamp 1621261055
transform 1 0 37536 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_383
timestamp 1621261055
transform 1 0 37920 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_386
timestamp 1621261055
transform 1 0 38208 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_388
timestamp 1621261055
transform 1 0 38400 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_394
timestamp 1621261055
transform 1 0 38976 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_402
timestamp 1621261055
transform 1 0 39744 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_410
timestamp 1621261055
transform 1 0 40512 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_418
timestamp 1621261055
transform 1 0 41280 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_738
timestamp 1621261055
transform 1 0 43392 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_426
timestamp 1621261055
transform 1 0 42048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_434
timestamp 1621261055
transform 1 0 42816 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_438
timestamp 1621261055
transform 1 0 43200 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_441
timestamp 1621261055
transform 1 0 43488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_449
timestamp 1621261055
transform 1 0 44256 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_457
timestamp 1621261055
transform 1 0 45024 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_465
timestamp 1621261055
transform 1 0 45792 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_473
timestamp 1621261055
transform 1 0 46560 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_481
timestamp 1621261055
transform 1 0 47328 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_739
timestamp 1621261055
transform 1 0 48672 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_489
timestamp 1621261055
transform 1 0 48096 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_493
timestamp 1621261055
transform 1 0 48480 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_496
timestamp 1621261055
transform 1 0 48768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_504
timestamp 1621261055
transform 1 0 49536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_512
timestamp 1621261055
transform 1 0 50304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_520
timestamp 1621261055
transform 1 0 51072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_528
timestamp 1621261055
transform 1 0 51840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_536
timestamp 1621261055
transform 1 0 52608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_544
timestamp 1621261055
transform 1 0 53376 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_740
timestamp 1621261055
transform 1 0 53952 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_548
timestamp 1621261055
transform 1 0 53760 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_551
timestamp 1621261055
transform 1 0 54048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_559
timestamp 1621261055
transform 1 0 54816 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_567
timestamp 1621261055
transform 1 0 55584 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_575
timestamp 1621261055
transform 1 0 56352 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_583
timestamp 1621261055
transform 1 0 57120 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_107
timestamp 1621261055
transform -1 0 58848 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_53_591
timestamp 1621261055
transform 1 0 57888 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_595
timestamp 1621261055
transform 1 0 58272 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_108
timestamp 1621261055
transform 1 0 1152 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_110
timestamp 1621261055
transform 1 0 1152 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_4
timestamp 1621261055
transform 1 0 1536 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_12
timestamp 1621261055
transform 1 0 2304 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_20
timestamp 1621261055
transform 1 0 3072 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_4
timestamp 1621261055
transform 1 0 1536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_12
timestamp 1621261055
transform 1 0 2304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_20
timestamp 1621261055
transform 1 0 3072 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_741
timestamp 1621261055
transform 1 0 3840 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_29
timestamp 1621261055
transform 1 0 3936 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_37
timestamp 1621261055
transform 1 0 4704 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_28
timestamp 1621261055
transform 1 0 3840 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_36
timestamp 1621261055
transform 1 0 4608 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_44
timestamp 1621261055
transform 1 0 5376 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_45
timestamp 1621261055
transform 1 0 5472 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_56
timestamp 1621261055
transform 1 0 6528 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_55_54
timestamp 1621261055
transform 1 0 6336 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_52
timestamp 1621261055
transform 1 0 6144 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_53
timestamp 1621261055
transform 1 0 6240 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_165
timestamp 1621261055
transform 1 0 6720 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_752
timestamp 1621261055
transform 1 0 6432 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_63
timestamp 1621261055
transform 1 0 7200 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_61
timestamp 1621261055
transform 1 0 7008 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _105_
timestamp 1621261055
transform 1 0 6912 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_742
timestamp 1621261055
transform 1 0 9120 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_69
timestamp 1621261055
transform 1 0 7776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_77
timestamp 1621261055
transform 1 0 8544 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_81
timestamp 1621261055
transform 1 0 8928 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_84
timestamp 1621261055
transform 1 0 9216 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_71
timestamp 1621261055
transform 1 0 7968 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_79
timestamp 1621261055
transform 1 0 8736 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_92
timestamp 1621261055
transform 1 0 9984 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_100
timestamp 1621261055
transform 1 0 10752 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_87
timestamp 1621261055
transform 1 0 9504 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_95
timestamp 1621261055
transform 1 0 10272 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_103
timestamp 1621261055
transform 1 0 11040 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_753
timestamp 1621261055
transform 1 0 11712 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_108
timestamp 1621261055
transform 1 0 11520 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_116
timestamp 1621261055
transform 1 0 12288 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_124
timestamp 1621261055
transform 1 0 13056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_107
timestamp 1621261055
transform 1 0 11424 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_55_109
timestamp 1621261055
transform 1 0 11616 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_111
timestamp 1621261055
transform 1 0 11808 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_119
timestamp 1621261055
transform 1 0 12576 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _045_
timestamp 1621261055
transform 1 0 15072 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_743
timestamp 1621261055
transform 1 0 14400 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_132
timestamp 1621261055
transform 1 0 13824 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_136
timestamp 1621261055
transform 1 0 14208 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_139
timestamp 1621261055
transform 1 0 14496 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_143
timestamp 1621261055
transform 1 0 14880 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_127
timestamp 1621261055
transform 1 0 13344 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_135
timestamp 1621261055
transform 1 0 14112 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_143
timestamp 1621261055
transform 1 0 14880 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_754
timestamp 1621261055
transform 1 0 16992 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_148
timestamp 1621261055
transform 1 0 15360 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_156
timestamp 1621261055
transform 1 0 16128 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_164
timestamp 1621261055
transform 1 0 16896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_151
timestamp 1621261055
transform 1 0 15648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_159
timestamp 1621261055
transform 1 0 16416 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_163
timestamp 1621261055
transform 1 0 16800 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_166
timestamp 1621261055
transform 1 0 17088 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_172
timestamp 1621261055
transform 1 0 17664 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_180
timestamp 1621261055
transform 1 0 18432 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_188
timestamp 1621261055
transform 1 0 19200 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_174
timestamp 1621261055
transform 1 0 17856 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_182
timestamp 1621261055
transform 1 0 18624 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_744
timestamp 1621261055
transform 1 0 19680 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_54_192
timestamp 1621261055
transform 1 0 19584 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_194
timestamp 1621261055
transform 1 0 19776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_202
timestamp 1621261055
transform 1 0 20544 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_210
timestamp 1621261055
transform 1 0 21312 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_190
timestamp 1621261055
transform 1 0 19392 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_198
timestamp 1621261055
transform 1 0 20160 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_206
timestamp 1621261055
transform 1 0 20928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_755
timestamp 1621261055
transform 1 0 22272 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_218
timestamp 1621261055
transform 1 0 22080 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_226
timestamp 1621261055
transform 1 0 22848 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_214
timestamp 1621261055
transform 1 0 21696 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_218
timestamp 1621261055
transform 1 0 22080 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_221
timestamp 1621261055
transform 1 0 22368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_229
timestamp 1621261055
transform 1 0 23136 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_55_231
timestamp 1621261055
transform 1 0 23328 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _028_
timestamp 1621261055
transform 1 0 23424 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_745
timestamp 1621261055
transform 1 0 24960 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_234
timestamp 1621261055
transform 1 0 23616 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_242
timestamp 1621261055
transform 1 0 24384 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_246
timestamp 1621261055
transform 1 0 24768 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_249
timestamp 1621261055
transform 1 0 25056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_235
timestamp 1621261055
transform 1 0 23712 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_243
timestamp 1621261055
transform 1 0 24480 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_251
timestamp 1621261055
transform 1 0 25248 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_257
timestamp 1621261055
transform 1 0 25824 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_265
timestamp 1621261055
transform 1 0 26592 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_273
timestamp 1621261055
transform 1 0 27360 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_259
timestamp 1621261055
transform 1 0 26016 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_267
timestamp 1621261055
transform 1 0 26784 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_756
timestamp 1621261055
transform 1 0 27552 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_281
timestamp 1621261055
transform 1 0 28128 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_289
timestamp 1621261055
transform 1 0 28896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_276
timestamp 1621261055
transform 1 0 27648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_284
timestamp 1621261055
transform 1 0 28416 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_292
timestamp 1621261055
transform 1 0 29184 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_746
timestamp 1621261055
transform 1 0 30240 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_297
timestamp 1621261055
transform 1 0 29664 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_301
timestamp 1621261055
transform 1 0 30048 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_304
timestamp 1621261055
transform 1 0 30336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_312
timestamp 1621261055
transform 1 0 31104 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_300
timestamp 1621261055
transform 1 0 29952 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_308
timestamp 1621261055
transform 1 0 30720 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_757
timestamp 1621261055
transform 1 0 32832 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_320
timestamp 1621261055
transform 1 0 31872 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_328
timestamp 1621261055
transform 1 0 32640 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_336
timestamp 1621261055
transform 1 0 33408 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_316
timestamp 1621261055
transform 1 0 31488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_324
timestamp 1621261055
transform 1 0 32256 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_328
timestamp 1621261055
transform 1 0 32640 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_331
timestamp 1621261055
transform 1 0 32928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_344
timestamp 1621261055
transform 1 0 34176 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_352
timestamp 1621261055
transform 1 0 34944 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_356
timestamp 1621261055
transform 1 0 35328 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_339
timestamp 1621261055
transform 1 0 33696 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_347
timestamp 1621261055
transform 1 0 34464 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_355
timestamp 1621261055
transform 1 0 35232 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_747
timestamp 1621261055
transform 1 0 35520 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_359
timestamp 1621261055
transform 1 0 35616 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_367
timestamp 1621261055
transform 1 0 36384 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_375
timestamp 1621261055
transform 1 0 37152 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_363
timestamp 1621261055
transform 1 0 36000 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_371
timestamp 1621261055
transform 1 0 36768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_758
timestamp 1621261055
transform 1 0 38112 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_383
timestamp 1621261055
transform 1 0 37920 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_391
timestamp 1621261055
transform 1 0 38688 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_399
timestamp 1621261055
transform 1 0 39456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_379
timestamp 1621261055
transform 1 0 37536 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_383
timestamp 1621261055
transform 1 0 37920 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_386
timestamp 1621261055
transform 1 0 38208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_394
timestamp 1621261055
transform 1 0 38976 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_748
timestamp 1621261055
transform 1 0 40800 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_407
timestamp 1621261055
transform 1 0 40224 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_411
timestamp 1621261055
transform 1 0 40608 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_414
timestamp 1621261055
transform 1 0 40896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_402
timestamp 1621261055
transform 1 0 39744 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_410
timestamp 1621261055
transform 1 0 40512 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_418
timestamp 1621261055
transform 1 0 41280 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_759
timestamp 1621261055
transform 1 0 43392 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_422
timestamp 1621261055
transform 1 0 41664 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_430
timestamp 1621261055
transform 1 0 42432 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_438
timestamp 1621261055
transform 1 0 43200 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_426
timestamp 1621261055
transform 1 0 42048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_434
timestamp 1621261055
transform 1 0 42816 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_438
timestamp 1621261055
transform 1 0 43200 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_441
timestamp 1621261055
transform 1 0 43488 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _162_
timestamp 1621261055
transform 1 0 43872 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_107
timestamp 1621261055
transform 1 0 43680 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_446
timestamp 1621261055
transform 1 0 43968 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_454
timestamp 1621261055
transform 1 0 44736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_462
timestamp 1621261055
transform 1 0 45504 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_448
timestamp 1621261055
transform 1 0 44160 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_456
timestamp 1621261055
transform 1 0 44928 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_460
timestamp 1621261055
transform 1 0 45312 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_55_462
timestamp 1621261055
transform 1 0 45504 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _032_
timestamp 1621261055
transform 1 0 45600 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_749
timestamp 1621261055
transform 1 0 46080 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_466
timestamp 1621261055
transform 1 0 45888 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_469
timestamp 1621261055
transform 1 0 46176 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_477
timestamp 1621261055
transform 1 0 46944 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_466
timestamp 1621261055
transform 1 0 45888 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_474
timestamp 1621261055
transform 1 0 46656 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_482
timestamp 1621261055
transform 1 0 47424 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_490
timestamp 1621261055
transform 1 0 48192 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_491
timestamp 1621261055
transform 1 0 48288 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_485
timestamp 1621261055
transform 1 0 47712 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_136
timestamp 1621261055
transform -1 0 48000 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _076_
timestamp 1621261055
transform -1 0 48288 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_500
timestamp 1621261055
transform 1 0 49152 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_55_496
timestamp 1621261055
transform 1 0 48768 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_55_494
timestamp 1621261055
transform 1 0 48576 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_499
timestamp 1621261055
transform 1 0 49056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_760
timestamp 1621261055
transform 1 0 48672 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_150
timestamp 1621261055
transform -1 0 49536 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _097_
timestamp 1621261055
transform -1 0 49824 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_750
timestamp 1621261055
transform 1 0 51360 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_507
timestamp 1621261055
transform 1 0 49824 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_515
timestamp 1621261055
transform 1 0 50592 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_524
timestamp 1621261055
transform 1 0 51456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_507
timestamp 1621261055
transform 1 0 49824 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_515
timestamp 1621261055
transform 1 0 50592 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_523
timestamp 1621261055
transform 1 0 51360 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_532
timestamp 1621261055
transform 1 0 52224 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_540
timestamp 1621261055
transform 1 0 52992 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_531
timestamp 1621261055
transform 1 0 52128 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_539
timestamp 1621261055
transform 1 0 52896 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_761
timestamp 1621261055
transform 1 0 53952 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_548
timestamp 1621261055
transform 1 0 53760 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_556
timestamp 1621261055
transform 1 0 54528 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_564
timestamp 1621261055
transform 1 0 55296 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_547
timestamp 1621261055
transform 1 0 53664 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_55_549
timestamp 1621261055
transform 1 0 53856 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_551
timestamp 1621261055
transform 1 0 54048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_559
timestamp 1621261055
transform 1 0 54816 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_567
timestamp 1621261055
transform 1 0 55584 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _171_
timestamp 1621261055
transform -1 0 57408 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_751
timestamp 1621261055
transform 1 0 56640 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_118
timestamp 1621261055
transform -1 0 57120 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_572
timestamp 1621261055
transform 1 0 56064 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_576
timestamp 1621261055
transform 1 0 56448 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_579
timestamp 1621261055
transform 1 0 56736 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_586
timestamp 1621261055
transform 1 0 57408 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_575
timestamp 1621261055
transform 1 0 56352 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_583
timestamp 1621261055
transform 1 0 57120 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_109
timestamp 1621261055
transform -1 0 58848 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_111
timestamp 1621261055
transform -1 0 58848 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_594
timestamp 1621261055
transform 1 0 58176 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_54_596
timestamp 1621261055
transform 1 0 58368 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_55_591
timestamp 1621261055
transform 1 0 57888 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_595
timestamp 1621261055
transform 1 0 58272 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_112
timestamp 1621261055
transform 1 0 1152 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_56_4
timestamp 1621261055
transform 1 0 1536 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_12
timestamp 1621261055
transform 1 0 2304 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_20
timestamp 1621261055
transform 1 0 3072 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_762
timestamp 1621261055
transform 1 0 3840 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_29
timestamp 1621261055
transform 1 0 3936 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_37
timestamp 1621261055
transform 1 0 4704 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_45
timestamp 1621261055
transform 1 0 5472 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_53
timestamp 1621261055
transform 1 0 6240 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_61
timestamp 1621261055
transform 1 0 7008 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_763
timestamp 1621261055
transform 1 0 9120 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_69
timestamp 1621261055
transform 1 0 7776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_77
timestamp 1621261055
transform 1 0 8544 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_81
timestamp 1621261055
transform 1 0 8928 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_84
timestamp 1621261055
transform 1 0 9216 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_92
timestamp 1621261055
transform 1 0 9984 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_100
timestamp 1621261055
transform 1 0 10752 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_108
timestamp 1621261055
transform 1 0 11520 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_116
timestamp 1621261055
transform 1 0 12288 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_124
timestamp 1621261055
transform 1 0 13056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_764
timestamp 1621261055
transform 1 0 14400 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_132
timestamp 1621261055
transform 1 0 13824 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_136
timestamp 1621261055
transform 1 0 14208 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_139
timestamp 1621261055
transform 1 0 14496 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_147
timestamp 1621261055
transform 1 0 15264 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_155
timestamp 1621261055
transform 1 0 16032 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_163
timestamp 1621261055
transform 1 0 16800 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_171
timestamp 1621261055
transform 1 0 17568 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_179
timestamp 1621261055
transform 1 0 18336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_187
timestamp 1621261055
transform 1 0 19104 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_765
timestamp 1621261055
transform 1 0 19680 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_191
timestamp 1621261055
transform 1 0 19488 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_194
timestamp 1621261055
transform 1 0 19776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_202
timestamp 1621261055
transform 1 0 20544 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_210
timestamp 1621261055
transform 1 0 21312 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_218
timestamp 1621261055
transform 1 0 22080 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_226
timestamp 1621261055
transform 1 0 22848 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_766
timestamp 1621261055
transform 1 0 24960 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_234
timestamp 1621261055
transform 1 0 23616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_242
timestamp 1621261055
transform 1 0 24384 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_246
timestamp 1621261055
transform 1 0 24768 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_249
timestamp 1621261055
transform 1 0 25056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_257
timestamp 1621261055
transform 1 0 25824 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_265
timestamp 1621261055
transform 1 0 26592 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_273
timestamp 1621261055
transform 1 0 27360 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_281
timestamp 1621261055
transform 1 0 28128 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_289
timestamp 1621261055
transform 1 0 28896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_767
timestamp 1621261055
transform 1 0 30240 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_297
timestamp 1621261055
transform 1 0 29664 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_301
timestamp 1621261055
transform 1 0 30048 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_304
timestamp 1621261055
transform 1 0 30336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_312
timestamp 1621261055
transform 1 0 31104 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_320
timestamp 1621261055
transform 1 0 31872 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_328
timestamp 1621261055
transform 1 0 32640 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_336
timestamp 1621261055
transform 1 0 33408 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_344
timestamp 1621261055
transform 1 0 34176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_352
timestamp 1621261055
transform 1 0 34944 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_356
timestamp 1621261055
transform 1 0 35328 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_768
timestamp 1621261055
transform 1 0 35520 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_359
timestamp 1621261055
transform 1 0 35616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_367
timestamp 1621261055
transform 1 0 36384 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_375
timestamp 1621261055
transform 1 0 37152 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_383
timestamp 1621261055
transform 1 0 37920 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_391
timestamp 1621261055
transform 1 0 38688 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_399
timestamp 1621261055
transform 1 0 39456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_769
timestamp 1621261055
transform 1 0 40800 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_407
timestamp 1621261055
transform 1 0 40224 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_411
timestamp 1621261055
transform 1 0 40608 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_414
timestamp 1621261055
transform 1 0 40896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_422
timestamp 1621261055
transform 1 0 41664 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_430
timestamp 1621261055
transform 1 0 42432 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_438
timestamp 1621261055
transform 1 0 43200 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _098_
timestamp 1621261055
transform -1 0 45504 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_152
timestamp 1621261055
transform -1 0 45216 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_446
timestamp 1621261055
transform 1 0 43968 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_454
timestamp 1621261055
transform 1 0 44736 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_56_456
timestamp 1621261055
transform 1 0 44928 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_462
timestamp 1621261055
transform 1 0 45504 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_770
timestamp 1621261055
transform 1 0 46080 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_466
timestamp 1621261055
transform 1 0 45888 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_469
timestamp 1621261055
transform 1 0 46176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_477
timestamp 1621261055
transform 1 0 46944 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_485
timestamp 1621261055
transform 1 0 47712 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_493
timestamp 1621261055
transform 1 0 48480 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_501
timestamp 1621261055
transform 1 0 49248 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_771
timestamp 1621261055
transform 1 0 51360 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_509
timestamp 1621261055
transform 1 0 50016 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_517
timestamp 1621261055
transform 1 0 50784 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_521
timestamp 1621261055
transform 1 0 51168 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_524
timestamp 1621261055
transform 1 0 51456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_532
timestamp 1621261055
transform 1 0 52224 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_540
timestamp 1621261055
transform 1 0 52992 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_548
timestamp 1621261055
transform 1 0 53760 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_556
timestamp 1621261055
transform 1 0 54528 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_564
timestamp 1621261055
transform 1 0 55296 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_772
timestamp 1621261055
transform 1 0 56640 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_572
timestamp 1621261055
transform 1 0 56064 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_576
timestamp 1621261055
transform 1 0 56448 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_579
timestamp 1621261055
transform 1 0 56736 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_587
timestamp 1621261055
transform 1 0 57504 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_113
timestamp 1621261055
transform -1 0 58848 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_595
timestamp 1621261055
transform 1 0 58272 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_114
timestamp 1621261055
transform 1 0 1152 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_57_4
timestamp 1621261055
transform 1 0 1536 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_12
timestamp 1621261055
transform 1 0 2304 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_20
timestamp 1621261055
transform 1 0 3072 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_28
timestamp 1621261055
transform 1 0 3840 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_36
timestamp 1621261055
transform 1 0 4608 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_773
timestamp 1621261055
transform 1 0 6432 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_44
timestamp 1621261055
transform 1 0 5376 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_52
timestamp 1621261055
transform 1 0 6144 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_54
timestamp 1621261055
transform 1 0 6336 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_56
timestamp 1621261055
transform 1 0 6528 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _136_
timestamp 1621261055
transform 1 0 8352 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_186
timestamp 1621261055
transform 1 0 8160 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_64
timestamp 1621261055
transform 1 0 7296 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_57_72
timestamp 1621261055
transform 1 0 8064 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_78
timestamp 1621261055
transform 1 0 8640 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_86
timestamp 1621261055
transform 1 0 9408 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_94
timestamp 1621261055
transform 1 0 10176 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_102
timestamp 1621261055
transform 1 0 10944 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _193_
timestamp 1621261055
transform -1 0 12480 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_774
timestamp 1621261055
transform 1 0 11712 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_210
timestamp 1621261055
transform -1 0 12192 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_111
timestamp 1621261055
transform 1 0 11808 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_118
timestamp 1621261055
transform 1 0 12480 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_126
timestamp 1621261055
transform 1 0 13248 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_134
timestamp 1621261055
transform 1 0 14016 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_142
timestamp 1621261055
transform 1 0 14784 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_775
timestamp 1621261055
transform 1 0 16992 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_150
timestamp 1621261055
transform 1 0 15552 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_158
timestamp 1621261055
transform 1 0 16320 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_162
timestamp 1621261055
transform 1 0 16704 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_164
timestamp 1621261055
transform 1 0 16896 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_166
timestamp 1621261055
transform 1 0 17088 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_174
timestamp 1621261055
transform 1 0 17856 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_182
timestamp 1621261055
transform 1 0 18624 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _088_
timestamp 1621261055
transform 1 0 19680 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_140
timestamp 1621261055
transform 1 0 19488 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_190
timestamp 1621261055
transform 1 0 19392 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_196
timestamp 1621261055
transform 1 0 19968 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_204
timestamp 1621261055
transform 1 0 20736 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_776
timestamp 1621261055
transform 1 0 22272 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_212
timestamp 1621261055
transform 1 0 21504 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_221
timestamp 1621261055
transform 1 0 22368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_229
timestamp 1621261055
transform 1 0 23136 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_237
timestamp 1621261055
transform 1 0 23904 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_245
timestamp 1621261055
transform 1 0 24672 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_253
timestamp 1621261055
transform 1 0 25440 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_261
timestamp 1621261055
transform 1 0 26208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_269
timestamp 1621261055
transform 1 0 26976 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_273
timestamp 1621261055
transform 1 0 27360 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_777
timestamp 1621261055
transform 1 0 27552 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_276
timestamp 1621261055
transform 1 0 27648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_284
timestamp 1621261055
transform 1 0 28416 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_292
timestamp 1621261055
transform 1 0 29184 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_300
timestamp 1621261055
transform 1 0 29952 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_308
timestamp 1621261055
transform 1 0 30720 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_778
timestamp 1621261055
transform 1 0 32832 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_316
timestamp 1621261055
transform 1 0 31488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_324
timestamp 1621261055
transform 1 0 32256 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_328
timestamp 1621261055
transform 1 0 32640 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_331
timestamp 1621261055
transform 1 0 32928 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_339
timestamp 1621261055
transform 1 0 33696 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_347
timestamp 1621261055
transform 1 0 34464 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_355
timestamp 1621261055
transform 1 0 35232 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_363
timestamp 1621261055
transform 1 0 36000 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_371
timestamp 1621261055
transform 1 0 36768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_779
timestamp 1621261055
transform 1 0 38112 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_379
timestamp 1621261055
transform 1 0 37536 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_383
timestamp 1621261055
transform 1 0 37920 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_386
timestamp 1621261055
transform 1 0 38208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_394
timestamp 1621261055
transform 1 0 38976 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _085_
timestamp 1621261055
transform -1 0 40800 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_138
timestamp 1621261055
transform -1 0 40512 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_57_402
timestamp 1621261055
transform 1 0 39744 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_406
timestamp 1621261055
transform 1 0 40128 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_413
timestamp 1621261055
transform 1 0 40800 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_780
timestamp 1621261055
transform 1 0 43392 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_421
timestamp 1621261055
transform 1 0 41568 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_429
timestamp 1621261055
transform 1 0 42336 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_437
timestamp 1621261055
transform 1 0 43104 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_439
timestamp 1621261055
transform 1 0 43296 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_441
timestamp 1621261055
transform 1 0 43488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_449
timestamp 1621261055
transform 1 0 44256 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_457
timestamp 1621261055
transform 1 0 45024 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_465
timestamp 1621261055
transform 1 0 45792 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_473
timestamp 1621261055
transform 1 0 46560 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_481
timestamp 1621261055
transform 1 0 47328 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_781
timestamp 1621261055
transform 1 0 48672 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_489
timestamp 1621261055
transform 1 0 48096 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_493
timestamp 1621261055
transform 1 0 48480 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_496
timestamp 1621261055
transform 1 0 48768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_504
timestamp 1621261055
transform 1 0 49536 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_512
timestamp 1621261055
transform 1 0 50304 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_520
timestamp 1621261055
transform 1 0 51072 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_528
timestamp 1621261055
transform 1 0 51840 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_536
timestamp 1621261055
transform 1 0 52608 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_544
timestamp 1621261055
transform 1 0 53376 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_782
timestamp 1621261055
transform 1 0 53952 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_548
timestamp 1621261055
transform 1 0 53760 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_551
timestamp 1621261055
transform 1 0 54048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_559
timestamp 1621261055
transform 1 0 54816 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_567
timestamp 1621261055
transform 1 0 55584 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_575
timestamp 1621261055
transform 1 0 56352 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_583
timestamp 1621261055
transform 1 0 57120 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_115
timestamp 1621261055
transform -1 0 58848 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_57_591
timestamp 1621261055
transform 1 0 57888 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_595
timestamp 1621261055
transform 1 0 58272 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_116
timestamp 1621261055
transform 1 0 1152 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_58_4
timestamp 1621261055
transform 1 0 1536 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_12
timestamp 1621261055
transform 1 0 2304 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_20
timestamp 1621261055
transform 1 0 3072 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _013_
timestamp 1621261055
transform 1 0 4704 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_783
timestamp 1621261055
transform 1 0 3840 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_29
timestamp 1621261055
transform 1 0 3936 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_40
timestamp 1621261055
transform 1 0 4992 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_48
timestamp 1621261055
transform 1 0 5760 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_56
timestamp 1621261055
transform 1 0 6528 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_784
timestamp 1621261055
transform 1 0 9120 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_64
timestamp 1621261055
transform 1 0 7296 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_72
timestamp 1621261055
transform 1 0 8064 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_80
timestamp 1621261055
transform 1 0 8832 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_82
timestamp 1621261055
transform 1 0 9024 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_84
timestamp 1621261055
transform 1 0 9216 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_92
timestamp 1621261055
transform 1 0 9984 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_100
timestamp 1621261055
transform 1 0 10752 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_108
timestamp 1621261055
transform 1 0 11520 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_116
timestamp 1621261055
transform 1 0 12288 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_124
timestamp 1621261055
transform 1 0 13056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_785
timestamp 1621261055
transform 1 0 14400 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_132
timestamp 1621261055
transform 1 0 13824 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_136
timestamp 1621261055
transform 1 0 14208 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_139
timestamp 1621261055
transform 1 0 14496 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_147
timestamp 1621261055
transform 1 0 15264 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_155
timestamp 1621261055
transform 1 0 16032 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_163
timestamp 1621261055
transform 1 0 16800 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_171
timestamp 1621261055
transform 1 0 17568 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_179
timestamp 1621261055
transform 1 0 18336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_187
timestamp 1621261055
transform 1 0 19104 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_786
timestamp 1621261055
transform 1 0 19680 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_191
timestamp 1621261055
transform 1 0 19488 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_194
timestamp 1621261055
transform 1 0 19776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_202
timestamp 1621261055
transform 1 0 20544 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_210
timestamp 1621261055
transform 1 0 21312 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_218
timestamp 1621261055
transform 1 0 22080 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_226
timestamp 1621261055
transform 1 0 22848 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_787
timestamp 1621261055
transform 1 0 24960 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_234
timestamp 1621261055
transform 1 0 23616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_242
timestamp 1621261055
transform 1 0 24384 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_246
timestamp 1621261055
transform 1 0 24768 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_249
timestamp 1621261055
transform 1 0 25056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _157_
timestamp 1621261055
transform 1 0 27360 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_101
timestamp 1621261055
transform 1 0 27168 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_257
timestamp 1621261055
transform 1 0 25824 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_265
timestamp 1621261055
transform 1 0 26592 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_269
timestamp 1621261055
transform 1 0 26976 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_276
timestamp 1621261055
transform 1 0 27648 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_284
timestamp 1621261055
transform 1 0 28416 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_292
timestamp 1621261055
transform 1 0 29184 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_788
timestamp 1621261055
transform 1 0 30240 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_300
timestamp 1621261055
transform 1 0 29952 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_302
timestamp 1621261055
transform 1 0 30144 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_304
timestamp 1621261055
transform 1 0 30336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_312
timestamp 1621261055
transform 1 0 31104 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_320
timestamp 1621261055
transform 1 0 31872 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_328
timestamp 1621261055
transform 1 0 32640 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_336
timestamp 1621261055
transform 1 0 33408 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_344
timestamp 1621261055
transform 1 0 34176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_352
timestamp 1621261055
transform 1 0 34944 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_356
timestamp 1621261055
transform 1 0 35328 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_789
timestamp 1621261055
transform 1 0 35520 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_359
timestamp 1621261055
transform 1 0 35616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_367
timestamp 1621261055
transform 1 0 36384 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_375
timestamp 1621261055
transform 1 0 37152 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_383
timestamp 1621261055
transform 1 0 37920 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_391
timestamp 1621261055
transform 1 0 38688 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_399
timestamp 1621261055
transform 1 0 39456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_790
timestamp 1621261055
transform 1 0 40800 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_407
timestamp 1621261055
transform 1 0 40224 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_411
timestamp 1621261055
transform 1 0 40608 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_414
timestamp 1621261055
transform 1 0 40896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_422
timestamp 1621261055
transform 1 0 41664 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_430
timestamp 1621261055
transform 1 0 42432 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_438
timestamp 1621261055
transform 1 0 43200 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_446
timestamp 1621261055
transform 1 0 43968 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_454
timestamp 1621261055
transform 1 0 44736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_462
timestamp 1621261055
transform 1 0 45504 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_791
timestamp 1621261055
transform 1 0 46080 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_466
timestamp 1621261055
transform 1 0 45888 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_469
timestamp 1621261055
transform 1 0 46176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_477
timestamp 1621261055
transform 1 0 46944 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_485
timestamp 1621261055
transform 1 0 47712 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_493
timestamp 1621261055
transform 1 0 48480 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_501
timestamp 1621261055
transform 1 0 49248 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_792
timestamp 1621261055
transform 1 0 51360 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_509
timestamp 1621261055
transform 1 0 50016 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_517
timestamp 1621261055
transform 1 0 50784 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_521
timestamp 1621261055
transform 1 0 51168 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_524
timestamp 1621261055
transform 1 0 51456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_532
timestamp 1621261055
transform 1 0 52224 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_540
timestamp 1621261055
transform 1 0 52992 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_548
timestamp 1621261055
transform 1 0 53760 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_556
timestamp 1621261055
transform 1 0 54528 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_564
timestamp 1621261055
transform 1 0 55296 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_793
timestamp 1621261055
transform 1 0 56640 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_572
timestamp 1621261055
transform 1 0 56064 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_576
timestamp 1621261055
transform 1 0 56448 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_579
timestamp 1621261055
transform 1 0 56736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_587
timestamp 1621261055
transform 1 0 57504 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_117
timestamp 1621261055
transform -1 0 58848 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_595
timestamp 1621261055
transform 1 0 58272 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_118
timestamp 1621261055
transform 1 0 1152 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_4
timestamp 1621261055
transform 1 0 1536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_12
timestamp 1621261055
transform 1 0 2304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_20
timestamp 1621261055
transform 1 0 3072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_28
timestamp 1621261055
transform 1 0 3840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_36
timestamp 1621261055
transform 1 0 4608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_794
timestamp 1621261055
transform 1 0 6432 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_44
timestamp 1621261055
transform 1 0 5376 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_52
timestamp 1621261055
transform 1 0 6144 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_54
timestamp 1621261055
transform 1 0 6336 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_56
timestamp 1621261055
transform 1 0 6528 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _175_
timestamp 1621261055
transform 1 0 7776 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_122
timestamp 1621261055
transform 1 0 7584 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_64
timestamp 1621261055
transform 1 0 7296 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_66
timestamp 1621261055
transform 1 0 7488 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_72
timestamp 1621261055
transform 1 0 8064 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_80
timestamp 1621261055
transform 1 0 8832 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_88
timestamp 1621261055
transform 1 0 9600 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_96
timestamp 1621261055
transform 1 0 10368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_104
timestamp 1621261055
transform 1 0 11136 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_795
timestamp 1621261055
transform 1 0 11712 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_108
timestamp 1621261055
transform 1 0 11520 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_111
timestamp 1621261055
transform 1 0 11808 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_119
timestamp 1621261055
transform 1 0 12576 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_127
timestamp 1621261055
transform 1 0 13344 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_135
timestamp 1621261055
transform 1 0 14112 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_143
timestamp 1621261055
transform 1 0 14880 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_796
timestamp 1621261055
transform 1 0 16992 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_151
timestamp 1621261055
transform 1 0 15648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_159
timestamp 1621261055
transform 1 0 16416 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_163
timestamp 1621261055
transform 1 0 16800 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_166
timestamp 1621261055
transform 1 0 17088 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_174
timestamp 1621261055
transform 1 0 17856 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_182
timestamp 1621261055
transform 1 0 18624 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_190
timestamp 1621261055
transform 1 0 19392 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_198
timestamp 1621261055
transform 1 0 20160 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_206
timestamp 1621261055
transform 1 0 20928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_797
timestamp 1621261055
transform 1 0 22272 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_214
timestamp 1621261055
transform 1 0 21696 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_218
timestamp 1621261055
transform 1 0 22080 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_221
timestamp 1621261055
transform 1 0 22368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_229
timestamp 1621261055
transform 1 0 23136 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_237
timestamp 1621261055
transform 1 0 23904 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_245
timestamp 1621261055
transform 1 0 24672 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_253
timestamp 1621261055
transform 1 0 25440 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_261
timestamp 1621261055
transform 1 0 26208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_269
timestamp 1621261055
transform 1 0 26976 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_273
timestamp 1621261055
transform 1 0 27360 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_798
timestamp 1621261055
transform 1 0 27552 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_276
timestamp 1621261055
transform 1 0 27648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_284
timestamp 1621261055
transform 1 0 28416 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_292
timestamp 1621261055
transform 1 0 29184 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_300
timestamp 1621261055
transform 1 0 29952 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_308
timestamp 1621261055
transform 1 0 30720 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_799
timestamp 1621261055
transform 1 0 32832 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_316
timestamp 1621261055
transform 1 0 31488 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_324
timestamp 1621261055
transform 1 0 32256 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_328
timestamp 1621261055
transform 1 0 32640 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_331
timestamp 1621261055
transform 1 0 32928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_339
timestamp 1621261055
transform 1 0 33696 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_347
timestamp 1621261055
transform 1 0 34464 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_355
timestamp 1621261055
transform 1 0 35232 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_363
timestamp 1621261055
transform 1 0 36000 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_371
timestamp 1621261055
transform 1 0 36768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_800
timestamp 1621261055
transform 1 0 38112 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_379
timestamp 1621261055
transform 1 0 37536 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_383
timestamp 1621261055
transform 1 0 37920 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_386
timestamp 1621261055
transform 1 0 38208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_394
timestamp 1621261055
transform 1 0 38976 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_402
timestamp 1621261055
transform 1 0 39744 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_410
timestamp 1621261055
transform 1 0 40512 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_418
timestamp 1621261055
transform 1 0 41280 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_801
timestamp 1621261055
transform 1 0 43392 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_426
timestamp 1621261055
transform 1 0 42048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_434
timestamp 1621261055
transform 1 0 42816 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_438
timestamp 1621261055
transform 1 0 43200 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_441
timestamp 1621261055
transform 1 0 43488 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_449
timestamp 1621261055
transform 1 0 44256 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_457
timestamp 1621261055
transform 1 0 45024 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_465
timestamp 1621261055
transform 1 0 45792 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_473
timestamp 1621261055
transform 1 0 46560 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_481
timestamp 1621261055
transform 1 0 47328 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_802
timestamp 1621261055
transform 1 0 48672 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_489
timestamp 1621261055
transform 1 0 48096 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_493
timestamp 1621261055
transform 1 0 48480 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_496
timestamp 1621261055
transform 1 0 48768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_504
timestamp 1621261055
transform 1 0 49536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_512
timestamp 1621261055
transform 1 0 50304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_520
timestamp 1621261055
transform 1 0 51072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_528
timestamp 1621261055
transform 1 0 51840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_536
timestamp 1621261055
transform 1 0 52608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_544
timestamp 1621261055
transform 1 0 53376 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_803
timestamp 1621261055
transform 1 0 53952 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_548
timestamp 1621261055
transform 1 0 53760 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_551
timestamp 1621261055
transform 1 0 54048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_559
timestamp 1621261055
transform 1 0 54816 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_567
timestamp 1621261055
transform 1 0 55584 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_575
timestamp 1621261055
transform 1 0 56352 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_583
timestamp 1621261055
transform 1 0 57120 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_119
timestamp 1621261055
transform -1 0 58848 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_59_591
timestamp 1621261055
transform 1 0 57888 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_595
timestamp 1621261055
transform 1 0 58272 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_120
timestamp 1621261055
transform 1 0 1152 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_60_4
timestamp 1621261055
transform 1 0 1536 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_12
timestamp 1621261055
transform 1 0 2304 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_20
timestamp 1621261055
transform 1 0 3072 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_804
timestamp 1621261055
transform 1 0 3840 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_29
timestamp 1621261055
transform 1 0 3936 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_37
timestamp 1621261055
transform 1 0 4704 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _051_
timestamp 1621261055
transform 1 0 6336 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_60_45
timestamp 1621261055
transform 1 0 5472 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_60_53
timestamp 1621261055
transform 1 0 6240 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_57
timestamp 1621261055
transform 1 0 6624 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_805
timestamp 1621261055
transform 1 0 9120 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_65
timestamp 1621261055
transform 1 0 7392 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_73
timestamp 1621261055
transform 1 0 8160 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_81
timestamp 1621261055
transform 1 0 8928 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_84
timestamp 1621261055
transform 1 0 9216 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_92
timestamp 1621261055
transform 1 0 9984 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_100
timestamp 1621261055
transform 1 0 10752 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_108
timestamp 1621261055
transform 1 0 11520 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_116
timestamp 1621261055
transform 1 0 12288 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_124
timestamp 1621261055
transform 1 0 13056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_806
timestamp 1621261055
transform 1 0 14400 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_132
timestamp 1621261055
transform 1 0 13824 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_136
timestamp 1621261055
transform 1 0 14208 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_139
timestamp 1621261055
transform 1 0 14496 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_147
timestamp 1621261055
transform 1 0 15264 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_155
timestamp 1621261055
transform 1 0 16032 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_163
timestamp 1621261055
transform 1 0 16800 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_171
timestamp 1621261055
transform 1 0 17568 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_179
timestamp 1621261055
transform 1 0 18336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_187
timestamp 1621261055
transform 1 0 19104 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_807
timestamp 1621261055
transform 1 0 19680 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_191
timestamp 1621261055
transform 1 0 19488 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_194
timestamp 1621261055
transform 1 0 19776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_202
timestamp 1621261055
transform 1 0 20544 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_210
timestamp 1621261055
transform 1 0 21312 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_218
timestamp 1621261055
transform 1 0 22080 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_226
timestamp 1621261055
transform 1 0 22848 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_808
timestamp 1621261055
transform 1 0 24960 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_234
timestamp 1621261055
transform 1 0 23616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_242
timestamp 1621261055
transform 1 0 24384 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_246
timestamp 1621261055
transform 1 0 24768 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_249
timestamp 1621261055
transform 1 0 25056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_257
timestamp 1621261055
transform 1 0 25824 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_265
timestamp 1621261055
transform 1 0 26592 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_273
timestamp 1621261055
transform 1 0 27360 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_281
timestamp 1621261055
transform 1 0 28128 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_289
timestamp 1621261055
transform 1 0 28896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_809
timestamp 1621261055
transform 1 0 30240 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_297
timestamp 1621261055
transform 1 0 29664 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_301
timestamp 1621261055
transform 1 0 30048 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_304
timestamp 1621261055
transform 1 0 30336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_312
timestamp 1621261055
transform 1 0 31104 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_320
timestamp 1621261055
transform 1 0 31872 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_328
timestamp 1621261055
transform 1 0 32640 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_336
timestamp 1621261055
transform 1 0 33408 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_344
timestamp 1621261055
transform 1 0 34176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_352
timestamp 1621261055
transform 1 0 34944 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_356
timestamp 1621261055
transform 1 0 35328 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_810
timestamp 1621261055
transform 1 0 35520 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_359
timestamp 1621261055
transform 1 0 35616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_367
timestamp 1621261055
transform 1 0 36384 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_375
timestamp 1621261055
transform 1 0 37152 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_383
timestamp 1621261055
transform 1 0 37920 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_391
timestamp 1621261055
transform 1 0 38688 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_399
timestamp 1621261055
transform 1 0 39456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_811
timestamp 1621261055
transform 1 0 40800 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_407
timestamp 1621261055
transform 1 0 40224 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_411
timestamp 1621261055
transform 1 0 40608 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_414
timestamp 1621261055
transform 1 0 40896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_422
timestamp 1621261055
transform 1 0 41664 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_430
timestamp 1621261055
transform 1 0 42432 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_438
timestamp 1621261055
transform 1 0 43200 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_446
timestamp 1621261055
transform 1 0 43968 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_454
timestamp 1621261055
transform 1 0 44736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_462
timestamp 1621261055
transform 1 0 45504 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _149_
timestamp 1621261055
transform 1 0 46560 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_812
timestamp 1621261055
transform 1 0 46080 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_201
timestamp 1621261055
transform 1 0 46368 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_466
timestamp 1621261055
transform 1 0 45888 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_469
timestamp 1621261055
transform 1 0 46176 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_476
timestamp 1621261055
transform 1 0 46848 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_484
timestamp 1621261055
transform 1 0 47616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_492
timestamp 1621261055
transform 1 0 48384 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_500
timestamp 1621261055
transform 1 0 49152 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_813
timestamp 1621261055
transform 1 0 51360 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_508
timestamp 1621261055
transform 1 0 49920 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_516
timestamp 1621261055
transform 1 0 50688 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_520
timestamp 1621261055
transform 1 0 51072 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_522
timestamp 1621261055
transform 1 0 51264 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_524
timestamp 1621261055
transform 1 0 51456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_532
timestamp 1621261055
transform 1 0 52224 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_540
timestamp 1621261055
transform 1 0 52992 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _104_
timestamp 1621261055
transform -1 0 54432 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_163
timestamp 1621261055
transform -1 0 54144 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_548
timestamp 1621261055
transform 1 0 53760 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_555
timestamp 1621261055
transform 1 0 54432 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_563
timestamp 1621261055
transform 1 0 55200 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_814
timestamp 1621261055
transform 1 0 56640 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_571
timestamp 1621261055
transform 1 0 55968 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_575
timestamp 1621261055
transform 1 0 56352 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_577
timestamp 1621261055
transform 1 0 56544 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_579
timestamp 1621261055
transform 1 0 56736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_587
timestamp 1621261055
transform 1 0 57504 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_121
timestamp 1621261055
transform -1 0 58848 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_595
timestamp 1621261055
transform 1 0 58272 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_122
timestamp 1621261055
transform 1 0 1152 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_124
timestamp 1621261055
transform 1 0 1152 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_4
timestamp 1621261055
transform 1 0 1536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_12
timestamp 1621261055
transform 1 0 2304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_20
timestamp 1621261055
transform 1 0 3072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_4
timestamp 1621261055
transform 1 0 1536 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_12
timestamp 1621261055
transform 1 0 2304 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_20
timestamp 1621261055
transform 1 0 3072 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_825
timestamp 1621261055
transform 1 0 3840 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_28
timestamp 1621261055
transform 1 0 3840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_36
timestamp 1621261055
transform 1 0 4608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_29
timestamp 1621261055
transform 1 0 3936 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_37
timestamp 1621261055
transform 1 0 4704 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_815
timestamp 1621261055
transform 1 0 6432 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_44
timestamp 1621261055
transform 1 0 5376 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_52
timestamp 1621261055
transform 1 0 6144 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_61_54
timestamp 1621261055
transform 1 0 6336 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_56
timestamp 1621261055
transform 1 0 6528 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_45
timestamp 1621261055
transform 1 0 5472 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_53
timestamp 1621261055
transform 1 0 6240 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_61
timestamp 1621261055
transform 1 0 7008 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_826
timestamp 1621261055
transform 1 0 9120 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_64
timestamp 1621261055
transform 1 0 7296 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_72
timestamp 1621261055
transform 1 0 8064 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_80
timestamp 1621261055
transform 1 0 8832 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_69
timestamp 1621261055
transform 1 0 7776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_77
timestamp 1621261055
transform 1 0 8544 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_81
timestamp 1621261055
transform 1 0 8928 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_84
timestamp 1621261055
transform 1 0 9216 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _140_
timestamp 1621261055
transform 1 0 11136 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_190
timestamp 1621261055
transform 1 0 10944 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_88
timestamp 1621261055
transform 1 0 9600 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_96
timestamp 1621261055
transform 1 0 10368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_104
timestamp 1621261055
transform 1 0 11136 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_92
timestamp 1621261055
transform 1 0 9984 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_100
timestamp 1621261055
transform 1 0 10752 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_107
timestamp 1621261055
transform 1 0 11424 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_111
timestamp 1621261055
transform 1 0 11808 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_108
timestamp 1621261055
transform 1 0 11520 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_816
timestamp 1621261055
transform 1 0 11712 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_115
timestamp 1621261055
transform 1 0 12192 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_121
timestamp 1621261055
transform 1 0 12768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_115
timestamp 1621261055
transform 1 0 12192 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_184
timestamp 1621261055
transform 1 0 12288 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _065_
timestamp 1621261055
transform 1 0 12480 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_123
timestamp 1621261055
transform 1 0 12960 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_827
timestamp 1621261055
transform 1 0 14400 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_129
timestamp 1621261055
transform 1 0 13536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_137
timestamp 1621261055
transform 1 0 14304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_145
timestamp 1621261055
transform 1 0 15072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_131
timestamp 1621261055
transform 1 0 13728 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_135
timestamp 1621261055
transform 1 0 14112 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_62_137
timestamp 1621261055
transform 1 0 14304 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_139
timestamp 1621261055
transform 1 0 14496 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_147
timestamp 1621261055
transform 1 0 15264 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_817
timestamp 1621261055
transform 1 0 16992 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_153
timestamp 1621261055
transform 1 0 15840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_161
timestamp 1621261055
transform 1 0 16608 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_166
timestamp 1621261055
transform 1 0 17088 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_155
timestamp 1621261055
transform 1 0 16032 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_163
timestamp 1621261055
transform 1 0 16800 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_174
timestamp 1621261055
transform 1 0 17856 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_182
timestamp 1621261055
transform 1 0 18624 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_171
timestamp 1621261055
transform 1 0 17568 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_179
timestamp 1621261055
transform 1 0 18336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_187
timestamp 1621261055
transform 1 0 19104 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_828
timestamp 1621261055
transform 1 0 19680 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_190
timestamp 1621261055
transform 1 0 19392 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_198
timestamp 1621261055
transform 1 0 20160 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_206
timestamp 1621261055
transform 1 0 20928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_191
timestamp 1621261055
transform 1 0 19488 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_194
timestamp 1621261055
transform 1 0 19776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_202
timestamp 1621261055
transform 1 0 20544 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_210
timestamp 1621261055
transform 1 0 21312 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_818
timestamp 1621261055
transform 1 0 22272 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_214
timestamp 1621261055
transform 1 0 21696 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_218
timestamp 1621261055
transform 1 0 22080 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_221
timestamp 1621261055
transform 1 0 22368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_229
timestamp 1621261055
transform 1 0 23136 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_218
timestamp 1621261055
transform 1 0 22080 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_226
timestamp 1621261055
transform 1 0 22848 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_829
timestamp 1621261055
transform 1 0 24960 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_237
timestamp 1621261055
transform 1 0 23904 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_245
timestamp 1621261055
transform 1 0 24672 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_234
timestamp 1621261055
transform 1 0 23616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_242
timestamp 1621261055
transform 1 0 24384 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_246
timestamp 1621261055
transform 1 0 24768 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_249
timestamp 1621261055
transform 1 0 25056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_253
timestamp 1621261055
transform 1 0 25440 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_261
timestamp 1621261055
transform 1 0 26208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_269
timestamp 1621261055
transform 1 0 26976 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_273
timestamp 1621261055
transform 1 0 27360 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_257
timestamp 1621261055
transform 1 0 25824 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_265
timestamp 1621261055
transform 1 0 26592 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_273
timestamp 1621261055
transform 1 0 27360 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_819
timestamp 1621261055
transform 1 0 27552 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_276
timestamp 1621261055
transform 1 0 27648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_284
timestamp 1621261055
transform 1 0 28416 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_292
timestamp 1621261055
transform 1 0 29184 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_281
timestamp 1621261055
transform 1 0 28128 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_289
timestamp 1621261055
transform 1 0 28896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_830
timestamp 1621261055
transform 1 0 30240 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_300
timestamp 1621261055
transform 1 0 29952 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_308
timestamp 1621261055
transform 1 0 30720 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_297
timestamp 1621261055
transform 1 0 29664 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_301
timestamp 1621261055
transform 1 0 30048 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_304
timestamp 1621261055
transform 1 0 30336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_312
timestamp 1621261055
transform 1 0 31104 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_820
timestamp 1621261055
transform 1 0 32832 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_316
timestamp 1621261055
transform 1 0 31488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_324
timestamp 1621261055
transform 1 0 32256 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_328
timestamp 1621261055
transform 1 0 32640 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_331
timestamp 1621261055
transform 1 0 32928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_320
timestamp 1621261055
transform 1 0 31872 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_328
timestamp 1621261055
transform 1 0 32640 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_336
timestamp 1621261055
transform 1 0 33408 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_339
timestamp 1621261055
transform 1 0 33696 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_347
timestamp 1621261055
transform 1 0 34464 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_355
timestamp 1621261055
transform 1 0 35232 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_344
timestamp 1621261055
transform 1 0 34176 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_352
timestamp 1621261055
transform 1 0 34944 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_356
timestamp 1621261055
transform 1 0 35328 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_831
timestamp 1621261055
transform 1 0 35520 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_363
timestamp 1621261055
transform 1 0 36000 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_371
timestamp 1621261055
transform 1 0 36768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_359
timestamp 1621261055
transform 1 0 35616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_367
timestamp 1621261055
transform 1 0 36384 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_375
timestamp 1621261055
transform 1 0 37152 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_821
timestamp 1621261055
transform 1 0 38112 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_379
timestamp 1621261055
transform 1 0 37536 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_383
timestamp 1621261055
transform 1 0 37920 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_386
timestamp 1621261055
transform 1 0 38208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_394
timestamp 1621261055
transform 1 0 38976 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_383
timestamp 1621261055
transform 1 0 37920 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_391
timestamp 1621261055
transform 1 0 38688 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_399
timestamp 1621261055
transform 1 0 39456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_832
timestamp 1621261055
transform 1 0 40800 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_402
timestamp 1621261055
transform 1 0 39744 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_410
timestamp 1621261055
transform 1 0 40512 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_418
timestamp 1621261055
transform 1 0 41280 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_407
timestamp 1621261055
transform 1 0 40224 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_411
timestamp 1621261055
transform 1 0 40608 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_414
timestamp 1621261055
transform 1 0 40896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_822
timestamp 1621261055
transform 1 0 43392 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_426
timestamp 1621261055
transform 1 0 42048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_434
timestamp 1621261055
transform 1 0 42816 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_438
timestamp 1621261055
transform 1 0 43200 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_441
timestamp 1621261055
transform 1 0 43488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_422
timestamp 1621261055
transform 1 0 41664 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_430
timestamp 1621261055
transform 1 0 42432 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_438
timestamp 1621261055
transform 1 0 43200 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_449
timestamp 1621261055
transform 1 0 44256 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_457
timestamp 1621261055
transform 1 0 45024 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_446
timestamp 1621261055
transform 1 0 43968 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_454
timestamp 1621261055
transform 1 0 44736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_462
timestamp 1621261055
transform 1 0 45504 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_833
timestamp 1621261055
transform 1 0 46080 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_465
timestamp 1621261055
transform 1 0 45792 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_473
timestamp 1621261055
transform 1 0 46560 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_481
timestamp 1621261055
transform 1 0 47328 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_466
timestamp 1621261055
transform 1 0 45888 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_469
timestamp 1621261055
transform 1 0 46176 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_477
timestamp 1621261055
transform 1 0 46944 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_823
timestamp 1621261055
transform 1 0 48672 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_489
timestamp 1621261055
transform 1 0 48096 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_493
timestamp 1621261055
transform 1 0 48480 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_496
timestamp 1621261055
transform 1 0 48768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_504
timestamp 1621261055
transform 1 0 49536 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_485
timestamp 1621261055
transform 1 0 47712 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_493
timestamp 1621261055
transform 1 0 48480 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_501
timestamp 1621261055
transform 1 0 49248 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_509
timestamp 1621261055
transform 1 0 50016 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_512
timestamp 1621261055
transform 1 0 50304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_506
timestamp 1621261055
transform 1 0 49728 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_208
timestamp 1621261055
transform -1 0 50016 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _183_
timestamp 1621261055
transform -1 0 50304 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_521
timestamp 1621261055
transform 1 0 51168 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_517
timestamp 1621261055
transform 1 0 50784 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_520
timestamp 1621261055
transform 1 0 51072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_524
timestamp 1621261055
transform 1 0 51456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_834
timestamp 1621261055
transform 1 0 51360 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_528
timestamp 1621261055
transform 1 0 51840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_536
timestamp 1621261055
transform 1 0 52608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_544
timestamp 1621261055
transform 1 0 53376 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_532
timestamp 1621261055
transform 1 0 52224 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_540
timestamp 1621261055
transform 1 0 52992 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_824
timestamp 1621261055
transform 1 0 53952 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_548
timestamp 1621261055
transform 1 0 53760 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_551
timestamp 1621261055
transform 1 0 54048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_559
timestamp 1621261055
transform 1 0 54816 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_567
timestamp 1621261055
transform 1 0 55584 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_548
timestamp 1621261055
transform 1 0 53760 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_556
timestamp 1621261055
transform 1 0 54528 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_564
timestamp 1621261055
transform 1 0 55296 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_835
timestamp 1621261055
transform 1 0 56640 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_575
timestamp 1621261055
transform 1 0 56352 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_583
timestamp 1621261055
transform 1 0 57120 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_572
timestamp 1621261055
transform 1 0 56064 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_576
timestamp 1621261055
transform 1 0 56448 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_579
timestamp 1621261055
transform 1 0 56736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_587
timestamp 1621261055
transform 1 0 57504 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_123
timestamp 1621261055
transform -1 0 58848 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_125
timestamp 1621261055
transform -1 0 58848 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_61_591
timestamp 1621261055
transform 1 0 57888 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_595
timestamp 1621261055
transform 1 0 58272 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_595
timestamp 1621261055
transform 1 0 58272 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_126
timestamp 1621261055
transform 1 0 1152 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_4
timestamp 1621261055
transform 1 0 1536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_12
timestamp 1621261055
transform 1 0 2304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_20
timestamp 1621261055
transform 1 0 3072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_28
timestamp 1621261055
transform 1 0 3840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_36
timestamp 1621261055
transform 1 0 4608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_836
timestamp 1621261055
transform 1 0 6432 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_44
timestamp 1621261055
transform 1 0 5376 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_52
timestamp 1621261055
transform 1 0 6144 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_54
timestamp 1621261055
transform 1 0 6336 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_56
timestamp 1621261055
transform 1 0 6528 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _008_
timestamp 1621261055
transform 1 0 7584 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _205_
timestamp 1621261055
transform 1 0 8256 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_226
timestamp 1621261055
transform 1 0 8064 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_64
timestamp 1621261055
transform 1 0 7296 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_66
timestamp 1621261055
transform 1 0 7488 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_70
timestamp 1621261055
transform 1 0 7872 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_77
timestamp 1621261055
transform 1 0 8544 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_85
timestamp 1621261055
transform 1 0 9312 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_93
timestamp 1621261055
transform 1 0 10080 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_101
timestamp 1621261055
transform 1 0 10848 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_837
timestamp 1621261055
transform 1 0 11712 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_63_109
timestamp 1621261055
transform 1 0 11616 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_111
timestamp 1621261055
transform 1 0 11808 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_119
timestamp 1621261055
transform 1 0 12576 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_127
timestamp 1621261055
transform 1 0 13344 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_135
timestamp 1621261055
transform 1 0 14112 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_143
timestamp 1621261055
transform 1 0 14880 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_838
timestamp 1621261055
transform 1 0 16992 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_151
timestamp 1621261055
transform 1 0 15648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_159
timestamp 1621261055
transform 1 0 16416 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_163
timestamp 1621261055
transform 1 0 16800 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_166
timestamp 1621261055
transform 1 0 17088 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_174
timestamp 1621261055
transform 1 0 17856 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_182
timestamp 1621261055
transform 1 0 18624 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _142_
timestamp 1621261055
transform 1 0 21120 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_194
timestamp 1621261055
transform 1 0 20928 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_190
timestamp 1621261055
transform 1 0 19392 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_198
timestamp 1621261055
transform 1 0 20160 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_839
timestamp 1621261055
transform 1 0 22272 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_211
timestamp 1621261055
transform 1 0 21408 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_63_219
timestamp 1621261055
transform 1 0 22176 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_221
timestamp 1621261055
transform 1 0 22368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_229
timestamp 1621261055
transform 1 0 23136 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_237
timestamp 1621261055
transform 1 0 23904 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_245
timestamp 1621261055
transform 1 0 24672 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_253
timestamp 1621261055
transform 1 0 25440 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_261
timestamp 1621261055
transform 1 0 26208 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_269
timestamp 1621261055
transform 1 0 26976 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_273
timestamp 1621261055
transform 1 0 27360 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_840
timestamp 1621261055
transform 1 0 27552 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_276
timestamp 1621261055
transform 1 0 27648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_284
timestamp 1621261055
transform 1 0 28416 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_292
timestamp 1621261055
transform 1 0 29184 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_300
timestamp 1621261055
transform 1 0 29952 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_308
timestamp 1621261055
transform 1 0 30720 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_841
timestamp 1621261055
transform 1 0 32832 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_316
timestamp 1621261055
transform 1 0 31488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_324
timestamp 1621261055
transform 1 0 32256 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_328
timestamp 1621261055
transform 1 0 32640 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_331
timestamp 1621261055
transform 1 0 32928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_339
timestamp 1621261055
transform 1 0 33696 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_347
timestamp 1621261055
transform 1 0 34464 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_355
timestamp 1621261055
transform 1 0 35232 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_363
timestamp 1621261055
transform 1 0 36000 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_371
timestamp 1621261055
transform 1 0 36768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _056_
timestamp 1621261055
transform 1 0 38592 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_842
timestamp 1621261055
transform 1 0 38112 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_379
timestamp 1621261055
transform 1 0 37536 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_383
timestamp 1621261055
transform 1 0 37920 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_63_386
timestamp 1621261055
transform 1 0 38208 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_393
timestamp 1621261055
transform 1 0 38880 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _070_
timestamp 1621261055
transform -1 0 41472 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_128
timestamp 1621261055
transform -1 0 41184 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_401
timestamp 1621261055
transform 1 0 39648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_409
timestamp 1621261055
transform 1 0 40416 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_413
timestamp 1621261055
transform 1 0 40800 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_420
timestamp 1621261055
transform 1 0 41472 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_843
timestamp 1621261055
transform 1 0 43392 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_428
timestamp 1621261055
transform 1 0 42240 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_436
timestamp 1621261055
transform 1 0 43008 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_441
timestamp 1621261055
transform 1 0 43488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_449
timestamp 1621261055
transform 1 0 44256 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_457
timestamp 1621261055
transform 1 0 45024 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_465
timestamp 1621261055
transform 1 0 45792 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_473
timestamp 1621261055
transform 1 0 46560 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_481
timestamp 1621261055
transform 1 0 47328 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_844
timestamp 1621261055
transform 1 0 48672 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_489
timestamp 1621261055
transform 1 0 48096 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_493
timestamp 1621261055
transform 1 0 48480 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_496
timestamp 1621261055
transform 1 0 48768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_504
timestamp 1621261055
transform 1 0 49536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_512
timestamp 1621261055
transform 1 0 50304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_520
timestamp 1621261055
transform 1 0 51072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _039_
timestamp 1621261055
transform 1 0 53280 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_63_528
timestamp 1621261055
transform 1 0 51840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_536
timestamp 1621261055
transform 1 0 52608 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_540
timestamp 1621261055
transform 1 0 52992 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_542
timestamp 1621261055
transform 1 0 53184 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_546
timestamp 1621261055
transform 1 0 53568 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_845
timestamp 1621261055
transform 1 0 53952 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_551
timestamp 1621261055
transform 1 0 54048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_559
timestamp 1621261055
transform 1 0 54816 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_567
timestamp 1621261055
transform 1 0 55584 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_575
timestamp 1621261055
transform 1 0 56352 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_583
timestamp 1621261055
transform 1 0 57120 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_127
timestamp 1621261055
transform -1 0 58848 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_63_591
timestamp 1621261055
transform 1 0 57888 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_595
timestamp 1621261055
transform 1 0 58272 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_128
timestamp 1621261055
transform 1 0 1152 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_64_4
timestamp 1621261055
transform 1 0 1536 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_12
timestamp 1621261055
transform 1 0 2304 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_20
timestamp 1621261055
transform 1 0 3072 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_846
timestamp 1621261055
transform 1 0 3840 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_29
timestamp 1621261055
transform 1 0 3936 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_37
timestamp 1621261055
transform 1 0 4704 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_45
timestamp 1621261055
transform 1 0 5472 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_53
timestamp 1621261055
transform 1 0 6240 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_61
timestamp 1621261055
transform 1 0 7008 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_847
timestamp 1621261055
transform 1 0 9120 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_69
timestamp 1621261055
transform 1 0 7776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_77
timestamp 1621261055
transform 1 0 8544 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_81
timestamp 1621261055
transform 1 0 8928 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_84
timestamp 1621261055
transform 1 0 9216 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_92
timestamp 1621261055
transform 1 0 9984 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_100
timestamp 1621261055
transform 1 0 10752 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_108
timestamp 1621261055
transform 1 0 11520 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_116
timestamp 1621261055
transform 1 0 12288 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_124
timestamp 1621261055
transform 1 0 13056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_848
timestamp 1621261055
transform 1 0 14400 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_132
timestamp 1621261055
transform 1 0 13824 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_136
timestamp 1621261055
transform 1 0 14208 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_139
timestamp 1621261055
transform 1 0 14496 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_147
timestamp 1621261055
transform 1 0 15264 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_155
timestamp 1621261055
transform 1 0 16032 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_163
timestamp 1621261055
transform 1 0 16800 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_171
timestamp 1621261055
transform 1 0 17568 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_179
timestamp 1621261055
transform 1 0 18336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_187
timestamp 1621261055
transform 1 0 19104 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_849
timestamp 1621261055
transform 1 0 19680 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_191
timestamp 1621261055
transform 1 0 19488 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_194
timestamp 1621261055
transform 1 0 19776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_202
timestamp 1621261055
transform 1 0 20544 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_210
timestamp 1621261055
transform 1 0 21312 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_218
timestamp 1621261055
transform 1 0 22080 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_226
timestamp 1621261055
transform 1 0 22848 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_850
timestamp 1621261055
transform 1 0 24960 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_234
timestamp 1621261055
transform 1 0 23616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_242
timestamp 1621261055
transform 1 0 24384 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_246
timestamp 1621261055
transform 1 0 24768 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_249
timestamp 1621261055
transform 1 0 25056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_257
timestamp 1621261055
transform 1 0 25824 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_265
timestamp 1621261055
transform 1 0 26592 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_273
timestamp 1621261055
transform 1 0 27360 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_281
timestamp 1621261055
transform 1 0 28128 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_289
timestamp 1621261055
transform 1 0 28896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_851
timestamp 1621261055
transform 1 0 30240 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_297
timestamp 1621261055
transform 1 0 29664 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_301
timestamp 1621261055
transform 1 0 30048 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_304
timestamp 1621261055
transform 1 0 30336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_312
timestamp 1621261055
transform 1 0 31104 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_320
timestamp 1621261055
transform 1 0 31872 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_328
timestamp 1621261055
transform 1 0 32640 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_336
timestamp 1621261055
transform 1 0 33408 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _054_
timestamp 1621261055
transform 1 0 34848 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_64_344
timestamp 1621261055
transform 1 0 34176 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_348
timestamp 1621261055
transform 1 0 34560 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_64_350
timestamp 1621261055
transform 1 0 34752 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_354
timestamp 1621261055
transform 1 0 35136 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_852
timestamp 1621261055
transform 1 0 35520 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_359
timestamp 1621261055
transform 1 0 35616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_367
timestamp 1621261055
transform 1 0 36384 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_375
timestamp 1621261055
transform 1 0 37152 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_383
timestamp 1621261055
transform 1 0 37920 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_391
timestamp 1621261055
transform 1 0 38688 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_399
timestamp 1621261055
transform 1 0 39456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_853
timestamp 1621261055
transform 1 0 40800 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_407
timestamp 1621261055
transform 1 0 40224 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_411
timestamp 1621261055
transform 1 0 40608 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_414
timestamp 1621261055
transform 1 0 40896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_422
timestamp 1621261055
transform 1 0 41664 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_430
timestamp 1621261055
transform 1 0 42432 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_438
timestamp 1621261055
transform 1 0 43200 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_446
timestamp 1621261055
transform 1 0 43968 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_454
timestamp 1621261055
transform 1 0 44736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_462
timestamp 1621261055
transform 1 0 45504 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_854
timestamp 1621261055
transform 1 0 46080 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_466
timestamp 1621261055
transform 1 0 45888 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_469
timestamp 1621261055
transform 1 0 46176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_477
timestamp 1621261055
transform 1 0 46944 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_485
timestamp 1621261055
transform 1 0 47712 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_493
timestamp 1621261055
transform 1 0 48480 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_501
timestamp 1621261055
transform 1 0 49248 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_855
timestamp 1621261055
transform 1 0 51360 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_509
timestamp 1621261055
transform 1 0 50016 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_517
timestamp 1621261055
transform 1 0 50784 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_521
timestamp 1621261055
transform 1 0 51168 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_524
timestamp 1621261055
transform 1 0 51456 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _072_
timestamp 1621261055
transform -1 0 52128 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_132
timestamp 1621261055
transform -1 0 51840 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_531
timestamp 1621261055
transform 1 0 52128 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_539
timestamp 1621261055
transform 1 0 52896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_547
timestamp 1621261055
transform 1 0 53664 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_555
timestamp 1621261055
transform 1 0 54432 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_563
timestamp 1621261055
transform 1 0 55200 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_856
timestamp 1621261055
transform 1 0 56640 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_571
timestamp 1621261055
transform 1 0 55968 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_575
timestamp 1621261055
transform 1 0 56352 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_64_577
timestamp 1621261055
transform 1 0 56544 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_579
timestamp 1621261055
transform 1 0 56736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_587
timestamp 1621261055
transform 1 0 57504 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_129
timestamp 1621261055
transform -1 0 58848 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_595
timestamp 1621261055
transform 1 0 58272 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_130
timestamp 1621261055
transform 1 0 1152 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_4
timestamp 1621261055
transform 1 0 1536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_12
timestamp 1621261055
transform 1 0 2304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_20
timestamp 1621261055
transform 1 0 3072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_28
timestamp 1621261055
transform 1 0 3840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_36
timestamp 1621261055
transform 1 0 4608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_857
timestamp 1621261055
transform 1 0 6432 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_44
timestamp 1621261055
transform 1 0 5376 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_52
timestamp 1621261055
transform 1 0 6144 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_54
timestamp 1621261055
transform 1 0 6336 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_56
timestamp 1621261055
transform 1 0 6528 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_64
timestamp 1621261055
transform 1 0 7296 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_72
timestamp 1621261055
transform 1 0 8064 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_80
timestamp 1621261055
transform 1 0 8832 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_84
timestamp 1621261055
transform 1 0 9216 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _209_
timestamp 1621261055
transform 1 0 9696 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_228
timestamp 1621261055
transform 1 0 9504 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_86
timestamp 1621261055
transform 1 0 9408 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_92
timestamp 1621261055
transform 1 0 9984 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_100
timestamp 1621261055
transform 1 0 10752 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _017_
timestamp 1621261055
transform 1 0 12576 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_858
timestamp 1621261055
transform 1 0 11712 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_108
timestamp 1621261055
transform 1 0 11520 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_111
timestamp 1621261055
transform 1 0 11808 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_122
timestamp 1621261055
transform 1 0 12864 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_130
timestamp 1621261055
transform 1 0 13632 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_138
timestamp 1621261055
transform 1 0 14400 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_146
timestamp 1621261055
transform 1 0 15168 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_859
timestamp 1621261055
transform 1 0 16992 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_154
timestamp 1621261055
transform 1 0 15936 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_162
timestamp 1621261055
transform 1 0 16704 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_164
timestamp 1621261055
transform 1 0 16896 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_166
timestamp 1621261055
transform 1 0 17088 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_174
timestamp 1621261055
transform 1 0 17856 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_182
timestamp 1621261055
transform 1 0 18624 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_190
timestamp 1621261055
transform 1 0 19392 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_198
timestamp 1621261055
transform 1 0 20160 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_206
timestamp 1621261055
transform 1 0 20928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_860
timestamp 1621261055
transform 1 0 22272 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_214
timestamp 1621261055
transform 1 0 21696 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_218
timestamp 1621261055
transform 1 0 22080 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_221
timestamp 1621261055
transform 1 0 22368 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_229
timestamp 1621261055
transform 1 0 23136 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_237
timestamp 1621261055
transform 1 0 23904 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_245
timestamp 1621261055
transform 1 0 24672 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_253
timestamp 1621261055
transform 1 0 25440 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_261
timestamp 1621261055
transform 1 0 26208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_269
timestamp 1621261055
transform 1 0 26976 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_273
timestamp 1621261055
transform 1 0 27360 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_861
timestamp 1621261055
transform 1 0 27552 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_276
timestamp 1621261055
transform 1 0 27648 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_284
timestamp 1621261055
transform 1 0 28416 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_292
timestamp 1621261055
transform 1 0 29184 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_300
timestamp 1621261055
transform 1 0 29952 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_308
timestamp 1621261055
transform 1 0 30720 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_862
timestamp 1621261055
transform 1 0 32832 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_316
timestamp 1621261055
transform 1 0 31488 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_324
timestamp 1621261055
transform 1 0 32256 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_328
timestamp 1621261055
transform 1 0 32640 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_331
timestamp 1621261055
transform 1 0 32928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_339
timestamp 1621261055
transform 1 0 33696 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_347
timestamp 1621261055
transform 1 0 34464 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_355
timestamp 1621261055
transform 1 0 35232 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_363
timestamp 1621261055
transform 1 0 36000 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_371
timestamp 1621261055
transform 1 0 36768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_863
timestamp 1621261055
transform 1 0 38112 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_379
timestamp 1621261055
transform 1 0 37536 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_383
timestamp 1621261055
transform 1 0 37920 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_386
timestamp 1621261055
transform 1 0 38208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_394
timestamp 1621261055
transform 1 0 38976 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_402
timestamp 1621261055
transform 1 0 39744 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_410
timestamp 1621261055
transform 1 0 40512 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_418
timestamp 1621261055
transform 1 0 41280 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_864
timestamp 1621261055
transform 1 0 43392 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_426
timestamp 1621261055
transform 1 0 42048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_434
timestamp 1621261055
transform 1 0 42816 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_438
timestamp 1621261055
transform 1 0 43200 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_441
timestamp 1621261055
transform 1 0 43488 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_449
timestamp 1621261055
transform 1 0 44256 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_457
timestamp 1621261055
transform 1 0 45024 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_465
timestamp 1621261055
transform 1 0 45792 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_473
timestamp 1621261055
transform 1 0 46560 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_481
timestamp 1621261055
transform 1 0 47328 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_865
timestamp 1621261055
transform 1 0 48672 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_489
timestamp 1621261055
transform 1 0 48096 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_493
timestamp 1621261055
transform 1 0 48480 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_496
timestamp 1621261055
transform 1 0 48768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_504
timestamp 1621261055
transform 1 0 49536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_512
timestamp 1621261055
transform 1 0 50304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_520
timestamp 1621261055
transform 1 0 51072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_528
timestamp 1621261055
transform 1 0 51840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_536
timestamp 1621261055
transform 1 0 52608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_544
timestamp 1621261055
transform 1 0 53376 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_866
timestamp 1621261055
transform 1 0 53952 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_548
timestamp 1621261055
transform 1 0 53760 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_551
timestamp 1621261055
transform 1 0 54048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_559
timestamp 1621261055
transform 1 0 54816 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_567
timestamp 1621261055
transform 1 0 55584 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_575
timestamp 1621261055
transform 1 0 56352 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_583
timestamp 1621261055
transform 1 0 57120 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_131
timestamp 1621261055
transform -1 0 58848 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_65_591
timestamp 1621261055
transform 1 0 57888 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_595
timestamp 1621261055
transform 1 0 58272 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_132
timestamp 1621261055
transform 1 0 1152 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_66_4
timestamp 1621261055
transform 1 0 1536 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_12
timestamp 1621261055
transform 1 0 2304 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_20
timestamp 1621261055
transform 1 0 3072 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_867
timestamp 1621261055
transform 1 0 3840 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_29
timestamp 1621261055
transform 1 0 3936 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_37
timestamp 1621261055
transform 1 0 4704 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _026_
timestamp 1621261055
transform 1 0 6528 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_66_45
timestamp 1621261055
transform 1 0 5472 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_53
timestamp 1621261055
transform 1 0 6240 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_66_55
timestamp 1621261055
transform 1 0 6432 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_59
timestamp 1621261055
transform 1 0 6816 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_868
timestamp 1621261055
transform 1 0 9120 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_67
timestamp 1621261055
transform 1 0 7584 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_75
timestamp 1621261055
transform 1 0 8352 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_84
timestamp 1621261055
transform 1 0 9216 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_92
timestamp 1621261055
transform 1 0 9984 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_100
timestamp 1621261055
transform 1 0 10752 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_108
timestamp 1621261055
transform 1 0 11520 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_116
timestamp 1621261055
transform 1 0 12288 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_124
timestamp 1621261055
transform 1 0 13056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_869
timestamp 1621261055
transform 1 0 14400 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_132
timestamp 1621261055
transform 1 0 13824 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_136
timestamp 1621261055
transform 1 0 14208 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_139
timestamp 1621261055
transform 1 0 14496 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_147
timestamp 1621261055
transform 1 0 15264 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_155
timestamp 1621261055
transform 1 0 16032 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_163
timestamp 1621261055
transform 1 0 16800 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_171
timestamp 1621261055
transform 1 0 17568 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_179
timestamp 1621261055
transform 1 0 18336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_187
timestamp 1621261055
transform 1 0 19104 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_870
timestamp 1621261055
transform 1 0 19680 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_191
timestamp 1621261055
transform 1 0 19488 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_194
timestamp 1621261055
transform 1 0 19776 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_202
timestamp 1621261055
transform 1 0 20544 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_210
timestamp 1621261055
transform 1 0 21312 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_218
timestamp 1621261055
transform 1 0 22080 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_226
timestamp 1621261055
transform 1 0 22848 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_230
timestamp 1621261055
transform 1 0 23232 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _133_
timestamp 1621261055
transform 1 0 23712 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_871
timestamp 1621261055
transform 1 0 24960 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_182
timestamp 1621261055
transform 1 0 23520 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_66_232
timestamp 1621261055
transform 1 0 23424 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_238
timestamp 1621261055
transform 1 0 24000 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_246
timestamp 1621261055
transform 1 0 24768 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_249
timestamp 1621261055
transform 1 0 25056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_257
timestamp 1621261055
transform 1 0 25824 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_265
timestamp 1621261055
transform 1 0 26592 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_273
timestamp 1621261055
transform 1 0 27360 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_281
timestamp 1621261055
transform 1 0 28128 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_289
timestamp 1621261055
transform 1 0 28896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_872
timestamp 1621261055
transform 1 0 30240 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_297
timestamp 1621261055
transform 1 0 29664 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_301
timestamp 1621261055
transform 1 0 30048 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_304
timestamp 1621261055
transform 1 0 30336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_312
timestamp 1621261055
transform 1 0 31104 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_320
timestamp 1621261055
transform 1 0 31872 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_328
timestamp 1621261055
transform 1 0 32640 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_336
timestamp 1621261055
transform 1 0 33408 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_344
timestamp 1621261055
transform 1 0 34176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_352
timestamp 1621261055
transform 1 0 34944 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_356
timestamp 1621261055
transform 1 0 35328 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_873
timestamp 1621261055
transform 1 0 35520 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_359
timestamp 1621261055
transform 1 0 35616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_367
timestamp 1621261055
transform 1 0 36384 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_375
timestamp 1621261055
transform 1 0 37152 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_383
timestamp 1621261055
transform 1 0 37920 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_391
timestamp 1621261055
transform 1 0 38688 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_399
timestamp 1621261055
transform 1 0 39456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_874
timestamp 1621261055
transform 1 0 40800 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_407
timestamp 1621261055
transform 1 0 40224 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_411
timestamp 1621261055
transform 1 0 40608 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_414
timestamp 1621261055
transform 1 0 40896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_422
timestamp 1621261055
transform 1 0 41664 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_430
timestamp 1621261055
transform 1 0 42432 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_438
timestamp 1621261055
transform 1 0 43200 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_446
timestamp 1621261055
transform 1 0 43968 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_454
timestamp 1621261055
transform 1 0 44736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_462
timestamp 1621261055
transform 1 0 45504 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_875
timestamp 1621261055
transform 1 0 46080 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_466
timestamp 1621261055
transform 1 0 45888 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_469
timestamp 1621261055
transform 1 0 46176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_477
timestamp 1621261055
transform 1 0 46944 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_485
timestamp 1621261055
transform 1 0 47712 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_493
timestamp 1621261055
transform 1 0 48480 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_501
timestamp 1621261055
transform 1 0 49248 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_876
timestamp 1621261055
transform 1 0 51360 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_509
timestamp 1621261055
transform 1 0 50016 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_517
timestamp 1621261055
transform 1 0 50784 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_521
timestamp 1621261055
transform 1 0 51168 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_524
timestamp 1621261055
transform 1 0 51456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_532
timestamp 1621261055
transform 1 0 52224 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_540
timestamp 1621261055
transform 1 0 52992 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_548
timestamp 1621261055
transform 1 0 53760 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_556
timestamp 1621261055
transform 1 0 54528 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_564
timestamp 1621261055
transform 1 0 55296 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_877
timestamp 1621261055
transform 1 0 56640 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_572
timestamp 1621261055
transform 1 0 56064 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_576
timestamp 1621261055
transform 1 0 56448 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_579
timestamp 1621261055
transform 1 0 56736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_587
timestamp 1621261055
transform 1 0 57504 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_133
timestamp 1621261055
transform -1 0 58848 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_595
timestamp 1621261055
transform 1 0 58272 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_134
timestamp 1621261055
transform 1 0 1152 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_67_4
timestamp 1621261055
transform 1 0 1536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_12
timestamp 1621261055
transform 1 0 2304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_20
timestamp 1621261055
transform 1 0 3072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_28
timestamp 1621261055
transform 1 0 3840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_36
timestamp 1621261055
transform 1 0 4608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_878
timestamp 1621261055
transform 1 0 6432 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_44
timestamp 1621261055
transform 1 0 5376 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_52
timestamp 1621261055
transform 1 0 6144 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_54
timestamp 1621261055
transform 1 0 6336 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_56
timestamp 1621261055
transform 1 0 6528 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_64
timestamp 1621261055
transform 1 0 7296 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_72
timestamp 1621261055
transform 1 0 8064 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_80
timestamp 1621261055
transform 1 0 8832 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_88
timestamp 1621261055
transform 1 0 9600 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_96
timestamp 1621261055
transform 1 0 10368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_104
timestamp 1621261055
transform 1 0 11136 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_879
timestamp 1621261055
transform 1 0 11712 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_108
timestamp 1621261055
transform 1 0 11520 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_111
timestamp 1621261055
transform 1 0 11808 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_119
timestamp 1621261055
transform 1 0 12576 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_127
timestamp 1621261055
transform 1 0 13344 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_135
timestamp 1621261055
transform 1 0 14112 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_143
timestamp 1621261055
transform 1 0 14880 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_880
timestamp 1621261055
transform 1 0 16992 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_151
timestamp 1621261055
transform 1 0 15648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_159
timestamp 1621261055
transform 1 0 16416 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_163
timestamp 1621261055
transform 1 0 16800 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_166
timestamp 1621261055
transform 1 0 17088 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_174
timestamp 1621261055
transform 1 0 17856 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_182
timestamp 1621261055
transform 1 0 18624 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_190
timestamp 1621261055
transform 1 0 19392 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_198
timestamp 1621261055
transform 1 0 20160 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_206
timestamp 1621261055
transform 1 0 20928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_881
timestamp 1621261055
transform 1 0 22272 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_214
timestamp 1621261055
transform 1 0 21696 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_218
timestamp 1621261055
transform 1 0 22080 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_221
timestamp 1621261055
transform 1 0 22368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_229
timestamp 1621261055
transform 1 0 23136 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_237
timestamp 1621261055
transform 1 0 23904 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_245
timestamp 1621261055
transform 1 0 24672 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_253
timestamp 1621261055
transform 1 0 25440 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_261
timestamp 1621261055
transform 1 0 26208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_269
timestamp 1621261055
transform 1 0 26976 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_273
timestamp 1621261055
transform 1 0 27360 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_882
timestamp 1621261055
transform 1 0 27552 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_276
timestamp 1621261055
transform 1 0 27648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_284
timestamp 1621261055
transform 1 0 28416 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_292
timestamp 1621261055
transform 1 0 29184 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_300
timestamp 1621261055
transform 1 0 29952 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_308
timestamp 1621261055
transform 1 0 30720 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_883
timestamp 1621261055
transform 1 0 32832 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_316
timestamp 1621261055
transform 1 0 31488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_324
timestamp 1621261055
transform 1 0 32256 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_328
timestamp 1621261055
transform 1 0 32640 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_331
timestamp 1621261055
transform 1 0 32928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _112_
timestamp 1621261055
transform -1 0 34944 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_174
timestamp 1621261055
transform -1 0 34656 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_339
timestamp 1621261055
transform 1 0 33696 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_352
timestamp 1621261055
transform 1 0 34944 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_360
timestamp 1621261055
transform 1 0 35712 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_368
timestamp 1621261055
transform 1 0 36480 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_376
timestamp 1621261055
transform 1 0 37248 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_884
timestamp 1621261055
transform 1 0 38112 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_67_384
timestamp 1621261055
transform 1 0 38016 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_386
timestamp 1621261055
transform 1 0 38208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_394
timestamp 1621261055
transform 1 0 38976 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_402
timestamp 1621261055
transform 1 0 39744 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_410
timestamp 1621261055
transform 1 0 40512 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_418
timestamp 1621261055
transform 1 0 41280 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_885
timestamp 1621261055
transform 1 0 43392 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_426
timestamp 1621261055
transform 1 0 42048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_434
timestamp 1621261055
transform 1 0 42816 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_438
timestamp 1621261055
transform 1 0 43200 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_441
timestamp 1621261055
transform 1 0 43488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_449
timestamp 1621261055
transform 1 0 44256 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_457
timestamp 1621261055
transform 1 0 45024 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_465
timestamp 1621261055
transform 1 0 45792 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_473
timestamp 1621261055
transform 1 0 46560 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_481
timestamp 1621261055
transform 1 0 47328 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_886
timestamp 1621261055
transform 1 0 48672 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_489
timestamp 1621261055
transform 1 0 48096 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_493
timestamp 1621261055
transform 1 0 48480 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_496
timestamp 1621261055
transform 1 0 48768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_504
timestamp 1621261055
transform 1 0 49536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_512
timestamp 1621261055
transform 1 0 50304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_520
timestamp 1621261055
transform 1 0 51072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_528
timestamp 1621261055
transform 1 0 51840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_536
timestamp 1621261055
transform 1 0 52608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_544
timestamp 1621261055
transform 1 0 53376 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_887
timestamp 1621261055
transform 1 0 53952 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_548
timestamp 1621261055
transform 1 0 53760 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_551
timestamp 1621261055
transform 1 0 54048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_559
timestamp 1621261055
transform 1 0 54816 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_567
timestamp 1621261055
transform 1 0 55584 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_575
timestamp 1621261055
transform 1 0 56352 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_583
timestamp 1621261055
transform 1 0 57120 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_135
timestamp 1621261055
transform -1 0 58848 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_67_591
timestamp 1621261055
transform 1 0 57888 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_595
timestamp 1621261055
transform 1 0 58272 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_136
timestamp 1621261055
transform 1 0 1152 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_4
timestamp 1621261055
transform 1 0 1536 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_12
timestamp 1621261055
transform 1 0 2304 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_20
timestamp 1621261055
transform 1 0 3072 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _182_
timestamp 1621261055
transform -1 0 4704 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_888
timestamp 1621261055
transform 1 0 3840 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_206
timestamp 1621261055
transform -1 0 4416 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_29
timestamp 1621261055
transform 1 0 3936 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_68_31
timestamp 1621261055
transform 1 0 4128 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_37
timestamp 1621261055
transform 1 0 4704 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_45
timestamp 1621261055
transform 1 0 5472 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_53
timestamp 1621261055
transform 1 0 6240 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_61
timestamp 1621261055
transform 1 0 7008 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_889
timestamp 1621261055
transform 1 0 9120 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_69
timestamp 1621261055
transform 1 0 7776 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_77
timestamp 1621261055
transform 1 0 8544 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_81
timestamp 1621261055
transform 1 0 8928 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_84
timestamp 1621261055
transform 1 0 9216 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_92
timestamp 1621261055
transform 1 0 9984 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_100
timestamp 1621261055
transform 1 0 10752 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_108
timestamp 1621261055
transform 1 0 11520 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_116
timestamp 1621261055
transform 1 0 12288 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_124
timestamp 1621261055
transform 1 0 13056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_890
timestamp 1621261055
transform 1 0 14400 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_132
timestamp 1621261055
transform 1 0 13824 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_136
timestamp 1621261055
transform 1 0 14208 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_139
timestamp 1621261055
transform 1 0 14496 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_147
timestamp 1621261055
transform 1 0 15264 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_155
timestamp 1621261055
transform 1 0 16032 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_163
timestamp 1621261055
transform 1 0 16800 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_171
timestamp 1621261055
transform 1 0 17568 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_179
timestamp 1621261055
transform 1 0 18336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_187
timestamp 1621261055
transform 1 0 19104 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_891
timestamp 1621261055
transform 1 0 19680 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_191
timestamp 1621261055
transform 1 0 19488 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_194
timestamp 1621261055
transform 1 0 19776 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_202
timestamp 1621261055
transform 1 0 20544 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_210
timestamp 1621261055
transform 1 0 21312 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_218
timestamp 1621261055
transform 1 0 22080 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_226
timestamp 1621261055
transform 1 0 22848 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_892
timestamp 1621261055
transform 1 0 24960 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_234
timestamp 1621261055
transform 1 0 23616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_242
timestamp 1621261055
transform 1 0 24384 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_246
timestamp 1621261055
transform 1 0 24768 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_249
timestamp 1621261055
transform 1 0 25056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_257
timestamp 1621261055
transform 1 0 25824 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_265
timestamp 1621261055
transform 1 0 26592 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_273
timestamp 1621261055
transform 1 0 27360 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_281
timestamp 1621261055
transform 1 0 28128 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_289
timestamp 1621261055
transform 1 0 28896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_893
timestamp 1621261055
transform 1 0 30240 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_297
timestamp 1621261055
transform 1 0 29664 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_301
timestamp 1621261055
transform 1 0 30048 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_304
timestamp 1621261055
transform 1 0 30336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_312
timestamp 1621261055
transform 1 0 31104 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_320
timestamp 1621261055
transform 1 0 31872 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_328
timestamp 1621261055
transform 1 0 32640 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_336
timestamp 1621261055
transform 1 0 33408 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_344
timestamp 1621261055
transform 1 0 34176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_352
timestamp 1621261055
transform 1 0 34944 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_356
timestamp 1621261055
transform 1 0 35328 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_894
timestamp 1621261055
transform 1 0 35520 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_359
timestamp 1621261055
transform 1 0 35616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_367
timestamp 1621261055
transform 1 0 36384 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_375
timestamp 1621261055
transform 1 0 37152 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_383
timestamp 1621261055
transform 1 0 37920 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_391
timestamp 1621261055
transform 1 0 38688 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_399
timestamp 1621261055
transform 1 0 39456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _009_
timestamp 1621261055
transform 1 0 41280 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_895
timestamp 1621261055
transform 1 0 40800 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_407
timestamp 1621261055
transform 1 0 40224 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_411
timestamp 1621261055
transform 1 0 40608 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_68_414
timestamp 1621261055
transform 1 0 40896 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_421
timestamp 1621261055
transform 1 0 41568 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_429
timestamp 1621261055
transform 1 0 42336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_437
timestamp 1621261055
transform 1 0 43104 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_445
timestamp 1621261055
transform 1 0 43872 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_453
timestamp 1621261055
transform 1 0 44640 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_461
timestamp 1621261055
transform 1 0 45408 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_896
timestamp 1621261055
transform 1 0 46080 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_465
timestamp 1621261055
transform 1 0 45792 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_68_467
timestamp 1621261055
transform 1 0 45984 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_469
timestamp 1621261055
transform 1 0 46176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_477
timestamp 1621261055
transform 1 0 46944 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_485
timestamp 1621261055
transform 1 0 47712 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_493
timestamp 1621261055
transform 1 0 48480 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_501
timestamp 1621261055
transform 1 0 49248 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_897
timestamp 1621261055
transform 1 0 51360 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_509
timestamp 1621261055
transform 1 0 50016 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_517
timestamp 1621261055
transform 1 0 50784 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_521
timestamp 1621261055
transform 1 0 51168 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_524
timestamp 1621261055
transform 1 0 51456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _213_
timestamp 1621261055
transform -1 0 53088 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_232
timestamp 1621261055
transform -1 0 52800 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_68_532
timestamp 1621261055
transform 1 0 52224 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_541
timestamp 1621261055
transform 1 0 53088 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_549
timestamp 1621261055
transform 1 0 53856 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_557
timestamp 1621261055
transform 1 0 54624 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_565
timestamp 1621261055
transform 1 0 55392 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_898
timestamp 1621261055
transform 1 0 56640 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_573
timestamp 1621261055
transform 1 0 56160 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_68_577
timestamp 1621261055
transform 1 0 56544 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_579
timestamp 1621261055
transform 1 0 56736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_587
timestamp 1621261055
transform 1 0 57504 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_137
timestamp 1621261055
transform -1 0 58848 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_595
timestamp 1621261055
transform 1 0 58272 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_138
timestamp 1621261055
transform 1 0 1152 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_140
timestamp 1621261055
transform 1 0 1152 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_154
timestamp 1621261055
transform 1 0 3168 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_4
timestamp 1621261055
transform 1 0 1536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_12
timestamp 1621261055
transform 1 0 2304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_20
timestamp 1621261055
transform 1 0 3072 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_4
timestamp 1621261055
transform 1 0 1536 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_12
timestamp 1621261055
transform 1 0 2304 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_20
timestamp 1621261055
transform 1 0 3072 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _101_
timestamp 1621261055
transform 1 0 3360 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_909
timestamp 1621261055
transform 1 0 3840 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_26
timestamp 1621261055
transform 1 0 3648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_34
timestamp 1621261055
transform 1 0 4416 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_42
timestamp 1621261055
transform 1 0 5184 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_29
timestamp 1621261055
transform 1 0 3936 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_37
timestamp 1621261055
transform 1 0 4704 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_899
timestamp 1621261055
transform 1 0 6432 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_50
timestamp 1621261055
transform 1 0 5952 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_69_54
timestamp 1621261055
transform 1 0 6336 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_56
timestamp 1621261055
transform 1 0 6528 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_45
timestamp 1621261055
transform 1 0 5472 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_53
timestamp 1621261055
transform 1 0 6240 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_61
timestamp 1621261055
transform 1 0 7008 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_910
timestamp 1621261055
transform 1 0 9120 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_64
timestamp 1621261055
transform 1 0 7296 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_72
timestamp 1621261055
transform 1 0 8064 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_80
timestamp 1621261055
transform 1 0 8832 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_69
timestamp 1621261055
transform 1 0 7776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_77
timestamp 1621261055
transform 1 0 8544 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_81
timestamp 1621261055
transform 1 0 8928 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_84
timestamp 1621261055
transform 1 0 9216 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_88
timestamp 1621261055
transform 1 0 9600 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_96
timestamp 1621261055
transform 1 0 10368 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_104
timestamp 1621261055
transform 1 0 11136 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_92
timestamp 1621261055
transform 1 0 9984 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_100
timestamp 1621261055
transform 1 0 10752 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _184_
timestamp 1621261055
transform -1 0 12192 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_900
timestamp 1621261055
transform 1 0 11712 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_220
timestamp 1621261055
transform -1 0 11904 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_108
timestamp 1621261055
transform 1 0 11520 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_111
timestamp 1621261055
transform 1 0 11808 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_119
timestamp 1621261055
transform 1 0 12576 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_108
timestamp 1621261055
transform 1 0 11520 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_115
timestamp 1621261055
transform 1 0 12192 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_123
timestamp 1621261055
transform 1 0 12960 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_911
timestamp 1621261055
transform 1 0 14400 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_127
timestamp 1621261055
transform 1 0 13344 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_135
timestamp 1621261055
transform 1 0 14112 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_143
timestamp 1621261055
transform 1 0 14880 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_131
timestamp 1621261055
transform 1 0 13728 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_135
timestamp 1621261055
transform 1 0 14112 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_70_137
timestamp 1621261055
transform 1 0 14304 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_139
timestamp 1621261055
transform 1 0 14496 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_147
timestamp 1621261055
transform 1 0 15264 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _212_
timestamp 1621261055
transform -1 0 15936 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_901
timestamp 1621261055
transform 1 0 16992 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_230
timestamp 1621261055
transform -1 0 15648 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_151
timestamp 1621261055
transform 1 0 15648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_159
timestamp 1621261055
transform 1 0 16416 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_163
timestamp 1621261055
transform 1 0 16800 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_166
timestamp 1621261055
transform 1 0 17088 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_154
timestamp 1621261055
transform 1 0 15936 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_162
timestamp 1621261055
transform 1 0 16704 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _027_
timestamp 1621261055
transform 1 0 18336 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_69_174
timestamp 1621261055
transform 1 0 17856 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_69_178
timestamp 1621261055
transform 1 0 18240 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_182
timestamp 1621261055
transform 1 0 18624 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_170
timestamp 1621261055
transform 1 0 17472 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_178
timestamp 1621261055
transform 1 0 18240 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_186
timestamp 1621261055
transform 1 0 19008 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_912
timestamp 1621261055
transform 1 0 19680 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_190
timestamp 1621261055
transform 1 0 19392 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_198
timestamp 1621261055
transform 1 0 20160 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_206
timestamp 1621261055
transform 1 0 20928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_190
timestamp 1621261055
transform 1 0 19392 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_70_192
timestamp 1621261055
transform 1 0 19584 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_194
timestamp 1621261055
transform 1 0 19776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_202
timestamp 1621261055
transform 1 0 20544 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_210
timestamp 1621261055
transform 1 0 21312 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _010_
timestamp 1621261055
transform 1 0 22752 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_902
timestamp 1621261055
transform 1 0 22272 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_214
timestamp 1621261055
transform 1 0 21696 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_218
timestamp 1621261055
transform 1 0 22080 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_221
timestamp 1621261055
transform 1 0 22368 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_228
timestamp 1621261055
transform 1 0 23040 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_218
timestamp 1621261055
transform 1 0 22080 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_226
timestamp 1621261055
transform 1 0 22848 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_913
timestamp 1621261055
transform 1 0 24960 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_236
timestamp 1621261055
transform 1 0 23808 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_244
timestamp 1621261055
transform 1 0 24576 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_252
timestamp 1621261055
transform 1 0 25344 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_234
timestamp 1621261055
transform 1 0 23616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_242
timestamp 1621261055
transform 1 0 24384 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_246
timestamp 1621261055
transform 1 0 24768 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_249
timestamp 1621261055
transform 1 0 25056 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_260
timestamp 1621261055
transform 1 0 26112 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_268
timestamp 1621261055
transform 1 0 26880 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_272
timestamp 1621261055
transform 1 0 27264 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_257
timestamp 1621261055
transform 1 0 25824 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_265
timestamp 1621261055
transform 1 0 26592 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_273
timestamp 1621261055
transform 1 0 27360 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_903
timestamp 1621261055
transform 1 0 27552 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_69_274
timestamp 1621261055
transform 1 0 27456 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_276
timestamp 1621261055
transform 1 0 27648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_284
timestamp 1621261055
transform 1 0 28416 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_292
timestamp 1621261055
transform 1 0 29184 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_281
timestamp 1621261055
transform 1 0 28128 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_289
timestamp 1621261055
transform 1 0 28896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_914
timestamp 1621261055
transform 1 0 30240 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_300
timestamp 1621261055
transform 1 0 29952 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_308
timestamp 1621261055
transform 1 0 30720 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_297
timestamp 1621261055
transform 1 0 29664 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_301
timestamp 1621261055
transform 1 0 30048 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_304
timestamp 1621261055
transform 1 0 30336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_312
timestamp 1621261055
transform 1 0 31104 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_904
timestamp 1621261055
transform 1 0 32832 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_316
timestamp 1621261055
transform 1 0 31488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_324
timestamp 1621261055
transform 1 0 32256 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_328
timestamp 1621261055
transform 1 0 32640 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_331
timestamp 1621261055
transform 1 0 32928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_320
timestamp 1621261055
transform 1 0 31872 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_328
timestamp 1621261055
transform 1 0 32640 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_336
timestamp 1621261055
transform 1 0 33408 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_339
timestamp 1621261055
transform 1 0 33696 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_347
timestamp 1621261055
transform 1 0 34464 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_355
timestamp 1621261055
transform 1 0 35232 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_344
timestamp 1621261055
transform 1 0 34176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_352
timestamp 1621261055
transform 1 0 34944 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_356
timestamp 1621261055
transform 1 0 35328 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_915
timestamp 1621261055
transform 1 0 35520 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_363
timestamp 1621261055
transform 1 0 36000 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_371
timestamp 1621261055
transform 1 0 36768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_359
timestamp 1621261055
transform 1 0 35616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_367
timestamp 1621261055
transform 1 0 36384 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_375
timestamp 1621261055
transform 1 0 37152 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_905
timestamp 1621261055
transform 1 0 38112 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_379
timestamp 1621261055
transform 1 0 37536 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_383
timestamp 1621261055
transform 1 0 37920 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_386
timestamp 1621261055
transform 1 0 38208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_394
timestamp 1621261055
transform 1 0 38976 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_383
timestamp 1621261055
transform 1 0 37920 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_391
timestamp 1621261055
transform 1 0 38688 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_399
timestamp 1621261055
transform 1 0 39456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_916
timestamp 1621261055
transform 1 0 40800 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_402
timestamp 1621261055
transform 1 0 39744 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_410
timestamp 1621261055
transform 1 0 40512 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_418
timestamp 1621261055
transform 1 0 41280 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_407
timestamp 1621261055
transform 1 0 40224 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_411
timestamp 1621261055
transform 1 0 40608 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_414
timestamp 1621261055
transform 1 0 40896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_906
timestamp 1621261055
transform 1 0 43392 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_426
timestamp 1621261055
transform 1 0 42048 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_434
timestamp 1621261055
transform 1 0 42816 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_438
timestamp 1621261055
transform 1 0 43200 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_441
timestamp 1621261055
transform 1 0 43488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_422
timestamp 1621261055
transform 1 0 41664 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_430
timestamp 1621261055
transform 1 0 42432 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_438
timestamp 1621261055
transform 1 0 43200 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_449
timestamp 1621261055
transform 1 0 44256 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_457
timestamp 1621261055
transform 1 0 45024 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_446
timestamp 1621261055
transform 1 0 43968 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_454
timestamp 1621261055
transform 1 0 44736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_462
timestamp 1621261055
transform 1 0 45504 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_917
timestamp 1621261055
transform 1 0 46080 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_465
timestamp 1621261055
transform 1 0 45792 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_473
timestamp 1621261055
transform 1 0 46560 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_481
timestamp 1621261055
transform 1 0 47328 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_466
timestamp 1621261055
transform 1 0 45888 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_469
timestamp 1621261055
transform 1 0 46176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_477
timestamp 1621261055
transform 1 0 46944 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_485
timestamp 1621261055
transform 1 0 47712 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_489
timestamp 1621261055
transform 1 0 48096 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_493
timestamp 1621261055
transform 1 0 48480 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_496
timestamp 1621261055
transform 1 0 48768 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_493
timestamp 1621261055
transform 1 0 48480 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_105
timestamp 1621261055
transform 1 0 48960 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_907
timestamp 1621261055
transform 1 0 48672 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _159_
timestamp 1621261055
transform 1 0 49152 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_501
timestamp 1621261055
transform 1 0 49248 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_503
timestamp 1621261055
transform 1 0 49440 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_918
timestamp 1621261055
transform 1 0 51360 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_511
timestamp 1621261055
transform 1 0 50208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_519
timestamp 1621261055
transform 1 0 50976 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_509
timestamp 1621261055
transform 1 0 50016 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_517
timestamp 1621261055
transform 1 0 50784 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_521
timestamp 1621261055
transform 1 0 51168 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_524
timestamp 1621261055
transform 1 0 51456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _214_
timestamp 1621261055
transform 1 0 52224 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_69_527
timestamp 1621261055
transform 1 0 51744 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_535
timestamp 1621261055
transform 1 0 52512 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_543
timestamp 1621261055
transform 1 0 53280 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_535
timestamp 1621261055
transform 1 0 52512 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_543
timestamp 1621261055
transform 1 0 53280 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_908
timestamp 1621261055
transform 1 0 53952 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_547
timestamp 1621261055
transform 1 0 53664 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_69_549
timestamp 1621261055
transform 1 0 53856 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_551
timestamp 1621261055
transform 1 0 54048 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_559
timestamp 1621261055
transform 1 0 54816 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_567
timestamp 1621261055
transform 1 0 55584 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_551
timestamp 1621261055
transform 1 0 54048 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_559
timestamp 1621261055
transform 1 0 54816 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_567
timestamp 1621261055
transform 1 0 55584 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_919
timestamp 1621261055
transform 1 0 56640 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_575
timestamp 1621261055
transform 1 0 56352 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_583
timestamp 1621261055
transform 1 0 57120 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_575
timestamp 1621261055
transform 1 0 56352 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_70_577
timestamp 1621261055
transform 1 0 56544 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_579
timestamp 1621261055
transform 1 0 56736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_587
timestamp 1621261055
transform 1 0 57504 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_139
timestamp 1621261055
transform -1 0 58848 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_141
timestamp 1621261055
transform -1 0 58848 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_69_591
timestamp 1621261055
transform 1 0 57888 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_595
timestamp 1621261055
transform 1 0 58272 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_595
timestamp 1621261055
transform 1 0 58272 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_142
timestamp 1621261055
transform 1 0 1152 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_71_4
timestamp 1621261055
transform 1 0 1536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_12
timestamp 1621261055
transform 1 0 2304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_20
timestamp 1621261055
transform 1 0 3072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_28
timestamp 1621261055
transform 1 0 3840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_36
timestamp 1621261055
transform 1 0 4608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_920
timestamp 1621261055
transform 1 0 6432 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_44
timestamp 1621261055
transform 1 0 5376 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_52
timestamp 1621261055
transform 1 0 6144 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_54
timestamp 1621261055
transform 1 0 6336 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_56
timestamp 1621261055
transform 1 0 6528 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_64
timestamp 1621261055
transform 1 0 7296 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_72
timestamp 1621261055
transform 1 0 8064 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_80
timestamp 1621261055
transform 1 0 8832 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_88
timestamp 1621261055
transform 1 0 9600 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_96
timestamp 1621261055
transform 1 0 10368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_104
timestamp 1621261055
transform 1 0 11136 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_921
timestamp 1621261055
transform 1 0 11712 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_108
timestamp 1621261055
transform 1 0 11520 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_111
timestamp 1621261055
transform 1 0 11808 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_119
timestamp 1621261055
transform 1 0 12576 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_127
timestamp 1621261055
transform 1 0 13344 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_135
timestamp 1621261055
transform 1 0 14112 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_143
timestamp 1621261055
transform 1 0 14880 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_922
timestamp 1621261055
transform 1 0 16992 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_151
timestamp 1621261055
transform 1 0 15648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_159
timestamp 1621261055
transform 1 0 16416 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_163
timestamp 1621261055
transform 1 0 16800 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_166
timestamp 1621261055
transform 1 0 17088 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_174
timestamp 1621261055
transform 1 0 17856 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_182
timestamp 1621261055
transform 1 0 18624 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_190
timestamp 1621261055
transform 1 0 19392 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_198
timestamp 1621261055
transform 1 0 20160 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_206
timestamp 1621261055
transform 1 0 20928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_923
timestamp 1621261055
transform 1 0 22272 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_214
timestamp 1621261055
transform 1 0 21696 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_218
timestamp 1621261055
transform 1 0 22080 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_221
timestamp 1621261055
transform 1 0 22368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_229
timestamp 1621261055
transform 1 0 23136 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_237
timestamp 1621261055
transform 1 0 23904 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_245
timestamp 1621261055
transform 1 0 24672 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_253
timestamp 1621261055
transform 1 0 25440 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_261
timestamp 1621261055
transform 1 0 26208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_269
timestamp 1621261055
transform 1 0 26976 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_273
timestamp 1621261055
transform 1 0 27360 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_924
timestamp 1621261055
transform 1 0 27552 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_276
timestamp 1621261055
transform 1 0 27648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_284
timestamp 1621261055
transform 1 0 28416 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_292
timestamp 1621261055
transform 1 0 29184 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_300
timestamp 1621261055
transform 1 0 29952 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_308
timestamp 1621261055
transform 1 0 30720 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_925
timestamp 1621261055
transform 1 0 32832 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_316
timestamp 1621261055
transform 1 0 31488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_324
timestamp 1621261055
transform 1 0 32256 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_328
timestamp 1621261055
transform 1 0 32640 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_331
timestamp 1621261055
transform 1 0 32928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_339
timestamp 1621261055
transform 1 0 33696 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_347
timestamp 1621261055
transform 1 0 34464 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_355
timestamp 1621261055
transform 1 0 35232 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_363
timestamp 1621261055
transform 1 0 36000 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_371
timestamp 1621261055
transform 1 0 36768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _071_
timestamp 1621261055
transform -1 0 39744 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_926
timestamp 1621261055
transform 1 0 38112 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_130
timestamp 1621261055
transform -1 0 39456 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_71_379
timestamp 1621261055
transform 1 0 37536 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_383
timestamp 1621261055
transform 1 0 37920 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_386
timestamp 1621261055
transform 1 0 38208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_394
timestamp 1621261055
transform 1 0 38976 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_396
timestamp 1621261055
transform 1 0 39168 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_402
timestamp 1621261055
transform 1 0 39744 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_410
timestamp 1621261055
transform 1 0 40512 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_418
timestamp 1621261055
transform 1 0 41280 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_927
timestamp 1621261055
transform 1 0 43392 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_426
timestamp 1621261055
transform 1 0 42048 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_434
timestamp 1621261055
transform 1 0 42816 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_438
timestamp 1621261055
transform 1 0 43200 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_441
timestamp 1621261055
transform 1 0 43488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_449
timestamp 1621261055
transform 1 0 44256 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_457
timestamp 1621261055
transform 1 0 45024 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_465
timestamp 1621261055
transform 1 0 45792 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_473
timestamp 1621261055
transform 1 0 46560 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_481
timestamp 1621261055
transform 1 0 47328 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_928
timestamp 1621261055
transform 1 0 48672 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_489
timestamp 1621261055
transform 1 0 48096 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_493
timestamp 1621261055
transform 1 0 48480 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_496
timestamp 1621261055
transform 1 0 48768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_504
timestamp 1621261055
transform 1 0 49536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _024_
timestamp 1621261055
transform 1 0 51552 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_71_512
timestamp 1621261055
transform 1 0 50304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_520
timestamp 1621261055
transform 1 0 51072 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_71_524
timestamp 1621261055
transform 1 0 51456 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_528
timestamp 1621261055
transform 1 0 51840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_536
timestamp 1621261055
transform 1 0 52608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_544
timestamp 1621261055
transform 1 0 53376 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_929
timestamp 1621261055
transform 1 0 53952 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_548
timestamp 1621261055
transform 1 0 53760 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_551
timestamp 1621261055
transform 1 0 54048 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_559
timestamp 1621261055
transform 1 0 54816 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_567
timestamp 1621261055
transform 1 0 55584 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _093_
timestamp 1621261055
transform -1 0 57888 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_144
timestamp 1621261055
transform -1 0 57600 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_575
timestamp 1621261055
transform 1 0 56352 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_583
timestamp 1621261055
transform 1 0 57120 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_585
timestamp 1621261055
transform 1 0 57312 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_143
timestamp 1621261055
transform -1 0 58848 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_71_591
timestamp 1621261055
transform 1 0 57888 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_595
timestamp 1621261055
transform 1 0 58272 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_144
timestamp 1621261055
transform 1 0 1152 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_72_4
timestamp 1621261055
transform 1 0 1536 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_12
timestamp 1621261055
transform 1 0 2304 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_20
timestamp 1621261055
transform 1 0 3072 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_930
timestamp 1621261055
transform 1 0 3840 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_29
timestamp 1621261055
transform 1 0 3936 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_37
timestamp 1621261055
transform 1 0 4704 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_45
timestamp 1621261055
transform 1 0 5472 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_53
timestamp 1621261055
transform 1 0 6240 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_61
timestamp 1621261055
transform 1 0 7008 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_931
timestamp 1621261055
transform 1 0 9120 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_69
timestamp 1621261055
transform 1 0 7776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_77
timestamp 1621261055
transform 1 0 8544 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_81
timestamp 1621261055
transform 1 0 8928 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_84
timestamp 1621261055
transform 1 0 9216 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_92
timestamp 1621261055
transform 1 0 9984 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_100
timestamp 1621261055
transform 1 0 10752 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_108
timestamp 1621261055
transform 1 0 11520 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_116
timestamp 1621261055
transform 1 0 12288 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_124
timestamp 1621261055
transform 1 0 13056 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_932
timestamp 1621261055
transform 1 0 14400 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_132
timestamp 1621261055
transform 1 0 13824 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_136
timestamp 1621261055
transform 1 0 14208 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_139
timestamp 1621261055
transform 1 0 14496 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_147
timestamp 1621261055
transform 1 0 15264 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _141_
timestamp 1621261055
transform 1 0 15840 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_192
timestamp 1621261055
transform 1 0 15648 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_156
timestamp 1621261055
transform 1 0 16128 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_164
timestamp 1621261055
transform 1 0 16896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_172
timestamp 1621261055
transform 1 0 17664 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_180
timestamp 1621261055
transform 1 0 18432 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_188
timestamp 1621261055
transform 1 0 19200 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_933
timestamp 1621261055
transform 1 0 19680 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_72_192
timestamp 1621261055
transform 1 0 19584 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_194
timestamp 1621261055
transform 1 0 19776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_202
timestamp 1621261055
transform 1 0 20544 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_210
timestamp 1621261055
transform 1 0 21312 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_218
timestamp 1621261055
transform 1 0 22080 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_226
timestamp 1621261055
transform 1 0 22848 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_934
timestamp 1621261055
transform 1 0 24960 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_234
timestamp 1621261055
transform 1 0 23616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_242
timestamp 1621261055
transform 1 0 24384 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_246
timestamp 1621261055
transform 1 0 24768 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_249
timestamp 1621261055
transform 1 0 25056 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_257
timestamp 1621261055
transform 1 0 25824 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_265
timestamp 1621261055
transform 1 0 26592 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_273
timestamp 1621261055
transform 1 0 27360 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_281
timestamp 1621261055
transform 1 0 28128 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_289
timestamp 1621261055
transform 1 0 28896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_935
timestamp 1621261055
transform 1 0 30240 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_297
timestamp 1621261055
transform 1 0 29664 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_301
timestamp 1621261055
transform 1 0 30048 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_304
timestamp 1621261055
transform 1 0 30336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_312
timestamp 1621261055
transform 1 0 31104 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_320
timestamp 1621261055
transform 1 0 31872 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_328
timestamp 1621261055
transform 1 0 32640 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_336
timestamp 1621261055
transform 1 0 33408 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_344
timestamp 1621261055
transform 1 0 34176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_352
timestamp 1621261055
transform 1 0 34944 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_356
timestamp 1621261055
transform 1 0 35328 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_936
timestamp 1621261055
transform 1 0 35520 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_359
timestamp 1621261055
transform 1 0 35616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_367
timestamp 1621261055
transform 1 0 36384 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_375
timestamp 1621261055
transform 1 0 37152 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_383
timestamp 1621261055
transform 1 0 37920 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_391
timestamp 1621261055
transform 1 0 38688 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_399
timestamp 1621261055
transform 1 0 39456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_937
timestamp 1621261055
transform 1 0 40800 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_407
timestamp 1621261055
transform 1 0 40224 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_411
timestamp 1621261055
transform 1 0 40608 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_414
timestamp 1621261055
transform 1 0 40896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_422
timestamp 1621261055
transform 1 0 41664 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_430
timestamp 1621261055
transform 1 0 42432 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_438
timestamp 1621261055
transform 1 0 43200 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_446
timestamp 1621261055
transform 1 0 43968 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_454
timestamp 1621261055
transform 1 0 44736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_462
timestamp 1621261055
transform 1 0 45504 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_938
timestamp 1621261055
transform 1 0 46080 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_466
timestamp 1621261055
transform 1 0 45888 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_469
timestamp 1621261055
transform 1 0 46176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_477
timestamp 1621261055
transform 1 0 46944 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_485
timestamp 1621261055
transform 1 0 47712 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_493
timestamp 1621261055
transform 1 0 48480 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_501
timestamp 1621261055
transform 1 0 49248 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_939
timestamp 1621261055
transform 1 0 51360 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_509
timestamp 1621261055
transform 1 0 50016 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_517
timestamp 1621261055
transform 1 0 50784 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_521
timestamp 1621261055
transform 1 0 51168 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_524
timestamp 1621261055
transform 1 0 51456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_222
timestamp 1621261055
transform -1 0 53760 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_532
timestamp 1621261055
transform 1 0 52224 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_540
timestamp 1621261055
transform 1 0 52992 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_544
timestamp 1621261055
transform 1 0 53376 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _203_
timestamp 1621261055
transform -1 0 54048 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_72_551
timestamp 1621261055
transform 1 0 54048 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_559
timestamp 1621261055
transform 1 0 54816 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_567
timestamp 1621261055
transform 1 0 55584 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_940
timestamp 1621261055
transform 1 0 56640 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_575
timestamp 1621261055
transform 1 0 56352 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_72_577
timestamp 1621261055
transform 1 0 56544 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_579
timestamp 1621261055
transform 1 0 56736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_587
timestamp 1621261055
transform 1 0 57504 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_145
timestamp 1621261055
transform -1 0 58848 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_595
timestamp 1621261055
transform 1 0 58272 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_146
timestamp 1621261055
transform 1 0 1152 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_73_4
timestamp 1621261055
transform 1 0 1536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_12
timestamp 1621261055
transform 1 0 2304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_20
timestamp 1621261055
transform 1 0 3072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_28
timestamp 1621261055
transform 1 0 3840 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_36
timestamp 1621261055
transform 1 0 4608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_941
timestamp 1621261055
transform 1 0 6432 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_44
timestamp 1621261055
transform 1 0 5376 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_52
timestamp 1621261055
transform 1 0 6144 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_54
timestamp 1621261055
transform 1 0 6336 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_56
timestamp 1621261055
transform 1 0 6528 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_64
timestamp 1621261055
transform 1 0 7296 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_72
timestamp 1621261055
transform 1 0 8064 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_80
timestamp 1621261055
transform 1 0 8832 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _012_
timestamp 1621261055
transform 1 0 10272 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_73_88
timestamp 1621261055
transform 1 0 9600 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_92
timestamp 1621261055
transform 1 0 9984 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_94
timestamp 1621261055
transform 1 0 10176 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_98
timestamp 1621261055
transform 1 0 10560 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_942
timestamp 1621261055
transform 1 0 11712 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_106
timestamp 1621261055
transform 1 0 11328 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_73_111
timestamp 1621261055
transform 1 0 11808 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_119
timestamp 1621261055
transform 1 0 12576 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_127
timestamp 1621261055
transform 1 0 13344 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_135
timestamp 1621261055
transform 1 0 14112 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_143
timestamp 1621261055
transform 1 0 14880 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_943
timestamp 1621261055
transform 1 0 16992 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_151
timestamp 1621261055
transform 1 0 15648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_159
timestamp 1621261055
transform 1 0 16416 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_163
timestamp 1621261055
transform 1 0 16800 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_166
timestamp 1621261055
transform 1 0 17088 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_174
timestamp 1621261055
transform 1 0 17856 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_182
timestamp 1621261055
transform 1 0 18624 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_190
timestamp 1621261055
transform 1 0 19392 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_198
timestamp 1621261055
transform 1 0 20160 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_206
timestamp 1621261055
transform 1 0 20928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_944
timestamp 1621261055
transform 1 0 22272 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_214
timestamp 1621261055
transform 1 0 21696 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_218
timestamp 1621261055
transform 1 0 22080 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_221
timestamp 1621261055
transform 1 0 22368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_229
timestamp 1621261055
transform 1 0 23136 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_237
timestamp 1621261055
transform 1 0 23904 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_245
timestamp 1621261055
transform 1 0 24672 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_253
timestamp 1621261055
transform 1 0 25440 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_261
timestamp 1621261055
transform 1 0 26208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_269
timestamp 1621261055
transform 1 0 26976 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_273
timestamp 1621261055
transform 1 0 27360 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_945
timestamp 1621261055
transform 1 0 27552 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_276
timestamp 1621261055
transform 1 0 27648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_284
timestamp 1621261055
transform 1 0 28416 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_292
timestamp 1621261055
transform 1 0 29184 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_294
timestamp 1621261055
transform 1 0 29376 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _005_
timestamp 1621261055
transform 1 0 29472 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_73_298
timestamp 1621261055
transform 1 0 29760 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_306
timestamp 1621261055
transform 1 0 30528 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_314
timestamp 1621261055
transform 1 0 31296 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_946
timestamp 1621261055
transform 1 0 32832 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_322
timestamp 1621261055
transform 1 0 32064 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_331
timestamp 1621261055
transform 1 0 32928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_339
timestamp 1621261055
transform 1 0 33696 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_347
timestamp 1621261055
transform 1 0 34464 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_355
timestamp 1621261055
transform 1 0 35232 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_363
timestamp 1621261055
transform 1 0 36000 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_371
timestamp 1621261055
transform 1 0 36768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_947
timestamp 1621261055
transform 1 0 38112 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_379
timestamp 1621261055
transform 1 0 37536 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_383
timestamp 1621261055
transform 1 0 37920 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_386
timestamp 1621261055
transform 1 0 38208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_394
timestamp 1621261055
transform 1 0 38976 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_402
timestamp 1621261055
transform 1 0 39744 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_410
timestamp 1621261055
transform 1 0 40512 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_418
timestamp 1621261055
transform 1 0 41280 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_948
timestamp 1621261055
transform 1 0 43392 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_426
timestamp 1621261055
transform 1 0 42048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_434
timestamp 1621261055
transform 1 0 42816 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_438
timestamp 1621261055
transform 1 0 43200 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_441
timestamp 1621261055
transform 1 0 43488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_449
timestamp 1621261055
transform 1 0 44256 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_457
timestamp 1621261055
transform 1 0 45024 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_465
timestamp 1621261055
transform 1 0 45792 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_473
timestamp 1621261055
transform 1 0 46560 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_481
timestamp 1621261055
transform 1 0 47328 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_949
timestamp 1621261055
transform 1 0 48672 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_489
timestamp 1621261055
transform 1 0 48096 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_493
timestamp 1621261055
transform 1 0 48480 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_496
timestamp 1621261055
transform 1 0 48768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_504
timestamp 1621261055
transform 1 0 49536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_512
timestamp 1621261055
transform 1 0 50304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_520
timestamp 1621261055
transform 1 0 51072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_528
timestamp 1621261055
transform 1 0 51840 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_536
timestamp 1621261055
transform 1 0 52608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_544
timestamp 1621261055
transform 1 0 53376 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_950
timestamp 1621261055
transform 1 0 53952 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_548
timestamp 1621261055
transform 1 0 53760 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_551
timestamp 1621261055
transform 1 0 54048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_559
timestamp 1621261055
transform 1 0 54816 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_567
timestamp 1621261055
transform 1 0 55584 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_575
timestamp 1621261055
transform 1 0 56352 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_583
timestamp 1621261055
transform 1 0 57120 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_147
timestamp 1621261055
transform -1 0 58848 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_73_591
timestamp 1621261055
transform 1 0 57888 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_595
timestamp 1621261055
transform 1 0 58272 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _102_
timestamp 1621261055
transform 1 0 3168 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_148
timestamp 1621261055
transform 1 0 1152 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_157
timestamp 1621261055
transform 1 0 2976 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_4
timestamp 1621261055
transform 1 0 1536 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_12
timestamp 1621261055
transform 1 0 2304 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_16
timestamp 1621261055
transform 1 0 2688 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_74_18
timestamp 1621261055
transform 1 0 2880 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_951
timestamp 1621261055
transform 1 0 3840 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_24
timestamp 1621261055
transform 1 0 3456 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_74_29
timestamp 1621261055
transform 1 0 3936 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_37
timestamp 1621261055
transform 1 0 4704 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_45
timestamp 1621261055
transform 1 0 5472 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_53
timestamp 1621261055
transform 1 0 6240 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_61
timestamp 1621261055
transform 1 0 7008 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_952
timestamp 1621261055
transform 1 0 9120 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_69
timestamp 1621261055
transform 1 0 7776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_77
timestamp 1621261055
transform 1 0 8544 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_81
timestamp 1621261055
transform 1 0 8928 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_84
timestamp 1621261055
transform 1 0 9216 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_92
timestamp 1621261055
transform 1 0 9984 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_100
timestamp 1621261055
transform 1 0 10752 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_108
timestamp 1621261055
transform 1 0 11520 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_116
timestamp 1621261055
transform 1 0 12288 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_124
timestamp 1621261055
transform 1 0 13056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_953
timestamp 1621261055
transform 1 0 14400 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_132
timestamp 1621261055
transform 1 0 13824 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_136
timestamp 1621261055
transform 1 0 14208 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_139
timestamp 1621261055
transform 1 0 14496 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_147
timestamp 1621261055
transform 1 0 15264 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_155
timestamp 1621261055
transform 1 0 16032 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_163
timestamp 1621261055
transform 1 0 16800 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _109_
timestamp 1621261055
transform 1 0 18144 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_172
timestamp 1621261055
transform 1 0 17952 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_74_171
timestamp 1621261055
transform 1 0 17568 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_74_180
timestamp 1621261055
transform 1 0 18432 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_188
timestamp 1621261055
transform 1 0 19200 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_954
timestamp 1621261055
transform 1 0 19680 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_74_192
timestamp 1621261055
transform 1 0 19584 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_194
timestamp 1621261055
transform 1 0 19776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_202
timestamp 1621261055
transform 1 0 20544 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_210
timestamp 1621261055
transform 1 0 21312 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_218
timestamp 1621261055
transform 1 0 22080 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_226
timestamp 1621261055
transform 1 0 22848 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_955
timestamp 1621261055
transform 1 0 24960 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_234
timestamp 1621261055
transform 1 0 23616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_242
timestamp 1621261055
transform 1 0 24384 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_246
timestamp 1621261055
transform 1 0 24768 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_249
timestamp 1621261055
transform 1 0 25056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_257
timestamp 1621261055
transform 1 0 25824 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_265
timestamp 1621261055
transform 1 0 26592 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_273
timestamp 1621261055
transform 1 0 27360 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_281
timestamp 1621261055
transform 1 0 28128 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_289
timestamp 1621261055
transform 1 0 28896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_956
timestamp 1621261055
transform 1 0 30240 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_297
timestamp 1621261055
transform 1 0 29664 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_301
timestamp 1621261055
transform 1 0 30048 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_304
timestamp 1621261055
transform 1 0 30336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_312
timestamp 1621261055
transform 1 0 31104 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_320
timestamp 1621261055
transform 1 0 31872 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_328
timestamp 1621261055
transform 1 0 32640 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_336
timestamp 1621261055
transform 1 0 33408 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_344
timestamp 1621261055
transform 1 0 34176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_352
timestamp 1621261055
transform 1 0 34944 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_356
timestamp 1621261055
transform 1 0 35328 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_957
timestamp 1621261055
transform 1 0 35520 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_359
timestamp 1621261055
transform 1 0 35616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_367
timestamp 1621261055
transform 1 0 36384 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_375
timestamp 1621261055
transform 1 0 37152 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _057_
timestamp 1621261055
transform 1 0 37536 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_74_382
timestamp 1621261055
transform 1 0 37824 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_390
timestamp 1621261055
transform 1 0 38592 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_398
timestamp 1621261055
transform 1 0 39360 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _167_
timestamp 1621261055
transform 1 0 39840 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_958
timestamp 1621261055
transform 1 0 40800 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_112
timestamp 1621261055
transform 1 0 39648 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_74_400
timestamp 1621261055
transform 1 0 39552 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_406
timestamp 1621261055
transform 1 0 40128 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_410
timestamp 1621261055
transform 1 0 40512 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_74_412
timestamp 1621261055
transform 1 0 40704 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_414
timestamp 1621261055
transform 1 0 40896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_422
timestamp 1621261055
transform 1 0 41664 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_430
timestamp 1621261055
transform 1 0 42432 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_438
timestamp 1621261055
transform 1 0 43200 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_446
timestamp 1621261055
transform 1 0 43968 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_454
timestamp 1621261055
transform 1 0 44736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_462
timestamp 1621261055
transform 1 0 45504 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_959
timestamp 1621261055
transform 1 0 46080 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_466
timestamp 1621261055
transform 1 0 45888 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_469
timestamp 1621261055
transform 1 0 46176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_477
timestamp 1621261055
transform 1 0 46944 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_485
timestamp 1621261055
transform 1 0 47712 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_493
timestamp 1621261055
transform 1 0 48480 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_501
timestamp 1621261055
transform 1 0 49248 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_960
timestamp 1621261055
transform 1 0 51360 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_509
timestamp 1621261055
transform 1 0 50016 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_517
timestamp 1621261055
transform 1 0 50784 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_521
timestamp 1621261055
transform 1 0 51168 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_524
timestamp 1621261055
transform 1 0 51456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_532
timestamp 1621261055
transform 1 0 52224 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_540
timestamp 1621261055
transform 1 0 52992 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_548
timestamp 1621261055
transform 1 0 53760 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_556
timestamp 1621261055
transform 1 0 54528 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_564
timestamp 1621261055
transform 1 0 55296 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_961
timestamp 1621261055
transform 1 0 56640 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_572
timestamp 1621261055
transform 1 0 56064 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_576
timestamp 1621261055
transform 1 0 56448 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_579
timestamp 1621261055
transform 1 0 56736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_587
timestamp 1621261055
transform 1 0 57504 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_149
timestamp 1621261055
transform -1 0 58848 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_595
timestamp 1621261055
transform 1 0 58272 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_150
timestamp 1621261055
transform 1 0 1152 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_75_4
timestamp 1621261055
transform 1 0 1536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_12
timestamp 1621261055
transform 1 0 2304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_20
timestamp 1621261055
transform 1 0 3072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_28
timestamp 1621261055
transform 1 0 3840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_36
timestamp 1621261055
transform 1 0 4608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _158_
timestamp 1621261055
transform 1 0 7008 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_962
timestamp 1621261055
transform 1 0 6432 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_103
timestamp 1621261055
transform 1 0 6816 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_44
timestamp 1621261055
transform 1 0 5376 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_52
timestamp 1621261055
transform 1 0 6144 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_54
timestamp 1621261055
transform 1 0 6336 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_56
timestamp 1621261055
transform 1 0 6528 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_58
timestamp 1621261055
transform 1 0 6720 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_64
timestamp 1621261055
transform 1 0 7296 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_72
timestamp 1621261055
transform 1 0 8064 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_80
timestamp 1621261055
transform 1 0 8832 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_88
timestamp 1621261055
transform 1 0 9600 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_96
timestamp 1621261055
transform 1 0 10368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_104
timestamp 1621261055
transform 1 0 11136 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_963
timestamp 1621261055
transform 1 0 11712 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_108
timestamp 1621261055
transform 1 0 11520 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_111
timestamp 1621261055
transform 1 0 11808 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_119
timestamp 1621261055
transform 1 0 12576 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_127
timestamp 1621261055
transform 1 0 13344 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_135
timestamp 1621261055
transform 1 0 14112 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_143
timestamp 1621261055
transform 1 0 14880 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_964
timestamp 1621261055
transform 1 0 16992 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_151
timestamp 1621261055
transform 1 0 15648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_159
timestamp 1621261055
transform 1 0 16416 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_163
timestamp 1621261055
transform 1 0 16800 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_75_166
timestamp 1621261055
transform 1 0 17088 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _023_
timestamp 1621261055
transform 1 0 17664 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_170
timestamp 1621261055
transform 1 0 17472 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_175
timestamp 1621261055
transform 1 0 17952 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_183
timestamp 1621261055
transform 1 0 18720 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_191
timestamp 1621261055
transform 1 0 19488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_199
timestamp 1621261055
transform 1 0 20256 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_207
timestamp 1621261055
transform 1 0 21024 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_965
timestamp 1621261055
transform 1 0 22272 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_215
timestamp 1621261055
transform 1 0 21792 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_75_219
timestamp 1621261055
transform 1 0 22176 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_221
timestamp 1621261055
transform 1 0 22368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_229
timestamp 1621261055
transform 1 0 23136 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_237
timestamp 1621261055
transform 1 0 23904 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_245
timestamp 1621261055
transform 1 0 24672 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_253
timestamp 1621261055
transform 1 0 25440 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_261
timestamp 1621261055
transform 1 0 26208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_269
timestamp 1621261055
transform 1 0 26976 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_273
timestamp 1621261055
transform 1 0 27360 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_966
timestamp 1621261055
transform 1 0 27552 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_276
timestamp 1621261055
transform 1 0 27648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_284
timestamp 1621261055
transform 1 0 28416 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_292
timestamp 1621261055
transform 1 0 29184 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_300
timestamp 1621261055
transform 1 0 29952 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_308
timestamp 1621261055
transform 1 0 30720 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_967
timestamp 1621261055
transform 1 0 32832 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_316
timestamp 1621261055
transform 1 0 31488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_324
timestamp 1621261055
transform 1 0 32256 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_328
timestamp 1621261055
transform 1 0 32640 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_331
timestamp 1621261055
transform 1 0 32928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_339
timestamp 1621261055
transform 1 0 33696 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_347
timestamp 1621261055
transform 1 0 34464 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_355
timestamp 1621261055
transform 1 0 35232 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_363
timestamp 1621261055
transform 1 0 36000 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_371
timestamp 1621261055
transform 1 0 36768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_968
timestamp 1621261055
transform 1 0 38112 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_379
timestamp 1621261055
transform 1 0 37536 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_383
timestamp 1621261055
transform 1 0 37920 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_386
timestamp 1621261055
transform 1 0 38208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_394
timestamp 1621261055
transform 1 0 38976 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_402
timestamp 1621261055
transform 1 0 39744 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_410
timestamp 1621261055
transform 1 0 40512 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_418
timestamp 1621261055
transform 1 0 41280 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_969
timestamp 1621261055
transform 1 0 43392 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_426
timestamp 1621261055
transform 1 0 42048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_434
timestamp 1621261055
transform 1 0 42816 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_438
timestamp 1621261055
transform 1 0 43200 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_441
timestamp 1621261055
transform 1 0 43488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_449
timestamp 1621261055
transform 1 0 44256 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_457
timestamp 1621261055
transform 1 0 45024 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_465
timestamp 1621261055
transform 1 0 45792 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_473
timestamp 1621261055
transform 1 0 46560 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_481
timestamp 1621261055
transform 1 0 47328 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_970
timestamp 1621261055
transform 1 0 48672 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_489
timestamp 1621261055
transform 1 0 48096 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_493
timestamp 1621261055
transform 1 0 48480 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_496
timestamp 1621261055
transform 1 0 48768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_504
timestamp 1621261055
transform 1 0 49536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_512
timestamp 1621261055
transform 1 0 50304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_520
timestamp 1621261055
transform 1 0 51072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_528
timestamp 1621261055
transform 1 0 51840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_536
timestamp 1621261055
transform 1 0 52608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_544
timestamp 1621261055
transform 1 0 53376 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_971
timestamp 1621261055
transform 1 0 53952 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_548
timestamp 1621261055
transform 1 0 53760 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_551
timestamp 1621261055
transform 1 0 54048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_559
timestamp 1621261055
transform 1 0 54816 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_567
timestamp 1621261055
transform 1 0 55584 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_575
timestamp 1621261055
transform 1 0 56352 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_583
timestamp 1621261055
transform 1 0 57120 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_151
timestamp 1621261055
transform -1 0 58848 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_75_591
timestamp 1621261055
transform 1 0 57888 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_595
timestamp 1621261055
transform 1 0 58272 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _103_
timestamp 1621261055
transform 1 0 2400 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_152
timestamp 1621261055
transform 1 0 1152 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_160
timestamp 1621261055
transform 1 0 2208 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_76_4
timestamp 1621261055
transform 1 0 1536 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_8
timestamp 1621261055
transform 1 0 1920 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_76_10
timestamp 1621261055
transform 1 0 2112 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_16
timestamp 1621261055
transform 1 0 2688 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_972
timestamp 1621261055
transform 1 0 3840 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_24
timestamp 1621261055
transform 1 0 3456 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_76_29
timestamp 1621261055
transform 1 0 3936 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_37
timestamp 1621261055
transform 1 0 4704 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_45
timestamp 1621261055
transform 1 0 5472 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_53
timestamp 1621261055
transform 1 0 6240 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_61
timestamp 1621261055
transform 1 0 7008 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_973
timestamp 1621261055
transform 1 0 9120 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_69
timestamp 1621261055
transform 1 0 7776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_77
timestamp 1621261055
transform 1 0 8544 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_81
timestamp 1621261055
transform 1 0 8928 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_84
timestamp 1621261055
transform 1 0 9216 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_92
timestamp 1621261055
transform 1 0 9984 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_100
timestamp 1621261055
transform 1 0 10752 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_108
timestamp 1621261055
transform 1 0 11520 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_116
timestamp 1621261055
transform 1 0 12288 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_124
timestamp 1621261055
transform 1 0 13056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_974
timestamp 1621261055
transform 1 0 14400 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_132
timestamp 1621261055
transform 1 0 13824 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_136
timestamp 1621261055
transform 1 0 14208 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_139
timestamp 1621261055
transform 1 0 14496 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_147
timestamp 1621261055
transform 1 0 15264 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_155
timestamp 1621261055
transform 1 0 16032 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_163
timestamp 1621261055
transform 1 0 16800 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _129_
timestamp 1621261055
transform 1 0 17760 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_180
timestamp 1621261055
transform 1 0 17568 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_176
timestamp 1621261055
transform 1 0 18048 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_184
timestamp 1621261055
transform 1 0 18816 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_975
timestamp 1621261055
transform 1 0 19680 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_76_192
timestamp 1621261055
transform 1 0 19584 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_194
timestamp 1621261055
transform 1 0 19776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_202
timestamp 1621261055
transform 1 0 20544 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_210
timestamp 1621261055
transform 1 0 21312 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_218
timestamp 1621261055
transform 1 0 22080 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_226
timestamp 1621261055
transform 1 0 22848 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_976
timestamp 1621261055
transform 1 0 24960 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_234
timestamp 1621261055
transform 1 0 23616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_242
timestamp 1621261055
transform 1 0 24384 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_246
timestamp 1621261055
transform 1 0 24768 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_249
timestamp 1621261055
transform 1 0 25056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_257
timestamp 1621261055
transform 1 0 25824 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_265
timestamp 1621261055
transform 1 0 26592 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_273
timestamp 1621261055
transform 1 0 27360 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_281
timestamp 1621261055
transform 1 0 28128 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_289
timestamp 1621261055
transform 1 0 28896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_977
timestamp 1621261055
transform 1 0 30240 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_297
timestamp 1621261055
transform 1 0 29664 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_301
timestamp 1621261055
transform 1 0 30048 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_304
timestamp 1621261055
transform 1 0 30336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_312
timestamp 1621261055
transform 1 0 31104 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _137_
timestamp 1621261055
transform 1 0 32256 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_188
timestamp 1621261055
transform 1 0 32064 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_320
timestamp 1621261055
transform 1 0 31872 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_327
timestamp 1621261055
transform 1 0 32544 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_335
timestamp 1621261055
transform 1 0 33312 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_343
timestamp 1621261055
transform 1 0 34080 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_351
timestamp 1621261055
transform 1 0 34848 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_355
timestamp 1621261055
transform 1 0 35232 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_76_357
timestamp 1621261055
transform 1 0 35424 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_978
timestamp 1621261055
transform 1 0 35520 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_359
timestamp 1621261055
transform 1 0 35616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_367
timestamp 1621261055
transform 1 0 36384 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_375
timestamp 1621261055
transform 1 0 37152 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_218
timestamp 1621261055
transform -1 0 39552 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_383
timestamp 1621261055
transform 1 0 37920 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_391
timestamp 1621261055
transform 1 0 38688 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_395
timestamp 1621261055
transform 1 0 39072 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_76_397
timestamp 1621261055
transform 1 0 39264 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _202_
timestamp 1621261055
transform -1 0 39840 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_979
timestamp 1621261055
transform 1 0 40800 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_403
timestamp 1621261055
transform 1 0 39840 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_411
timestamp 1621261055
transform 1 0 40608 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_414
timestamp 1621261055
transform 1 0 40896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _108_
timestamp 1621261055
transform -1 0 43392 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_170
timestamp 1621261055
transform -1 0 43104 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_422
timestamp 1621261055
transform 1 0 41664 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_430
timestamp 1621261055
transform 1 0 42432 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_76_434
timestamp 1621261055
transform 1 0 42816 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_440
timestamp 1621261055
transform 1 0 43392 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_448
timestamp 1621261055
transform 1 0 44160 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_456
timestamp 1621261055
transform 1 0 44928 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_980
timestamp 1621261055
transform 1 0 46080 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_464
timestamp 1621261055
transform 1 0 45696 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_76_469
timestamp 1621261055
transform 1 0 46176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_477
timestamp 1621261055
transform 1 0 46944 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_485
timestamp 1621261055
transform 1 0 47712 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_493
timestamp 1621261055
transform 1 0 48480 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_501
timestamp 1621261055
transform 1 0 49248 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_981
timestamp 1621261055
transform 1 0 51360 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_509
timestamp 1621261055
transform 1 0 50016 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_517
timestamp 1621261055
transform 1 0 50784 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_521
timestamp 1621261055
transform 1 0 51168 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_524
timestamp 1621261055
transform 1 0 51456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_532
timestamp 1621261055
transform 1 0 52224 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_540
timestamp 1621261055
transform 1 0 52992 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_548
timestamp 1621261055
transform 1 0 53760 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_556
timestamp 1621261055
transform 1 0 54528 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_564
timestamp 1621261055
transform 1 0 55296 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _188_
timestamp 1621261055
transform -1 0 56256 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_982
timestamp 1621261055
transform 1 0 56640 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_84
timestamp 1621261055
transform -1 0 57696 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_234
timestamp 1621261055
transform -1 0 55968 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_76_568
timestamp 1621261055
transform 1 0 55680 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_574
timestamp 1621261055
transform 1 0 56256 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_76_579
timestamp 1621261055
transform 1 0 56736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_153
timestamp 1621261055
transform -1 0 58848 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output436
timestamp 1621261055
transform -1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_76_593
timestamp 1621261055
transform 1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_154
timestamp 1621261055
transform 1 0 1152 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_156
timestamp 1621261055
transform 1 0 1152 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_4
timestamp 1621261055
transform 1 0 1536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_12
timestamp 1621261055
transform 1 0 2304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_20
timestamp 1621261055
transform 1 0 3072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_4
timestamp 1621261055
transform 1 0 1536 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_12
timestamp 1621261055
transform 1 0 2304 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_20
timestamp 1621261055
transform 1 0 3072 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_993
timestamp 1621261055
transform 1 0 3840 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_28
timestamp 1621261055
transform 1 0 3840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_36
timestamp 1621261055
transform 1 0 4608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_29
timestamp 1621261055
transform 1 0 3936 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_37
timestamp 1621261055
transform 1 0 4704 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_983
timestamp 1621261055
transform 1 0 6432 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_44
timestamp 1621261055
transform 1 0 5376 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_52
timestamp 1621261055
transform 1 0 6144 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_77_54
timestamp 1621261055
transform 1 0 6336 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_56
timestamp 1621261055
transform 1 0 6528 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_45
timestamp 1621261055
transform 1 0 5472 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_53
timestamp 1621261055
transform 1 0 6240 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_61
timestamp 1621261055
transform 1 0 7008 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_994
timestamp 1621261055
transform 1 0 9120 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_64
timestamp 1621261055
transform 1 0 7296 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_72
timestamp 1621261055
transform 1 0 8064 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_80
timestamp 1621261055
transform 1 0 8832 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_69
timestamp 1621261055
transform 1 0 7776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_77
timestamp 1621261055
transform 1 0 8544 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_81
timestamp 1621261055
transform 1 0 8928 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_84
timestamp 1621261055
transform 1 0 9216 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_88
timestamp 1621261055
transform 1 0 9600 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_96
timestamp 1621261055
transform 1 0 10368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_104
timestamp 1621261055
transform 1 0 11136 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_92
timestamp 1621261055
transform 1 0 9984 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_100
timestamp 1621261055
transform 1 0 10752 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_984
timestamp 1621261055
transform 1 0 11712 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_108
timestamp 1621261055
transform 1 0 11520 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_111
timestamp 1621261055
transform 1 0 11808 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_119
timestamp 1621261055
transform 1 0 12576 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_108
timestamp 1621261055
transform 1 0 11520 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_116
timestamp 1621261055
transform 1 0 12288 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_124
timestamp 1621261055
transform 1 0 13056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_995
timestamp 1621261055
transform 1 0 14400 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_127
timestamp 1621261055
transform 1 0 13344 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_135
timestamp 1621261055
transform 1 0 14112 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_143
timestamp 1621261055
transform 1 0 14880 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_132
timestamp 1621261055
transform 1 0 13824 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_136
timestamp 1621261055
transform 1 0 14208 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_139
timestamp 1621261055
transform 1 0 14496 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_147
timestamp 1621261055
transform 1 0 15264 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_985
timestamp 1621261055
transform 1 0 16992 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_151
timestamp 1621261055
transform 1 0 15648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_159
timestamp 1621261055
transform 1 0 16416 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_163
timestamp 1621261055
transform 1 0 16800 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_166
timestamp 1621261055
transform 1 0 17088 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_155
timestamp 1621261055
transform 1 0 16032 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_163
timestamp 1621261055
transform 1 0 16800 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_174
timestamp 1621261055
transform 1 0 17856 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_182
timestamp 1621261055
transform 1 0 18624 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_171
timestamp 1621261055
transform 1 0 17568 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_179
timestamp 1621261055
transform 1 0 18336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_187
timestamp 1621261055
transform 1 0 19104 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_996
timestamp 1621261055
transform 1 0 19680 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_190
timestamp 1621261055
transform 1 0 19392 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_198
timestamp 1621261055
transform 1 0 20160 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_206
timestamp 1621261055
transform 1 0 20928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_191
timestamp 1621261055
transform 1 0 19488 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_194
timestamp 1621261055
transform 1 0 19776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_202
timestamp 1621261055
transform 1 0 20544 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_210
timestamp 1621261055
transform 1 0 21312 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_986
timestamp 1621261055
transform 1 0 22272 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_77_214
timestamp 1621261055
transform 1 0 21696 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_218
timestamp 1621261055
transform 1 0 22080 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_221
timestamp 1621261055
transform 1 0 22368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_229
timestamp 1621261055
transform 1 0 23136 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_218
timestamp 1621261055
transform 1 0 22080 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_226
timestamp 1621261055
transform 1 0 22848 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_997
timestamp 1621261055
transform 1 0 24960 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_203
timestamp 1621261055
transform 1 0 25248 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_237
timestamp 1621261055
transform 1 0 23904 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_245
timestamp 1621261055
transform 1 0 24672 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_234
timestamp 1621261055
transform 1 0 23616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_242
timestamp 1621261055
transform 1 0 24384 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_246
timestamp 1621261055
transform 1 0 24768 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_249
timestamp 1621261055
transform 1 0 25056 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_256
timestamp 1621261055
transform 1 0 25728 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_253
timestamp 1621261055
transform 1 0 25440 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _150_
timestamp 1621261055
transform 1 0 25440 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_269
timestamp 1621261055
transform 1 0 26976 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_269
timestamp 1621261055
transform 1 0 26976 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_261
timestamp 1621261055
transform 1 0 26208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_27
timestamp 1621261055
transform 1 0 26496 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _034_
timestamp 1621261055
transform 1 0 26688 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_273
timestamp 1621261055
transform 1 0 27360 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_97
timestamp 1621261055
transform 1 0 27168 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _155_
timestamp 1621261055
transform 1 0 27360 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_987
timestamp 1621261055
transform 1 0 27552 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_276
timestamp 1621261055
transform 1 0 27648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_284
timestamp 1621261055
transform 1 0 28416 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_292
timestamp 1621261055
transform 1 0 29184 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_276
timestamp 1621261055
transform 1 0 27648 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_284
timestamp 1621261055
transform 1 0 28416 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_292
timestamp 1621261055
transform 1 0 29184 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_998
timestamp 1621261055
transform 1 0 30240 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_300
timestamp 1621261055
transform 1 0 29952 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_308
timestamp 1621261055
transform 1 0 30720 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_300
timestamp 1621261055
transform 1 0 29952 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_78_302
timestamp 1621261055
transform 1 0 30144 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_304
timestamp 1621261055
transform 1 0 30336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_312
timestamp 1621261055
transform 1 0 31104 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_988
timestamp 1621261055
transform 1 0 32832 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_316
timestamp 1621261055
transform 1 0 31488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_324
timestamp 1621261055
transform 1 0 32256 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_328
timestamp 1621261055
transform 1 0 32640 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_331
timestamp 1621261055
transform 1 0 32928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_320
timestamp 1621261055
transform 1 0 31872 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_328
timestamp 1621261055
transform 1 0 32640 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_336
timestamp 1621261055
transform 1 0 33408 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_339
timestamp 1621261055
transform 1 0 33696 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_347
timestamp 1621261055
transform 1 0 34464 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_355
timestamp 1621261055
transform 1 0 35232 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_344
timestamp 1621261055
transform 1 0 34176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_352
timestamp 1621261055
transform 1 0 34944 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_356
timestamp 1621261055
transform 1 0 35328 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_999
timestamp 1621261055
transform 1 0 35520 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_363
timestamp 1621261055
transform 1 0 36000 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_371
timestamp 1621261055
transform 1 0 36768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_359
timestamp 1621261055
transform 1 0 35616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_367
timestamp 1621261055
transform 1 0 36384 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_375
timestamp 1621261055
transform 1 0 37152 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_989
timestamp 1621261055
transform 1 0 38112 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_77_379
timestamp 1621261055
transform 1 0 37536 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_383
timestamp 1621261055
transform 1 0 37920 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_386
timestamp 1621261055
transform 1 0 38208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_394
timestamp 1621261055
transform 1 0 38976 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_383
timestamp 1621261055
transform 1 0 37920 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_391
timestamp 1621261055
transform 1 0 38688 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_399
timestamp 1621261055
transform 1 0 39456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1000
timestamp 1621261055
transform 1 0 40800 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_402
timestamp 1621261055
transform 1 0 39744 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_410
timestamp 1621261055
transform 1 0 40512 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_418
timestamp 1621261055
transform 1 0 41280 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_407
timestamp 1621261055
transform 1 0 40224 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_411
timestamp 1621261055
transform 1 0 40608 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_414
timestamp 1621261055
transform 1 0 40896 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_990
timestamp 1621261055
transform 1 0 43392 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_426
timestamp 1621261055
transform 1 0 42048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_434
timestamp 1621261055
transform 1 0 42816 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_438
timestamp 1621261055
transform 1 0 43200 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_441
timestamp 1621261055
transform 1 0 43488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_422
timestamp 1621261055
transform 1 0 41664 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_430
timestamp 1621261055
transform 1 0 42432 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_438
timestamp 1621261055
transform 1 0 43200 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_449
timestamp 1621261055
transform 1 0 44256 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_457
timestamp 1621261055
transform 1 0 45024 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_446
timestamp 1621261055
transform 1 0 43968 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_454
timestamp 1621261055
transform 1 0 44736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_462
timestamp 1621261055
transform 1 0 45504 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1001
timestamp 1621261055
transform 1 0 46080 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_465
timestamp 1621261055
transform 1 0 45792 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_473
timestamp 1621261055
transform 1 0 46560 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_481
timestamp 1621261055
transform 1 0 47328 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_466
timestamp 1621261055
transform 1 0 45888 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_469
timestamp 1621261055
transform 1 0 46176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_477
timestamp 1621261055
transform 1 0 46944 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_991
timestamp 1621261055
transform 1 0 48672 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_77_489
timestamp 1621261055
transform 1 0 48096 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_493
timestamp 1621261055
transform 1 0 48480 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_496
timestamp 1621261055
transform 1 0 48768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_504
timestamp 1621261055
transform 1 0 49536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_485
timestamp 1621261055
transform 1 0 47712 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_493
timestamp 1621261055
transform 1 0 48480 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_501
timestamp 1621261055
transform 1 0 49248 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1002
timestamp 1621261055
transform 1 0 51360 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_512
timestamp 1621261055
transform 1 0 50304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_520
timestamp 1621261055
transform 1 0 51072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_509
timestamp 1621261055
transform 1 0 50016 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_517
timestamp 1621261055
transform 1 0 50784 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_521
timestamp 1621261055
transform 1 0 51168 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_524
timestamp 1621261055
transform 1 0 51456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_528
timestamp 1621261055
transform 1 0 51840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_536
timestamp 1621261055
transform 1 0 52608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_544
timestamp 1621261055
transform 1 0 53376 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_532
timestamp 1621261055
transform 1 0 52224 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_540
timestamp 1621261055
transform 1 0 52992 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_992
timestamp 1621261055
transform 1 0 53952 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_548
timestamp 1621261055
transform 1 0 53760 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_551
timestamp 1621261055
transform 1 0 54048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_559
timestamp 1621261055
transform 1 0 54816 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_567
timestamp 1621261055
transform 1 0 55584 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_548
timestamp 1621261055
transform 1 0 53760 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_556
timestamp 1621261055
transform 1 0 54528 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_564
timestamp 1621261055
transform 1 0 55296 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_576
timestamp 1621261055
transform 1 0 56448 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_572
timestamp 1621261055
transform 1 0 56064 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_224
timestamp 1621261055
transform -1 0 56544 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_579
timestamp 1621261055
transform 1 0 56736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_584
timestamp 1621261055
transform 1 0 57216 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_580
timestamp 1621261055
transform 1 0 56832 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1003
timestamp 1621261055
transform 1 0 56640 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _204_
timestamp 1621261055
transform -1 0 56832 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_77_586
timestamp 1621261055
transform 1 0 57408 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_81
timestamp 1621261055
transform -1 0 57696 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_28
timestamp 1621261055
transform -1 0 57696 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_155
timestamp 1621261055
transform -1 0 58848 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_157
timestamp 1621261055
transform -1 0 58848 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output398
timestamp 1621261055
transform -1 0 58080 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output435
timestamp 1621261055
transform -1 0 58080 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_82
timestamp 1621261055
transform -1 0 58272 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_595
timestamp 1621261055
transform 1 0 58272 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_593
timestamp 1621261055
transform 1 0 58080 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_158
timestamp 1621261055
transform 1 0 1152 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output406
timestamp 1621261055
transform 1 0 1536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_8
timestamp 1621261055
transform 1 0 1920 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_16
timestamp 1621261055
transform 1 0 2688 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output428
timestamp 1621261055
transform 1 0 4320 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_72
timestamp 1621261055
transform 1 0 4128 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_24
timestamp 1621261055
transform 1 0 3456 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_28
timestamp 1621261055
transform 1 0 3840 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_30
timestamp 1621261055
transform 1 0 4032 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_37
timestamp 1621261055
transform 1 0 4704 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1004
timestamp 1621261055
transform 1 0 6432 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_45
timestamp 1621261055
transform 1 0 5472 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_53
timestamp 1621261055
transform 1 0 6240 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_56
timestamp 1621261055
transform 1 0 6528 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output438
timestamp 1621261055
transform 1 0 7488 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output439
timestamp 1621261055
transform -1 0 9504 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_88
timestamp 1621261055
transform 1 0 7296 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_90
timestamp 1621261055
transform -1 0 9120 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_70
timestamp 1621261055
transform 1 0 7872 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_78
timestamp 1621261055
transform 1 0 8640 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_80
timestamp 1621261055
transform 1 0 8832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_87
timestamp 1621261055
transform 1 0 9504 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_95
timestamp 1621261055
transform 1 0 10272 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_103
timestamp 1621261055
transform 1 0 11040 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1005
timestamp 1621261055
transform 1 0 11712 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_107
timestamp 1621261055
transform 1 0 11424 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_109
timestamp 1621261055
transform 1 0 11616 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_111
timestamp 1621261055
transform 1 0 11808 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_119
timestamp 1621261055
transform 1 0 12576 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output442
timestamp 1621261055
transform 1 0 13824 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_92
timestamp 1621261055
transform 1 0 13632 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_127
timestamp 1621261055
transform 1 0 13344 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_129
timestamp 1621261055
transform 1 0 13536 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_136
timestamp 1621261055
transform 1 0 14208 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_144
timestamp 1621261055
transform 1 0 14976 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1006
timestamp 1621261055
transform 1 0 16992 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_152
timestamp 1621261055
transform 1 0 15744 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_160
timestamp 1621261055
transform 1 0 16512 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_164
timestamp 1621261055
transform 1 0 16896 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_166
timestamp 1621261055
transform 1 0 17088 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_174
timestamp 1621261055
transform 1 0 17856 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_182
timestamp 1621261055
transform 1 0 18624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output409
timestamp 1621261055
transform 1 0 20160 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_42
timestamp 1621261055
transform 1 0 19968 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_190
timestamp 1621261055
transform 1 0 19392 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_194
timestamp 1621261055
transform 1 0 19776 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_202
timestamp 1621261055
transform 1 0 20544 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_210
timestamp 1621261055
transform 1 0 21312 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1007
timestamp 1621261055
transform 1 0 22272 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output411
timestamp 1621261055
transform -1 0 23712 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_44
timestamp 1621261055
transform -1 0 23328 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_218
timestamp 1621261055
transform 1 0 22080 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_221
timestamp 1621261055
transform 1 0 22368 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output412
timestamp 1621261055
transform 1 0 24864 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_46
timestamp 1621261055
transform 1 0 24672 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_235
timestamp 1621261055
transform 1 0 23712 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_243
timestamp 1621261055
transform 1 0 24480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_251
timestamp 1621261055
transform 1 0 25248 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_259
timestamp 1621261055
transform 1 0 26016 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_267
timestamp 1621261055
transform 1 0 26784 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _073_
timestamp 1621261055
transform -1 0 29280 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _169_
timestamp 1621261055
transform 1 0 28032 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1008
timestamp 1621261055
transform 1 0 27552 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_115
timestamp 1621261055
transform 1 0 27840 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_134
timestamp 1621261055
transform -1 0 28992 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_276
timestamp 1621261055
transform 1 0 27648 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_283
timestamp 1621261055
transform 1 0 28320 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_287
timestamp 1621261055
transform 1 0 28704 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_293
timestamp 1621261055
transform 1 0 29280 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_301
timestamp 1621261055
transform 1 0 30048 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_309
timestamp 1621261055
transform 1 0 30816 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1009
timestamp 1621261055
transform 1 0 32832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_317
timestamp 1621261055
transform 1 0 31584 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_325
timestamp 1621261055
transform 1 0 32352 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_329
timestamp 1621261055
transform 1 0 32736 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_331
timestamp 1621261055
transform 1 0 32928 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_339
timestamp 1621261055
transform 1 0 33696 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_347
timestamp 1621261055
transform 1 0 34464 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_355
timestamp 1621261055
transform 1 0 35232 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_363
timestamp 1621261055
transform 1 0 36000 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_371
timestamp 1621261055
transform 1 0 36768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1010
timestamp 1621261055
transform 1 0 38112 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output422
timestamp 1621261055
transform -1 0 39456 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_66
timestamp 1621261055
transform -1 0 39072 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_379
timestamp 1621261055
transform 1 0 37536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_383
timestamp 1621261055
transform 1 0 37920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_386
timestamp 1621261055
transform 1 0 38208 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_390
timestamp 1621261055
transform 1 0 38592 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_392
timestamp 1621261055
transform 1 0 38784 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_399
timestamp 1621261055
transform 1 0 39456 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output423
timestamp 1621261055
transform -1 0 41088 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_67
timestamp 1621261055
transform -1 0 40704 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_407
timestamp 1621261055
transform 1 0 40224 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_409
timestamp 1621261055
transform 1 0 40416 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_416
timestamp 1621261055
transform 1 0 41088 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1011
timestamp 1621261055
transform 1 0 43392 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_424
timestamp 1621261055
transform 1 0 41856 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_432
timestamp 1621261055
transform 1 0 42624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_441
timestamp 1621261055
transform 1 0 43488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output426
timestamp 1621261055
transform -1 0 45792 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_70
timestamp 1621261055
transform -1 0 45408 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_449
timestamp 1621261055
transform 1 0 44256 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_457
timestamp 1621261055
transform 1 0 45024 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output427
timestamp 1621261055
transform 1 0 46944 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_465
timestamp 1621261055
transform 1 0 45792 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_473
timestamp 1621261055
transform 1 0 46560 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_481
timestamp 1621261055
transform 1 0 47328 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _127_
timestamp 1621261055
transform -1 0 49440 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1012
timestamp 1621261055
transform 1 0 48672 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_178
timestamp 1621261055
transform -1 0 49152 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_489
timestamp 1621261055
transform 1 0 48096 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_493
timestamp 1621261055
transform 1 0 48480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_496
timestamp 1621261055
transform 1 0 48768 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_503
timestamp 1621261055
transform 1 0 49440 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_511
timestamp 1621261055
transform 1 0 50208 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_519
timestamp 1621261055
transform 1 0 50976 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output431
timestamp 1621261055
transform 1 0 51744 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_531
timestamp 1621261055
transform 1 0 52128 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_539
timestamp 1621261055
transform 1 0 52896 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1013
timestamp 1621261055
transform 1 0 53952 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_547
timestamp 1621261055
transform 1 0 53664 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_549
timestamp 1621261055
transform 1 0 53856 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_551
timestamp 1621261055
transform 1 0 54048 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_559
timestamp 1621261055
transform 1 0 54816 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_567
timestamp 1621261055
transform 1 0 55584 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output397
timestamp 1621261055
transform -1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output434
timestamp 1621261055
transform -1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_26
timestamp 1621261055
transform -1 0 57504 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_79
timestamp 1621261055
transform -1 0 56448 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_571
timestamp 1621261055
transform 1 0 55968 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_573
timestamp 1621261055
transform 1 0 56160 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_79_580
timestamp 1621261055
transform 1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_584
timestamp 1621261055
transform 1 0 57216 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_159
timestamp 1621261055
transform -1 0 58848 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_79_591
timestamp 1621261055
transform 1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_595
timestamp 1621261055
transform 1 0 58272 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_160
timestamp 1621261055
transform 1 0 1152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output368
timestamp 1621261055
transform 1 0 1536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output379
timestamp 1621261055
transform 1 0 2304 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output417
timestamp 1621261055
transform 1 0 3072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_1
timestamp 1621261055
transform 1 0 1920 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_56
timestamp 1621261055
transform 1 0 2880 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_10
timestamp 1621261055
transform 1 0 2112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_16
timestamp 1621261055
transform 1 0 2688 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1014
timestamp 1621261055
transform 1 0 3840 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output390
timestamp 1621261055
transform 1 0 4320 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_17
timestamp 1621261055
transform 1 0 4128 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_30
timestamp 1621261055
transform 1 0 5184 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_24
timestamp 1621261055
transform 1 0 3456 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_29
timestamp 1621261055
transform 1 0 3936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_37
timestamp 1621261055
transform 1 0 4704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_41
timestamp 1621261055
transform 1 0 5088 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output399
timestamp 1621261055
transform 1 0 5376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output400
timestamp 1621261055
transform 1 0 7008 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output437
timestamp 1621261055
transform 1 0 6144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_32
timestamp 1621261055
transform 1 0 6816 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_86
timestamp 1621261055
transform 1 0 5952 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_48
timestamp 1621261055
transform 1 0 5760 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_56
timestamp 1621261055
transform 1 0 6528 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_58
timestamp 1621261055
transform 1 0 6720 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1015
timestamp 1621261055
transform 1 0 9120 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output401
timestamp 1621261055
transform 1 0 8352 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_65
timestamp 1621261055
transform 1 0 7392 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_73
timestamp 1621261055
transform 1 0 8160 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_79
timestamp 1621261055
transform 1 0 8736 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_84
timestamp 1621261055
transform 1 0 9216 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output402
timestamp 1621261055
transform 1 0 10176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output440
timestamp 1621261055
transform 1 0 10944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_34
timestamp 1621261055
transform 1 0 9984 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_98
timestamp 1621261055
transform 1 0 10560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output403
timestamp 1621261055
transform 1 0 11712 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output441
timestamp 1621261055
transform 1 0 12480 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_36
timestamp 1621261055
transform 1 0 11520 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_106
timestamp 1621261055
transform 1 0 11328 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_114
timestamp 1621261055
transform 1 0 12096 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_122
timestamp 1621261055
transform 1 0 12864 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_126
timestamp 1621261055
transform 1 0 13248 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1016
timestamp 1621261055
transform 1 0 14400 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output404
timestamp 1621261055
transform 1 0 13344 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output405
timestamp 1621261055
transform -1 0 15264 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_38
timestamp 1621261055
transform -1 0 14880 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_131
timestamp 1621261055
transform 1 0 13728 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_135
timestamp 1621261055
transform 1 0 14112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_137
timestamp 1621261055
transform 1 0 14304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_139
timestamp 1621261055
transform 1 0 14496 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_147
timestamp 1621261055
transform 1 0 15264 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output407
timestamp 1621261055
transform -1 0 17376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output443
timestamp 1621261055
transform -1 0 16032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_40
timestamp 1621261055
transform -1 0 16992 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_94
timestamp 1621261055
transform -1 0 15648 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_155
timestamp 1621261055
transform 1 0 16032 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output370
timestamp 1621261055
transform 1 0 18048 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output408
timestamp 1621261055
transform 1 0 18816 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_169
timestamp 1621261055
transform 1 0 17376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_173
timestamp 1621261055
transform 1 0 17760 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_175
timestamp 1621261055
transform 1 0 17952 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_180
timestamp 1621261055
transform 1 0 18432 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_188
timestamp 1621261055
transform 1 0 19200 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1017
timestamp 1621261055
transform 1 0 19680 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output371
timestamp 1621261055
transform 1 0 20160 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output372
timestamp 1621261055
transform -1 0 21600 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_3
timestamp 1621261055
transform -1 0 21216 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_192
timestamp 1621261055
transform 1 0 19584 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_194
timestamp 1621261055
transform 1 0 19776 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_202
timestamp 1621261055
transform 1 0 20544 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_206
timestamp 1621261055
transform 1 0 20928 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output373
timestamp 1621261055
transform -1 0 23136 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output410
timestamp 1621261055
transform 1 0 21984 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_5
timestamp 1621261055
transform -1 0 22752 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_213
timestamp 1621261055
transform 1 0 21600 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_221
timestamp 1621261055
transform 1 0 22368 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_229
timestamp 1621261055
transform 1 0 23136 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1018
timestamp 1621261055
transform 1 0 24960 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output374
timestamp 1621261055
transform -1 0 24576 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_7
timestamp 1621261055
transform -1 0 24192 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_237
timestamp 1621261055
transform 1 0 23904 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_244
timestamp 1621261055
transform 1 0 24576 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_249
timestamp 1621261055
transform 1 0 25056 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output375
timestamp 1621261055
transform 1 0 25920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output413
timestamp 1621261055
transform -1 0 27072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_9
timestamp 1621261055
transform -1 0 27552 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_48
timestamp 1621261055
transform -1 0 26688 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_257
timestamp 1621261055
transform 1 0 25824 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_262
timestamp 1621261055
transform 1 0 26304 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_270
timestamp 1621261055
transform 1 0 27072 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_272
timestamp 1621261055
transform 1 0 27264 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output376
timestamp 1621261055
transform -1 0 27936 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output414
timestamp 1621261055
transform 1 0 28320 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_50
timestamp 1621261055
transform 1 0 28128 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_52
timestamp 1621261055
transform -1 0 29472 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_279
timestamp 1621261055
transform 1 0 27936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_287
timestamp 1621261055
transform 1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_291
timestamp 1621261055
transform 1 0 29088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1019
timestamp 1621261055
transform 1 0 30240 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output378
timestamp 1621261055
transform 1 0 30720 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output415
timestamp 1621261055
transform -1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_54
timestamp 1621261055
transform 1 0 31296 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_299
timestamp 1621261055
transform 1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_304
timestamp 1621261055
transform 1 0 30336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_312
timestamp 1621261055
transform 1 0 31104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output380
timestamp 1621261055
transform 1 0 32256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output416
timestamp 1621261055
transform 1 0 31488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output418
timestamp 1621261055
transform -1 0 33408 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_58
timestamp 1621261055
transform -1 0 33024 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_320
timestamp 1621261055
transform 1 0 31872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_328
timestamp 1621261055
transform 1 0 32640 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_336
timestamp 1621261055
transform 1 0 33408 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output381
timestamp 1621261055
transform 1 0 33792 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output419
timestamp 1621261055
transform -1 0 34944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_60
timestamp 1621261055
transform -1 0 34560 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_344
timestamp 1621261055
transform 1 0 34176 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_352
timestamp 1621261055
transform 1 0 34944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_356
timestamp 1621261055
transform 1 0 35328 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1020
timestamp 1621261055
transform 1 0 35520 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output382
timestamp 1621261055
transform 1 0 36000 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output420
timestamp 1621261055
transform -1 0 37152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_11
timestamp 1621261055
transform 1 0 35808 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_62
timestamp 1621261055
transform -1 0 36768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_64
timestamp 1621261055
transform -1 0 37536 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_359
timestamp 1621261055
transform 1 0 35616 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_367
timestamp 1621261055
transform 1 0 36384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_375
timestamp 1621261055
transform 1 0 37152 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output384
timestamp 1621261055
transform 1 0 38592 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output421
timestamp 1621261055
transform -1 0 37920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_383
timestamp 1621261055
transform 1 0 37920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_387
timestamp 1621261055
transform 1 0 38304 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_389
timestamp 1621261055
transform 1 0 38496 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_394
timestamp 1621261055
transform 1 0 38976 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1021
timestamp 1621261055
transform 1 0 40800 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output385
timestamp 1621261055
transform 1 0 40032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_15
timestamp 1621261055
transform 1 0 39840 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_402
timestamp 1621261055
transform 1 0 39744 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_409
timestamp 1621261055
transform 1 0 40416 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_414
timestamp 1621261055
transform 1 0 40896 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output386
timestamp 1621261055
transform 1 0 41760 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output387
timestamp 1621261055
transform 1 0 43296 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output424
timestamp 1621261055
transform -1 0 42912 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_69
timestamp 1621261055
transform -1 0 42528 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_422
timestamp 1621261055
transform 1 0 41664 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_427
timestamp 1621261055
transform 1 0 42144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_435
timestamp 1621261055
transform 1 0 42912 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output388
timestamp 1621261055
transform 1 0 44928 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output425
timestamp 1621261055
transform 1 0 44064 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_443
timestamp 1621261055
transform 1 0 43680 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_451
timestamp 1621261055
transform 1 0 44448 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_455
timestamp 1621261055
transform 1 0 44832 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_460
timestamp 1621261055
transform 1 0 45312 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1022
timestamp 1621261055
transform 1 0 46080 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output389
timestamp 1621261055
transform 1 0 46560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_469
timestamp 1621261055
transform 1 0 46176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_477
timestamp 1621261055
transform 1 0 46944 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output391
timestamp 1621261055
transform 1 0 48000 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output429
timestamp 1621261055
transform -1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_19
timestamp 1621261055
transform 1 0 49440 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_74
timestamp 1621261055
transform -1 0 48768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_485
timestamp 1621261055
transform 1 0 47712 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_487
timestamp 1621261055
transform 1 0 47904 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_492
timestamp 1621261055
transform 1 0 48384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_500
timestamp 1621261055
transform 1 0 49152 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_502
timestamp 1621261055
transform 1 0 49344 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1023
timestamp 1621261055
transform 1 0 51360 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output392
timestamp 1621261055
transform 1 0 49632 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output430
timestamp 1621261055
transform 1 0 50400 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_76
timestamp 1621261055
transform 1 0 50208 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_509
timestamp 1621261055
transform 1 0 50016 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_517
timestamp 1621261055
transform 1 0 50784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_521
timestamp 1621261055
transform 1 0 51168 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_524
timestamp 1621261055
transform 1 0 51456 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output393
timestamp 1621261055
transform 1 0 51840 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output394
timestamp 1621261055
transform -1 0 53184 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output432
timestamp 1621261055
transform -1 0 53952 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_21
timestamp 1621261055
transform -1 0 52800 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_22
timestamp 1621261055
transform -1 0 53376 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_78
timestamp 1621261055
transform -1 0 53568 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_532
timestamp 1621261055
transform 1 0 52224 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output395
timestamp 1621261055
transform 1 0 54336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output433
timestamp 1621261055
transform 1 0 55104 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_550
timestamp 1621261055
transform 1 0 53952 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_558
timestamp 1621261055
transform 1 0 54720 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_566
timestamp 1621261055
transform 1 0 55488 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1024
timestamp 1621261055
transform 1 0 56640 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output396
timestamp 1621261055
transform -1 0 56256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_24
timestamp 1621261055
transform -1 0 55872 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_574
timestamp 1621261055
transform 1 0 56256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_579
timestamp 1621261055
transform 1 0 56736 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_587
timestamp 1621261055
transform 1 0 57504 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_161
timestamp 1621261055
transform -1 0 58848 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input31
timestamp 1621261055
transform 1 0 57696 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_593
timestamp 1621261055
transform 1 0 58080 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_162
timestamp 1621261055
transform 1 0 1152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input12
timestamp 1621261055
transform 1 0 2400 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_9
timestamp 1621261055
transform 1 0 2016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_18
timestamp 1621261055
transform 1 0 2880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1025
timestamp 1621261055
transform 1 0 3840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input32
timestamp 1621261055
transform 1 0 4896 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_26
timestamp 1621261055
transform 1 0 3648 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_29
timestamp 1621261055
transform 1 0 3936 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_37
timestamp 1621261055
transform 1 0 4704 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1026
timestamp 1621261055
transform 1 0 6528 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input23
timestamp 1621261055
transform 1 0 5760 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input33
timestamp 1621261055
transform 1 0 7008 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_44
timestamp 1621261055
transform 1 0 5376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_52
timestamp 1621261055
transform 1 0 6144 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_57
timestamp 1621261055
transform 1 0 6624 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1027
timestamp 1621261055
transform 1 0 9216 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input34
timestamp 1621261055
transform 1 0 8064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_66
timestamp 1621261055
transform 1 0 7488 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_70
timestamp 1621261055
transform 1 0 7872 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_76
timestamp 1621261055
transform 1 0 8448 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  input35
timestamp 1621261055
transform 1 0 9696 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input36
timestamp 1621261055
transform 1 0 11040 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_85
timestamp 1621261055
transform 1 0 9312 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_93
timestamp 1621261055
transform 1 0 10080 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_101
timestamp 1621261055
transform 1 0 10848 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1028
timestamp 1621261055
transform 1 0 11904 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input37
timestamp 1621261055
transform 1 0 12768 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_108
timestamp 1621261055
transform 1 0 11520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_113
timestamp 1621261055
transform 1 0 12000 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_126
timestamp 1621261055
transform 1 0 13248 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1029
timestamp 1621261055
transform 1 0 14592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input38
timestamp 1621261055
transform 1 0 15072 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output369
timestamp 1621261055
transform 1 0 13824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_130
timestamp 1621261055
transform 1 0 13632 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_136
timestamp 1621261055
transform 1 0 14208 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_141
timestamp 1621261055
transform 1 0 14688 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1030
timestamp 1621261055
transform 1 0 17280 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input2
timestamp 1621261055
transform 1 0 15936 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_149
timestamp 1621261055
transform 1 0 15456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_153
timestamp 1621261055
transform 1 0 15840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_159
timestamp 1621261055
transform 1 0 16416 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_167
timestamp 1621261055
transform 1 0 17184 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input3
timestamp 1621261055
transform 1 0 17760 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input4
timestamp 1621261055
transform 1 0 19104 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_169
timestamp 1621261055
transform 1 0 17376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_178
timestamp 1621261055
transform 1 0 18240 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_186
timestamp 1621261055
transform 1 0 19008 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1031
timestamp 1621261055
transform 1 0 19968 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input5
timestamp 1621261055
transform 1 0 20640 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_192
timestamp 1621261055
transform 1 0 19584 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_197
timestamp 1621261055
transform 1 0 20064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_201
timestamp 1621261055
transform 1 0 20448 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_208
timestamp 1621261055
transform 1 0 21120 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1032
timestamp 1621261055
transform 1 0 22656 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input6
timestamp 1621261055
transform 1 0 21888 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_220
timestamp 1621261055
transform 1 0 22272 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_225
timestamp 1621261055
transform 1 0 22752 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1033
timestamp 1621261055
transform 1 0 25344 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input7
timestamp 1621261055
transform 1 0 23808 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_233
timestamp 1621261055
transform 1 0 23520 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_235
timestamp 1621261055
transform 1 0 23712 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_241
timestamp 1621261055
transform 1 0 24288 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_249
timestamp 1621261055
transform 1 0 25056 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_251
timestamp 1621261055
transform 1 0 25248 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input8
timestamp 1621261055
transform 1 0 25824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input9
timestamp 1621261055
transform 1 0 26976 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_253
timestamp 1621261055
transform 1 0 25440 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_261
timestamp 1621261055
transform 1 0 26208 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1034
timestamp 1621261055
transform 1 0 28032 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input10
timestamp 1621261055
transform 1 0 28608 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_274
timestamp 1621261055
transform 1 0 27456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_278
timestamp 1621261055
transform 1 0 27840 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_281
timestamp 1621261055
transform 1 0 28128 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_285
timestamp 1621261055
transform 1 0 28512 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_290
timestamp 1621261055
transform 1 0 28992 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1035
timestamp 1621261055
transform 1 0 30720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input11
timestamp 1621261055
transform 1 0 29856 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_1  FILLER_81_298
timestamp 1621261055
transform 1 0 29760 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_304
timestamp 1621261055
transform 1 0 30336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_309
timestamp 1621261055
transform 1 0 30816 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1036
timestamp 1621261055
transform 1 0 33408 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input13
timestamp 1621261055
transform 1 0 31680 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output377
timestamp 1621261055
transform 1 0 32448 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_317
timestamp 1621261055
transform 1 0 31584 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_322
timestamp 1621261055
transform 1 0 32064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_330
timestamp 1621261055
transform 1 0 32832 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_334
timestamp 1621261055
transform 1 0 33216 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__buf_2  input14
timestamp 1621261055
transform 1 0 33888 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input15
timestamp 1621261055
transform 1 0 34848 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_337
timestamp 1621261055
transform 1 0 33504 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_346
timestamp 1621261055
transform 1 0 34368 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_350
timestamp 1621261055
transform 1 0 34752 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_355
timestamp 1621261055
transform 1 0 35232 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1037
timestamp 1621261055
transform 1 0 36096 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input16 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 36576 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__fill_1  FILLER_81_363
timestamp 1621261055
transform 1 0 36000 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_365
timestamp 1621261055
transform 1 0 36192 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_375
timestamp 1621261055
transform 1 0 37152 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1038
timestamp 1621261055
transform 1 0 38784 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input17
timestamp 1621261055
transform 1 0 38016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_383
timestamp 1621261055
transform 1 0 37920 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_388
timestamp 1621261055
transform 1 0 38400 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_393
timestamp 1621261055
transform 1 0 38880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1039
timestamp 1621261055
transform 1 0 41472 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input18
timestamp 1621261055
transform 1 0 39648 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_2  output383
timestamp 1621261055
transform -1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_13
timestamp 1621261055
transform -1 0 40608 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_407
timestamp 1621261055
transform 1 0 40224 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_415
timestamp 1621261055
transform 1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_419
timestamp 1621261055
transform 1 0 41376 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input19
timestamp 1621261055
transform 1 0 41952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_4  input20
timestamp 1621261055
transform 1 0 42816 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_421
timestamp 1621261055
transform 1 0 41568 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_429
timestamp 1621261055
transform 1 0 42336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_433
timestamp 1621261055
transform 1 0 42720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_440
timestamp 1621261055
transform 1 0 43392 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1040
timestamp 1621261055
transform 1 0 44160 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input21
timestamp 1621261055
transform 1 0 44640 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_449
timestamp 1621261055
transform 1 0 44256 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_459
timestamp 1621261055
transform 1 0 45216 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1041
timestamp 1621261055
transform 1 0 46848 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input22
timestamp 1621261055
transform 1 0 45888 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input24
timestamp 1621261055
transform 1 0 47520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_463
timestamp 1621261055
transform 1 0 45600 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_465
timestamp 1621261055
transform 1 0 45792 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_472
timestamp 1621261055
transform 1 0 46464 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_477
timestamp 1621261055
transform 1 0 46944 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_481
timestamp 1621261055
transform 1 0 47328 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1042
timestamp 1621261055
transform 1 0 49536 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input25
timestamp 1621261055
transform 1 0 48576 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_487
timestamp 1621261055
transform 1 0 47904 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_491
timestamp 1621261055
transform 1 0 48288 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_493
timestamp 1621261055
transform 1 0 48480 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_500
timestamp 1621261055
transform 1 0 49152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_4  input26
timestamp 1621261055
transform 1 0 50688 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_8  FILLER_81_505
timestamp 1621261055
transform 1 0 49632 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_513
timestamp 1621261055
transform 1 0 50400 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_515
timestamp 1621261055
transform 1 0 50592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_522
timestamp 1621261055
transform 1 0 51264 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1043
timestamp 1621261055
transform 1 0 52224 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input27
timestamp 1621261055
transform 1 0 52704 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_530
timestamp 1621261055
transform 1 0 52032 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_533
timestamp 1621261055
transform 1 0 52320 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_541
timestamp 1621261055
transform 1 0 53088 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1044
timestamp 1621261055
transform 1 0 54912 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input28
timestamp 1621261055
transform 1 0 53856 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_4  input29
timestamp 1621261055
transform 1 0 55392 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_555
timestamp 1621261055
transform 1 0 54432 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_559
timestamp 1621261055
transform 1 0 54816 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_561
timestamp 1621261055
transform 1 0 55008 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1045
timestamp 1621261055
transform 1 0 57600 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input30
timestamp 1621261055
transform 1 0 56640 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_571
timestamp 1621261055
transform 1 0 55968 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_575
timestamp 1621261055
transform 1 0 56352 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_577
timestamp 1621261055
transform 1 0 56544 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_584
timestamp 1621261055
transform 1 0 57216 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_163
timestamp 1621261055
transform -1 0 58848 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_589
timestamp 1621261055
transform 1 0 57696 0 1 56610
box -38 -49 806 715
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 12980 0 13036 800 6 la_data_in[0]
port 114 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_data_in[100]
port 115 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_data_in[101]
port 116 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[102]
port 117 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[103]
port 118 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[104]
port 119 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_data_in[105]
port 120 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_data_in[106]
port 121 nsew signal input
rlabel metal2 s 52244 0 52300 800 6 la_data_in[107]
port 122 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[108]
port 123 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[109]
port 124 nsew signal input
rlabel metal2 s 16628 0 16684 800 6 la_data_in[10]
port 125 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[110]
port 126 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_data_in[111]
port 127 nsew signal input
rlabel metal2 s 54068 0 54124 800 6 la_data_in[112]
port 128 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[113]
port 129 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[114]
port 130 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[115]
port 131 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[116]
port 132 nsew signal input
rlabel metal2 s 55892 0 55948 800 6 la_data_in[117]
port 133 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[118]
port 134 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[119]
port 135 nsew signal input
rlabel metal2 s 17012 0 17068 800 6 la_data_in[11]
port 136 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[120]
port 137 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[121]
port 138 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[122]
port 139 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[123]
port 140 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[124]
port 141 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[125]
port 142 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[126]
port 143 nsew signal input
rlabel metal2 s 59636 0 59692 800 6 la_data_in[127]
port 144 nsew signal input
rlabel metal2 s 17396 0 17452 800 6 la_data_in[12]
port 145 nsew signal input
rlabel metal2 s 17684 0 17740 800 6 la_data_in[13]
port 146 nsew signal input
rlabel metal2 s 18068 0 18124 800 6 la_data_in[14]
port 147 nsew signal input
rlabel metal2 s 18452 0 18508 800 6 la_data_in[15]
port 148 nsew signal input
rlabel metal2 s 18836 0 18892 800 6 la_data_in[16]
port 149 nsew signal input
rlabel metal2 s 19220 0 19276 800 6 la_data_in[17]
port 150 nsew signal input
rlabel metal2 s 19604 0 19660 800 6 la_data_in[18]
port 151 nsew signal input
rlabel metal2 s 19892 0 19948 800 6 la_data_in[19]
port 152 nsew signal input
rlabel metal2 s 13364 0 13420 800 6 la_data_in[1]
port 153 nsew signal input
rlabel metal2 s 20276 0 20332 800 6 la_data_in[20]
port 154 nsew signal input
rlabel metal2 s 20660 0 20716 800 6 la_data_in[21]
port 155 nsew signal input
rlabel metal2 s 21044 0 21100 800 6 la_data_in[22]
port 156 nsew signal input
rlabel metal2 s 21428 0 21484 800 6 la_data_in[23]
port 157 nsew signal input
rlabel metal2 s 21812 0 21868 800 6 la_data_in[24]
port 158 nsew signal input
rlabel metal2 s 22100 0 22156 800 6 la_data_in[25]
port 159 nsew signal input
rlabel metal2 s 22484 0 22540 800 6 la_data_in[26]
port 160 nsew signal input
rlabel metal2 s 22868 0 22924 800 6 la_data_in[27]
port 161 nsew signal input
rlabel metal2 s 23252 0 23308 800 6 la_data_in[28]
port 162 nsew signal input
rlabel metal2 s 23636 0 23692 800 6 la_data_in[29]
port 163 nsew signal input
rlabel metal2 s 13652 0 13708 800 6 la_data_in[2]
port 164 nsew signal input
rlabel metal2 s 24020 0 24076 800 6 la_data_in[30]
port 165 nsew signal input
rlabel metal2 s 24308 0 24364 800 6 la_data_in[31]
port 166 nsew signal input
rlabel metal2 s 24692 0 24748 800 6 la_data_in[32]
port 167 nsew signal input
rlabel metal2 s 25076 0 25132 800 6 la_data_in[33]
port 168 nsew signal input
rlabel metal2 s 25460 0 25516 800 6 la_data_in[34]
port 169 nsew signal input
rlabel metal2 s 25844 0 25900 800 6 la_data_in[35]
port 170 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_in[36]
port 171 nsew signal input
rlabel metal2 s 26516 0 26572 800 6 la_data_in[37]
port 172 nsew signal input
rlabel metal2 s 26900 0 26956 800 6 la_data_in[38]
port 173 nsew signal input
rlabel metal2 s 27284 0 27340 800 6 la_data_in[39]
port 174 nsew signal input
rlabel metal2 s 14036 0 14092 800 6 la_data_in[3]
port 175 nsew signal input
rlabel metal2 s 27668 0 27724 800 6 la_data_in[40]
port 176 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_data_in[41]
port 177 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 la_data_in[42]
port 178 nsew signal input
rlabel metal2 s 28724 0 28780 800 6 la_data_in[43]
port 179 nsew signal input
rlabel metal2 s 29108 0 29164 800 6 la_data_in[44]
port 180 nsew signal input
rlabel metal2 s 29492 0 29548 800 6 la_data_in[45]
port 181 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_data_in[46]
port 182 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_data_in[47]
port 183 nsew signal input
rlabel metal2 s 30548 0 30604 800 6 la_data_in[48]
port 184 nsew signal input
rlabel metal2 s 30932 0 30988 800 6 la_data_in[49]
port 185 nsew signal input
rlabel metal2 s 14420 0 14476 800 6 la_data_in[4]
port 186 nsew signal input
rlabel metal2 s 31316 0 31372 800 6 la_data_in[50]
port 187 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_data_in[51]
port 188 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_data_in[52]
port 189 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_data_in[53]
port 190 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 la_data_in[54]
port 191 nsew signal input
rlabel metal2 s 33140 0 33196 800 6 la_data_in[55]
port 192 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_data_in[56]
port 193 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_data_in[57]
port 194 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_data_in[58]
port 195 nsew signal input
rlabel metal2 s 34580 0 34636 800 6 la_data_in[59]
port 196 nsew signal input
rlabel metal2 s 14804 0 14860 800 6 la_data_in[5]
port 197 nsew signal input
rlabel metal2 s 34964 0 35020 800 6 la_data_in[60]
port 198 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_data_in[61]
port 199 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_data_in[62]
port 200 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_data_in[63]
port 201 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_data_in[64]
port 202 nsew signal input
rlabel metal2 s 36788 0 36844 800 6 la_data_in[65]
port 203 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_data_in[66]
port 204 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_data_in[67]
port 205 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_data_in[68]
port 206 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_data_in[69]
port 207 nsew signal input
rlabel metal2 s 15188 0 15244 800 6 la_data_in[6]
port 208 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_data_in[70]
port 209 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_data_in[71]
port 210 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_data_in[72]
port 211 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_data_in[73]
port 212 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_data_in[74]
port 213 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_data_in[75]
port 214 nsew signal input
rlabel metal2 s 40916 0 40972 800 6 la_data_in[76]
port 215 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_data_in[77]
port 216 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_data_in[78]
port 217 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_data_in[79]
port 218 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 219 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_data_in[80]
port 220 nsew signal input
rlabel metal2 s 42740 0 42796 800 6 la_data_in[81]
port 221 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_data_in[82]
port 222 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_data_in[83]
port 223 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_data_in[84]
port 224 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_data_in[85]
port 225 nsew signal input
rlabel metal2 s 44564 0 44620 800 6 la_data_in[86]
port 226 nsew signal input
rlabel metal2 s 44948 0 45004 800 6 la_data_in[87]
port 227 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_data_in[88]
port 228 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_data_in[89]
port 229 nsew signal input
rlabel metal2 s 15860 0 15916 800 6 la_data_in[8]
port 230 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_data_in[90]
port 231 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_data_in[91]
port 232 nsew signal input
rlabel metal2 s 46772 0 46828 800 6 la_data_in[92]
port 233 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[93]
port 234 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_data_in[94]
port 235 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_data_in[95]
port 236 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_data_in[96]
port 237 nsew signal input
rlabel metal2 s 48596 0 48652 800 6 la_data_in[97]
port 238 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[98]
port 239 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[99]
port 240 nsew signal input
rlabel metal2 s 16244 0 16300 800 6 la_data_in[9]
port 241 nsew signal input
rlabel metal2 s 13076 0 13132 800 6 la_data_out[0]
port 242 nsew signal tristate
rlabel metal2 s 49844 0 49900 800 6 la_data_out[100]
port 243 nsew signal tristate
rlabel metal2 s 50132 0 50188 800 6 la_data_out[101]
port 244 nsew signal tristate
rlabel metal2 s 50516 0 50572 800 6 la_data_out[102]
port 245 nsew signal tristate
rlabel metal2 s 50900 0 50956 800 6 la_data_out[103]
port 246 nsew signal tristate
rlabel metal2 s 51284 0 51340 800 6 la_data_out[104]
port 247 nsew signal tristate
rlabel metal2 s 51668 0 51724 800 6 la_data_out[105]
port 248 nsew signal tristate
rlabel metal2 s 52052 0 52108 800 6 la_data_out[106]
port 249 nsew signal tristate
rlabel metal2 s 52340 0 52396 800 6 la_data_out[107]
port 250 nsew signal tristate
rlabel metal2 s 52724 0 52780 800 6 la_data_out[108]
port 251 nsew signal tristate
rlabel metal2 s 53108 0 53164 800 6 la_data_out[109]
port 252 nsew signal tristate
rlabel metal2 s 16724 0 16780 800 6 la_data_out[10]
port 253 nsew signal tristate
rlabel metal2 s 53492 0 53548 800 6 la_data_out[110]
port 254 nsew signal tristate
rlabel metal2 s 53876 0 53932 800 6 la_data_out[111]
port 255 nsew signal tristate
rlabel metal2 s 54260 0 54316 800 6 la_data_out[112]
port 256 nsew signal tristate
rlabel metal2 s 54548 0 54604 800 6 la_data_out[113]
port 257 nsew signal tristate
rlabel metal2 s 54932 0 54988 800 6 la_data_out[114]
port 258 nsew signal tristate
rlabel metal2 s 55316 0 55372 800 6 la_data_out[115]
port 259 nsew signal tristate
rlabel metal2 s 55700 0 55756 800 6 la_data_out[116]
port 260 nsew signal tristate
rlabel metal2 s 56084 0 56140 800 6 la_data_out[117]
port 261 nsew signal tristate
rlabel metal2 s 56468 0 56524 800 6 la_data_out[118]
port 262 nsew signal tristate
rlabel metal2 s 56756 0 56812 800 6 la_data_out[119]
port 263 nsew signal tristate
rlabel metal2 s 17108 0 17164 800 6 la_data_out[11]
port 264 nsew signal tristate
rlabel metal2 s 57140 0 57196 800 6 la_data_out[120]
port 265 nsew signal tristate
rlabel metal2 s 57524 0 57580 800 6 la_data_out[121]
port 266 nsew signal tristate
rlabel metal2 s 57908 0 57964 800 6 la_data_out[122]
port 267 nsew signal tristate
rlabel metal2 s 58292 0 58348 800 6 la_data_out[123]
port 268 nsew signal tristate
rlabel metal2 s 58580 0 58636 800 6 la_data_out[124]
port 269 nsew signal tristate
rlabel metal2 s 58964 0 59020 800 6 la_data_out[125]
port 270 nsew signal tristate
rlabel metal2 s 59348 0 59404 800 6 la_data_out[126]
port 271 nsew signal tristate
rlabel metal2 s 59732 0 59788 800 6 la_data_out[127]
port 272 nsew signal tristate
rlabel metal2 s 17492 0 17548 800 6 la_data_out[12]
port 273 nsew signal tristate
rlabel metal2 s 17876 0 17932 800 6 la_data_out[13]
port 274 nsew signal tristate
rlabel metal2 s 18260 0 18316 800 6 la_data_out[14]
port 275 nsew signal tristate
rlabel metal2 s 18548 0 18604 800 6 la_data_out[15]
port 276 nsew signal tristate
rlabel metal2 s 18932 0 18988 800 6 la_data_out[16]
port 277 nsew signal tristate
rlabel metal2 s 19316 0 19372 800 6 la_data_out[17]
port 278 nsew signal tristate
rlabel metal2 s 19700 0 19756 800 6 la_data_out[18]
port 279 nsew signal tristate
rlabel metal2 s 20084 0 20140 800 6 la_data_out[19]
port 280 nsew signal tristate
rlabel metal2 s 13460 0 13516 800 6 la_data_out[1]
port 281 nsew signal tristate
rlabel metal2 s 20468 0 20524 800 6 la_data_out[20]
port 282 nsew signal tristate
rlabel metal2 s 20756 0 20812 800 6 la_data_out[21]
port 283 nsew signal tristate
rlabel metal2 s 21140 0 21196 800 6 la_data_out[22]
port 284 nsew signal tristate
rlabel metal2 s 21524 0 21580 800 6 la_data_out[23]
port 285 nsew signal tristate
rlabel metal2 s 21908 0 21964 800 6 la_data_out[24]
port 286 nsew signal tristate
rlabel metal2 s 22292 0 22348 800 6 la_data_out[25]
port 287 nsew signal tristate
rlabel metal2 s 22580 0 22636 800 6 la_data_out[26]
port 288 nsew signal tristate
rlabel metal2 s 22964 0 23020 800 6 la_data_out[27]
port 289 nsew signal tristate
rlabel metal2 s 23348 0 23404 800 6 la_data_out[28]
port 290 nsew signal tristate
rlabel metal2 s 23732 0 23788 800 6 la_data_out[29]
port 291 nsew signal tristate
rlabel metal2 s 13844 0 13900 800 6 la_data_out[2]
port 292 nsew signal tristate
rlabel metal2 s 24116 0 24172 800 6 la_data_out[30]
port 293 nsew signal tristate
rlabel metal2 s 24500 0 24556 800 6 la_data_out[31]
port 294 nsew signal tristate
rlabel metal2 s 24788 0 24844 800 6 la_data_out[32]
port 295 nsew signal tristate
rlabel metal2 s 25172 0 25228 800 6 la_data_out[33]
port 296 nsew signal tristate
rlabel metal2 s 25556 0 25612 800 6 la_data_out[34]
port 297 nsew signal tristate
rlabel metal2 s 25940 0 25996 800 6 la_data_out[35]
port 298 nsew signal tristate
rlabel metal2 s 26324 0 26380 800 6 la_data_out[36]
port 299 nsew signal tristate
rlabel metal2 s 26708 0 26764 800 6 la_data_out[37]
port 300 nsew signal tristate
rlabel metal2 s 26996 0 27052 800 6 la_data_out[38]
port 301 nsew signal tristate
rlabel metal2 s 27380 0 27436 800 6 la_data_out[39]
port 302 nsew signal tristate
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 303 nsew signal tristate
rlabel metal2 s 27764 0 27820 800 6 la_data_out[40]
port 304 nsew signal tristate
rlabel metal2 s 28148 0 28204 800 6 la_data_out[41]
port 305 nsew signal tristate
rlabel metal2 s 28532 0 28588 800 6 la_data_out[42]
port 306 nsew signal tristate
rlabel metal2 s 28916 0 28972 800 6 la_data_out[43]
port 307 nsew signal tristate
rlabel metal2 s 29204 0 29260 800 6 la_data_out[44]
port 308 nsew signal tristate
rlabel metal2 s 29588 0 29644 800 6 la_data_out[45]
port 309 nsew signal tristate
rlabel metal2 s 29972 0 30028 800 6 la_data_out[46]
port 310 nsew signal tristate
rlabel metal2 s 30356 0 30412 800 6 la_data_out[47]
port 311 nsew signal tristate
rlabel metal2 s 30740 0 30796 800 6 la_data_out[48]
port 312 nsew signal tristate
rlabel metal2 s 31028 0 31084 800 6 la_data_out[49]
port 313 nsew signal tristate
rlabel metal2 s 14516 0 14572 800 6 la_data_out[4]
port 314 nsew signal tristate
rlabel metal2 s 31412 0 31468 800 6 la_data_out[50]
port 315 nsew signal tristate
rlabel metal2 s 31796 0 31852 800 6 la_data_out[51]
port 316 nsew signal tristate
rlabel metal2 s 32180 0 32236 800 6 la_data_out[52]
port 317 nsew signal tristate
rlabel metal2 s 32564 0 32620 800 6 la_data_out[53]
port 318 nsew signal tristate
rlabel metal2 s 32948 0 33004 800 6 la_data_out[54]
port 319 nsew signal tristate
rlabel metal2 s 33236 0 33292 800 6 la_data_out[55]
port 320 nsew signal tristate
rlabel metal2 s 33620 0 33676 800 6 la_data_out[56]
port 321 nsew signal tristate
rlabel metal2 s 34004 0 34060 800 6 la_data_out[57]
port 322 nsew signal tristate
rlabel metal2 s 34388 0 34444 800 6 la_data_out[58]
port 323 nsew signal tristate
rlabel metal2 s 34772 0 34828 800 6 la_data_out[59]
port 324 nsew signal tristate
rlabel metal2 s 14900 0 14956 800 6 la_data_out[5]
port 325 nsew signal tristate
rlabel metal2 s 35156 0 35212 800 6 la_data_out[60]
port 326 nsew signal tristate
rlabel metal2 s 35444 0 35500 800 6 la_data_out[61]
port 327 nsew signal tristate
rlabel metal2 s 35828 0 35884 800 6 la_data_out[62]
port 328 nsew signal tristate
rlabel metal2 s 36212 0 36268 800 6 la_data_out[63]
port 329 nsew signal tristate
rlabel metal2 s 36596 0 36652 800 6 la_data_out[64]
port 330 nsew signal tristate
rlabel metal2 s 36980 0 37036 800 6 la_data_out[65]
port 331 nsew signal tristate
rlabel metal2 s 37364 0 37420 800 6 la_data_out[66]
port 332 nsew signal tristate
rlabel metal2 s 37652 0 37708 800 6 la_data_out[67]
port 333 nsew signal tristate
rlabel metal2 s 38036 0 38092 800 6 la_data_out[68]
port 334 nsew signal tristate
rlabel metal2 s 38420 0 38476 800 6 la_data_out[69]
port 335 nsew signal tristate
rlabel metal2 s 15284 0 15340 800 6 la_data_out[6]
port 336 nsew signal tristate
rlabel metal2 s 38804 0 38860 800 6 la_data_out[70]
port 337 nsew signal tristate
rlabel metal2 s 39188 0 39244 800 6 la_data_out[71]
port 338 nsew signal tristate
rlabel metal2 s 39476 0 39532 800 6 la_data_out[72]
port 339 nsew signal tristate
rlabel metal2 s 39860 0 39916 800 6 la_data_out[73]
port 340 nsew signal tristate
rlabel metal2 s 40244 0 40300 800 6 la_data_out[74]
port 341 nsew signal tristate
rlabel metal2 s 40628 0 40684 800 6 la_data_out[75]
port 342 nsew signal tristate
rlabel metal2 s 41012 0 41068 800 6 la_data_out[76]
port 343 nsew signal tristate
rlabel metal2 s 41396 0 41452 800 6 la_data_out[77]
port 344 nsew signal tristate
rlabel metal2 s 41684 0 41740 800 6 la_data_out[78]
port 345 nsew signal tristate
rlabel metal2 s 42068 0 42124 800 6 la_data_out[79]
port 346 nsew signal tristate
rlabel metal2 s 15668 0 15724 800 6 la_data_out[7]
port 347 nsew signal tristate
rlabel metal2 s 42452 0 42508 800 6 la_data_out[80]
port 348 nsew signal tristate
rlabel metal2 s 42836 0 42892 800 6 la_data_out[81]
port 349 nsew signal tristate
rlabel metal2 s 43220 0 43276 800 6 la_data_out[82]
port 350 nsew signal tristate
rlabel metal2 s 43604 0 43660 800 6 la_data_out[83]
port 351 nsew signal tristate
rlabel metal2 s 43892 0 43948 800 6 la_data_out[84]
port 352 nsew signal tristate
rlabel metal2 s 44276 0 44332 800 6 la_data_out[85]
port 353 nsew signal tristate
rlabel metal2 s 44660 0 44716 800 6 la_data_out[86]
port 354 nsew signal tristate
rlabel metal2 s 45044 0 45100 800 6 la_data_out[87]
port 355 nsew signal tristate
rlabel metal2 s 45428 0 45484 800 6 la_data_out[88]
port 356 nsew signal tristate
rlabel metal2 s 45812 0 45868 800 6 la_data_out[89]
port 357 nsew signal tristate
rlabel metal2 s 16052 0 16108 800 6 la_data_out[8]
port 358 nsew signal tristate
rlabel metal2 s 46100 0 46156 800 6 la_data_out[90]
port 359 nsew signal tristate
rlabel metal2 s 46484 0 46540 800 6 la_data_out[91]
port 360 nsew signal tristate
rlabel metal2 s 46868 0 46924 800 6 la_data_out[92]
port 361 nsew signal tristate
rlabel metal2 s 47252 0 47308 800 6 la_data_out[93]
port 362 nsew signal tristate
rlabel metal2 s 47636 0 47692 800 6 la_data_out[94]
port 363 nsew signal tristate
rlabel metal2 s 48020 0 48076 800 6 la_data_out[95]
port 364 nsew signal tristate
rlabel metal2 s 48308 0 48364 800 6 la_data_out[96]
port 365 nsew signal tristate
rlabel metal2 s 48692 0 48748 800 6 la_data_out[97]
port 366 nsew signal tristate
rlabel metal2 s 49076 0 49132 800 6 la_data_out[98]
port 367 nsew signal tristate
rlabel metal2 s 49460 0 49516 800 6 la_data_out[99]
port 368 nsew signal tristate
rlabel metal2 s 16340 0 16396 800 6 la_data_out[9]
port 369 nsew signal tristate
rlabel metal2 s 13172 0 13228 800 6 la_oen[0]
port 370 nsew signal input
rlabel metal2 s 49940 0 49996 800 6 la_oen[100]
port 371 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oen[101]
port 372 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oen[102]
port 373 nsew signal input
rlabel metal2 s 50996 0 51052 800 6 la_oen[103]
port 374 nsew signal input
rlabel metal2 s 51380 0 51436 800 6 la_oen[104]
port 375 nsew signal input
rlabel metal2 s 51764 0 51820 800 6 la_oen[105]
port 376 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oen[106]
port 377 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oen[107]
port 378 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oen[108]
port 379 nsew signal input
rlabel metal2 s 53204 0 53260 800 6 la_oen[109]
port 380 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_oen[10]
port 381 nsew signal input
rlabel metal2 s 53588 0 53644 800 6 la_oen[110]
port 382 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oen[111]
port 383 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oen[112]
port 384 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oen[113]
port 385 nsew signal input
rlabel metal2 s 55028 0 55084 800 6 la_oen[114]
port 386 nsew signal input
rlabel metal2 s 55412 0 55468 800 6 la_oen[115]
port 387 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oen[116]
port 388 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oen[117]
port 389 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oen[118]
port 390 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oen[119]
port 391 nsew signal input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 392 nsew signal input
rlabel metal2 s 57236 0 57292 800 6 la_oen[120]
port 393 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oen[121]
port 394 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oen[122]
port 395 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oen[123]
port 396 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oen[124]
port 397 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oen[125]
port 398 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oen[126]
port 399 nsew signal input
rlabel metal2 s 59828 0 59884 800 6 la_oen[127]
port 400 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_oen[12]
port 401 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_oen[13]
port 402 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_oen[14]
port 403 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_oen[15]
port 404 nsew signal input
rlabel metal2 s 19028 0 19084 800 6 la_oen[16]
port 405 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 406 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_oen[18]
port 407 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_oen[19]
port 408 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_oen[1]
port 409 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_oen[20]
port 410 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_oen[21]
port 411 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_oen[22]
port 412 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 413 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_oen[24]
port 414 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_oen[25]
port 415 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_oen[26]
port 416 nsew signal input
rlabel metal2 s 23156 0 23212 800 6 la_oen[27]
port 417 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_oen[28]
port 418 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 419 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_oen[2]
port 420 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_oen[30]
port 421 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_oen[31]
port 422 nsew signal input
rlabel metal2 s 24980 0 25036 800 6 la_oen[32]
port 423 nsew signal input
rlabel metal2 s 25364 0 25420 800 6 la_oen[33]
port 424 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_oen[34]
port 425 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 426 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_oen[36]
port 427 nsew signal input
rlabel metal2 s 26804 0 26860 800 6 la_oen[37]
port 428 nsew signal input
rlabel metal2 s 27188 0 27244 800 6 la_oen[38]
port 429 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_oen[39]
port 430 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_oen[3]
port 431 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_oen[40]
port 432 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 433 nsew signal input
rlabel metal2 s 28628 0 28684 800 6 la_oen[42]
port 434 nsew signal input
rlabel metal2 s 29012 0 29068 800 6 la_oen[43]
port 435 nsew signal input
rlabel metal2 s 29396 0 29452 800 6 la_oen[44]
port 436 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_oen[45]
port 437 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_oen[46]
port 438 nsew signal input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 439 nsew signal input
rlabel metal2 s 30836 0 30892 800 6 la_oen[48]
port 440 nsew signal input
rlabel metal2 s 31220 0 31276 800 6 la_oen[49]
port 441 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_oen[4]
port 442 nsew signal input
rlabel metal2 s 31604 0 31660 800 6 la_oen[50]
port 443 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_oen[51]
port 444 nsew signal input
rlabel metal2 s 32276 0 32332 800 6 la_oen[52]
port 445 nsew signal input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 446 nsew signal input
rlabel metal2 s 33044 0 33100 800 6 la_oen[54]
port 447 nsew signal input
rlabel metal2 s 33428 0 33484 800 6 la_oen[55]
port 448 nsew signal input
rlabel metal2 s 33812 0 33868 800 6 la_oen[56]
port 449 nsew signal input
rlabel metal2 s 34100 0 34156 800 6 la_oen[57]
port 450 nsew signal input
rlabel metal2 s 34484 0 34540 800 6 la_oen[58]
port 451 nsew signal input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 452 nsew signal input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 453 nsew signal input
rlabel metal2 s 35252 0 35308 800 6 la_oen[60]
port 454 nsew signal input
rlabel metal2 s 35636 0 35692 800 6 la_oen[61]
port 455 nsew signal input
rlabel metal2 s 36020 0 36076 800 6 la_oen[62]
port 456 nsew signal input
rlabel metal2 s 36308 0 36364 800 6 la_oen[63]
port 457 nsew signal input
rlabel metal2 s 36692 0 36748 800 6 la_oen[64]
port 458 nsew signal input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 459 nsew signal input
rlabel metal2 s 37460 0 37516 800 6 la_oen[66]
port 460 nsew signal input
rlabel metal2 s 37844 0 37900 800 6 la_oen[67]
port 461 nsew signal input
rlabel metal2 s 38132 0 38188 800 6 la_oen[68]
port 462 nsew signal input
rlabel metal2 s 38516 0 38572 800 6 la_oen[69]
port 463 nsew signal input
rlabel metal2 s 15380 0 15436 800 6 la_oen[6]
port 464 nsew signal input
rlabel metal2 s 38900 0 38956 800 6 la_oen[70]
port 465 nsew signal input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 466 nsew signal input
rlabel metal2 s 39668 0 39724 800 6 la_oen[72]
port 467 nsew signal input
rlabel metal2 s 40052 0 40108 800 6 la_oen[73]
port 468 nsew signal input
rlabel metal2 s 40340 0 40396 800 6 la_oen[74]
port 469 nsew signal input
rlabel metal2 s 40724 0 40780 800 6 la_oen[75]
port 470 nsew signal input
rlabel metal2 s 41108 0 41164 800 6 la_oen[76]
port 471 nsew signal input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 472 nsew signal input
rlabel metal2 s 41876 0 41932 800 6 la_oen[78]
port 473 nsew signal input
rlabel metal2 s 42260 0 42316 800 6 la_oen[79]
port 474 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_oen[7]
port 475 nsew signal input
rlabel metal2 s 42548 0 42604 800 6 la_oen[80]
port 476 nsew signal input
rlabel metal2 s 42932 0 42988 800 6 la_oen[81]
port 477 nsew signal input
rlabel metal2 s 43316 0 43372 800 6 la_oen[82]
port 478 nsew signal input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 479 nsew signal input
rlabel metal2 s 44084 0 44140 800 6 la_oen[84]
port 480 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oen[85]
port 481 nsew signal input
rlabel metal2 s 44756 0 44812 800 6 la_oen[86]
port 482 nsew signal input
rlabel metal2 s 45140 0 45196 800 6 la_oen[87]
port 483 nsew signal input
rlabel metal2 s 45524 0 45580 800 6 la_oen[88]
port 484 nsew signal input
rlabel metal2 s 45908 0 45964 800 6 la_oen[89]
port 485 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_oen[8]
port 486 nsew signal input
rlabel metal2 s 46292 0 46348 800 6 la_oen[90]
port 487 nsew signal input
rlabel metal2 s 46580 0 46636 800 6 la_oen[91]
port 488 nsew signal input
rlabel metal2 s 46964 0 47020 800 6 la_oen[92]
port 489 nsew signal input
rlabel metal2 s 47348 0 47404 800 6 la_oen[93]
port 490 nsew signal input
rlabel metal2 s 47732 0 47788 800 6 la_oen[94]
port 491 nsew signal input
rlabel metal2 s 48116 0 48172 800 6 la_oen[95]
port 492 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oen[96]
port 493 nsew signal input
rlabel metal2 s 48788 0 48844 800 6 la_oen[97]
port 494 nsew signal input
rlabel metal2 s 49172 0 49228 800 6 la_oen[98]
port 495 nsew signal input
rlabel metal2 s 49556 0 49612 800 6 la_oen[99]
port 496 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_oen[9]
port 497 nsew signal input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 498 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 499 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 500 nsew signal tristate
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 501 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_adr_i[10]
port 502 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 503 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 504 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 505 nsew signal input
rlabel metal2 s 6356 0 6412 800 6 wbs_adr_i[14]
port 506 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_adr_i[15]
port 507 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 508 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 509 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 510 nsew signal input
rlabel metal2 s 8180 0 8236 800 6 wbs_adr_i[19]
port 511 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 512 nsew signal input
rlabel metal2 s 8564 0 8620 800 6 wbs_adr_i[20]
port 513 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_adr_i[21]
port 514 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 515 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 516 nsew signal input
rlabel metal2 s 10004 0 10060 800 6 wbs_adr_i[24]
port 517 nsew signal input
rlabel metal2 s 10388 0 10444 800 6 wbs_adr_i[25]
port 518 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_adr_i[26]
port 519 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_adr_i[27]
port 520 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 521 nsew signal input
rlabel metal2 s 11828 0 11884 800 6 wbs_adr_i[29]
port 522 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 523 nsew signal input
rlabel metal2 s 12212 0 12268 800 6 wbs_adr_i[30]
port 524 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_adr_i[31]
port 525 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 526 nsew signal input
rlabel metal2 s 2708 0 2764 800 6 wbs_adr_i[4]
port 527 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 528 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 529 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 530 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 531 nsew signal input
rlabel metal2 s 4532 0 4588 800 6 wbs_adr_i[9]
port 532 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 533 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 534 nsew signal input
rlabel metal2 s 5012 0 5068 800 6 wbs_dat_i[10]
port 535 nsew signal input
rlabel metal2 s 5396 0 5452 800 6 wbs_dat_i[11]
port 536 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 537 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 538 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 539 nsew signal input
rlabel metal2 s 6836 0 6892 800 6 wbs_dat_i[15]
port 540 nsew signal input
rlabel metal2 s 7220 0 7276 800 6 wbs_dat_i[16]
port 541 nsew signal input
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_i[17]
port 542 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 543 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 544 nsew signal input
rlabel metal2 s 1364 0 1420 800 6 wbs_dat_i[1]
port 545 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 546 nsew signal input
rlabel metal2 s 9044 0 9100 800 6 wbs_dat_i[21]
port 547 nsew signal input
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_i[22]
port 548 nsew signal input
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_i[23]
port 549 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 550 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 551 nsew signal input
rlabel metal2 s 10868 0 10924 800 6 wbs_dat_i[26]
port 552 nsew signal input
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_i[27]
port 553 nsew signal input
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_i[28]
port 554 nsew signal input
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_i[29]
port 555 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 556 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 557 nsew signal input
rlabel metal2 s 12692 0 12748 800 6 wbs_dat_i[31]
port 558 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 559 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 560 nsew signal input
rlabel metal2 s 3188 0 3244 800 6 wbs_dat_i[5]
port 561 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 562 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 563 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 564 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 565 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 566 nsew signal tristate
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 567 nsew signal tristate
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 568 nsew signal tristate
rlabel metal2 s 5876 0 5932 800 6 wbs_dat_o[12]
port 569 nsew signal tristate
rlabel metal2 s 6260 0 6316 800 6 wbs_dat_o[13]
port 570 nsew signal tristate
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 571 nsew signal tristate
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 572 nsew signal tristate
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 573 nsew signal tristate
rlabel metal2 s 7700 0 7756 800 6 wbs_dat_o[17]
port 574 nsew signal tristate
rlabel metal2 s 8084 0 8140 800 6 wbs_dat_o[18]
port 575 nsew signal tristate
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_o[19]
port 576 nsew signal tristate
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 577 nsew signal tristate
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 578 nsew signal tristate
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 579 nsew signal tristate
rlabel metal2 s 9524 0 9580 800 6 wbs_dat_o[22]
port 580 nsew signal tristate
rlabel metal2 s 9908 0 9964 800 6 wbs_dat_o[23]
port 581 nsew signal tristate
rlabel metal2 s 10292 0 10348 800 6 wbs_dat_o[24]
port 582 nsew signal tristate
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 583 nsew signal tristate
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 584 nsew signal tristate
rlabel metal2 s 11348 0 11404 800 6 wbs_dat_o[27]
port 585 nsew signal tristate
rlabel metal2 s 11732 0 11788 800 6 wbs_dat_o[28]
port 586 nsew signal tristate
rlabel metal2 s 12116 0 12172 800 6 wbs_dat_o[29]
port 587 nsew signal tristate
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 588 nsew signal tristate
rlabel metal2 s 12500 0 12556 800 6 wbs_dat_o[30]
port 589 nsew signal tristate
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 590 nsew signal tristate
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 591 nsew signal tristate
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 592 nsew signal tristate
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 593 nsew signal tristate
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 594 nsew signal tristate
rlabel metal2 s 4052 0 4108 800 6 wbs_dat_o[7]
port 595 nsew signal tristate
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 596 nsew signal tristate
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 597 nsew signal tristate
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 598 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 599 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 600 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 601 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 602 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 603 nsew signal input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 604 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 606 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 607 nsew ground bidirectional
rlabel metal4 s 35636 2664 35956 57276 6 vccd2
port 608 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 57276 6 vccd2
port 609 nsew power bidirectional
rlabel metal4 s 50996 2664 51316 57276 6 vssd2
port 610 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 57276 6 vssd2
port 611 nsew ground bidirectional
rlabel metal4 s 36296 2664 36616 57276 6 vdda1
port 612 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 57276 6 vdda1
port 613 nsew power bidirectional
rlabel metal4 s 51656 2664 51976 57276 6 vssa1
port 614 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 57276 6 vssa1
port 615 nsew ground bidirectional
rlabel metal4 s 36956 2664 37276 57276 6 vdda2
port 616 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 57276 6 vdda2
port 617 nsew power bidirectional
rlabel metal4 s 52316 2664 52636 57276 6 vssa2
port 618 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 57276 6 vssa2
port 619 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
