magic
tech sky130A
magscale 1 2
timestamp 1624892585
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1728 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 1027 134 1085 146
rect 1027 132 1039 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 102 561 132
rect 303 68 367 102
rect 401 68 561 102
rect 303 48 561 68
rect 591 48 849 132
rect 879 100 1039 132
rect 1073 132 1085 134
rect 1073 100 1137 132
rect 879 48 1137 100
rect 1167 48 1425 132
rect 1455 102 1613 132
rect 1455 68 1519 102
rect 1553 68 1613 102
rect 1455 48 1613 68
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 598 561 618
rect 303 564 367 598
rect 401 564 561 598
rect 303 450 561 564
rect 591 450 849 618
rect 879 485 1137 618
rect 879 451 1039 485
rect 1073 451 1137 485
rect 879 450 1137 451
rect 1167 450 1425 618
rect 1455 598 1613 618
rect 1455 564 1519 598
rect 1553 564 1613 598
rect 1455 450 1613 564
rect 115 439 173 450
rect 1027 439 1085 450
<< ndiffc >>
rect 127 100 161 134
rect 367 68 401 102
rect 1039 100 1073 134
rect 1519 68 1553 102
<< pdiffc >>
rect 127 451 161 485
rect 367 564 401 598
rect 1039 451 1073 485
rect 1519 564 1553 598
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 31 618 1697 649
rect 351 598 417 618
rect 351 564 367 598
rect 401 564 417 598
rect 351 548 417 564
rect 1503 598 1569 618
rect 1503 564 1519 598
rect 1553 564 1569 598
rect 1503 548 1569 564
rect 111 485 177 501
rect 1023 485 1089 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 271 418 305 451
rect 1023 451 1039 485
rect 1073 451 1089 485
rect 1023 435 1089 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 1123 402 1185 418
rect 1123 401 1135 402
rect 831 352 897 368
rect 1119 368 1135 401
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 271 323 305 352
rect 559 296 593 352
rect 559 231 593 262
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 831 215 897 231
rect 543 181 559 215
rect 593 181 609 215
rect 689 181 847 215
rect 881 181 897 215
rect 1119 215 1185 231
rect 1119 184 1135 215
rect 543 165 609 181
rect 831 165 897 181
rect 1123 181 1135 184
rect 1169 181 1185 215
rect 1123 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 1023 134 1089 150
rect 111 84 177 100
rect 351 102 417 118
rect 351 68 367 102
rect 401 68 417 102
rect 1023 100 1039 134
rect 1073 100 1089 134
rect 1023 84 1089 100
rect 1503 102 1569 118
rect 351 48 417 68
rect 1503 68 1519 102
rect 1553 68 1569 102
rect 1503 48 1569 68
rect 31 17 1697 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 367 564 401 598
rect 1519 564 1553 598
rect 127 451 161 485
rect 271 451 305 485
rect 1039 451 1073 485
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 271 289 305 323
rect 559 262 593 296
rect 271 181 305 215
rect 655 181 689 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 127 100 161 134
rect 367 68 401 102
rect 1039 100 1073 134
rect 1519 68 1553 102
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 714
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 618 1728 649
rect 355 598 413 618
rect 355 564 367 598
rect 401 564 413 598
rect 355 552 413 564
rect 1507 598 1565 618
rect 1507 564 1519 598
rect 1553 564 1565 598
rect 1507 552 1565 564
rect 115 485 173 497
rect 115 451 127 485
rect 161 451 173 485
rect 115 439 173 451
rect 259 485 317 497
rect 259 451 271 485
rect 305 482 317 485
rect 1027 485 1085 497
rect 305 454 974 482
rect 305 451 317 454
rect 259 439 317 451
rect 130 399 158 439
rect 835 402 893 414
rect 835 399 847 402
rect 130 371 847 399
rect 130 146 158 371
rect 835 368 847 371
rect 881 368 893 402
rect 946 399 974 454
rect 1027 451 1039 485
rect 1073 482 1085 485
rect 1073 454 1262 482
rect 1073 451 1085 454
rect 1027 439 1085 451
rect 1123 402 1181 414
rect 1123 399 1135 402
rect 946 371 1135 399
rect 835 356 893 368
rect 1123 368 1135 371
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 259 323 317 335
rect 259 289 271 323
rect 305 289 317 323
rect 259 277 317 289
rect 547 296 605 308
rect 274 227 302 277
rect 547 262 559 296
rect 593 262 605 296
rect 547 250 605 262
rect 259 215 317 227
rect 259 181 271 215
rect 305 212 317 215
rect 643 215 701 227
rect 643 212 655 215
rect 305 184 655 212
rect 305 181 317 184
rect 259 169 317 181
rect 643 181 655 184
rect 689 181 701 215
rect 850 212 878 356
rect 1123 215 1181 227
rect 1123 212 1135 215
rect 850 184 1135 212
rect 643 169 701 181
rect 1123 181 1135 184
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 1027 134 1085 146
rect 115 88 173 100
rect 355 102 413 114
rect 355 68 367 102
rect 401 68 413 102
rect 1027 100 1039 134
rect 1073 131 1085 134
rect 1234 131 1262 454
rect 1411 402 1469 414
rect 1411 368 1423 402
rect 1457 368 1469 402
rect 1411 356 1469 368
rect 1426 227 1454 356
rect 1411 215 1469 227
rect 1411 181 1423 215
rect 1457 181 1469 215
rect 1411 169 1469 181
rect 1073 103 1262 131
rect 1073 100 1085 103
rect 1027 88 1085 100
rect 1507 102 1565 114
rect 355 48 413 68
rect 1507 68 1519 102
rect 1553 68 1565 102
rect 1507 48 1565 68
rect 0 17 1728 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -48 1728 -17
<< labels >>
rlabel metal1 0 618 1728 714 0 VDD
port 4 se
rlabel metal1 0 618 1728 714 0 VDD
port 4 se
rlabel metal1 0 -48 1728 48 0 GND
port 2 se
rlabel metal1 0 -48 1728 48 0 GND
port 2 se
rlabel metal1 1027 88 1085 103 0 Y
port 5 se
rlabel metal1 1027 103 1262 131 0 Y
port 5 se
rlabel metal1 1027 131 1085 146 0 Y
port 5 se
rlabel metal1 1027 439 1085 454 0 Y
port 5 se
rlabel metal1 1234 131 1262 454 0 Y
port 5 se
rlabel metal1 1027 454 1262 482 0 Y
port 5 se
rlabel metal1 1027 482 1085 497 0 Y
port 5 se
rlabel metal1 259 169 317 184 0 S
port 3 se
rlabel metal1 643 169 701 184 0 S
port 3 se
rlabel metal1 259 184 701 212 0 S
port 3 se
rlabel metal1 259 212 317 227 0 S
port 3 se
rlabel metal1 643 212 701 227 0 S
port 3 se
rlabel metal1 274 227 302 277 0 S
port 3 se
rlabel metal1 259 277 317 335 0 S
port 3 se
rlabel metal1 547 250 605 308 0 A
port 0 se
rlabel metal1 1411 169 1469 227 0 B
port 1 se
rlabel metal1 1426 227 1454 356 0 B
port 1 se
rlabel metal1 1411 356 1469 414 0 B
port 1 se
rlabel locali 0 -17 1728 17 4 GND
port 2 se ground default abutment
rlabel locali 31 17 1697 48 4 GND
port 2 se ground default abutment
rlabel locali 0 649 1728 683 4 VDD
port 4 se power default abutment
rlabel locali 31 618 1697 649 4 VDD
port 4 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1728 666
<< end >>
