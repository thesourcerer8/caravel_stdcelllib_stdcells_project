magic
tech sky130A
magscale 1 2
timestamp 1636809601
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 2304 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
rect 2001 48 2031 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
rect 2001 450 2031 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 643 134 701 146
rect 643 132 655 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 48 561 132
rect 591 100 655 132
rect 689 132 701 134
rect 1027 134 1085 146
rect 1027 132 1039 134
rect 689 100 849 132
rect 591 48 849 100
rect 879 100 1039 132
rect 1073 132 1085 134
rect 1219 134 1277 146
rect 1219 132 1231 134
rect 1073 100 1137 132
rect 879 48 1137 100
rect 1167 100 1231 132
rect 1265 132 1277 134
rect 1555 134 1613 146
rect 1555 132 1567 134
rect 1265 100 1425 132
rect 1167 48 1425 100
rect 1455 100 1567 132
rect 1601 100 1613 134
rect 1455 48 1613 100
rect 1843 134 1901 146
rect 1843 100 1855 134
rect 1889 132 1901 134
rect 2083 134 2141 146
rect 2083 132 2095 134
rect 1889 100 2001 132
rect 1843 48 2001 100
rect 2031 100 2095 132
rect 2129 132 2141 134
rect 2129 100 2189 132
rect 2031 48 2189 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 450 561 618
rect 591 593 849 618
rect 591 559 655 593
rect 689 559 849 593
rect 591 450 849 559
rect 879 485 1137 618
rect 879 451 1039 485
rect 1073 451 1137 485
rect 879 450 1137 451
rect 1167 593 1425 618
rect 1167 559 1231 593
rect 1265 559 1425 593
rect 1167 450 1425 559
rect 1455 485 1613 618
rect 1455 451 1567 485
rect 1601 451 1613 485
rect 1455 450 1613 451
rect 115 439 173 450
rect 1027 439 1085 450
rect 1555 439 1613 450
rect 1843 485 2001 618
rect 1843 451 1855 485
rect 1889 451 2001 485
rect 1843 450 2001 451
rect 2031 485 2189 618
rect 2031 451 2095 485
rect 2129 451 2189 485
rect 2031 450 2189 451
rect 1843 439 1901 450
rect 2083 439 2141 450
<< ndiffc >>
rect 127 100 161 134
rect 655 100 689 134
rect 1039 100 1073 134
rect 1231 100 1265 134
rect 1567 100 1601 134
rect 1855 100 1889 134
rect 2095 100 2129 134
<< pdiffc >>
rect 127 451 161 485
rect 655 559 689 593
rect 1039 451 1073 485
rect 1231 559 1265 593
rect 1567 451 1601 485
rect 1855 451 1889 485
rect 2095 451 2129 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 2001 618 2031 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 2001 418 2031 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 2001 132 2031 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
rect 2001 22 2031 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1999 368 2033 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1999 181 2033 215
<< locali >>
rect 0 649 1231 683
rect 1265 649 2304 683
rect 31 643 2273 649
rect 31 618 1181 643
rect 1315 618 2273 643
rect 639 593 705 618
rect 639 559 655 593
rect 689 559 705 593
rect 639 543 705 559
rect 1215 593 1281 609
rect 1215 559 1231 593
rect 1265 559 1281 593
rect 1215 543 1281 559
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 1023 485 1089 501
rect 1023 451 1039 485
rect 1073 452 1089 485
rect 1551 485 1617 501
rect 1073 451 1085 452
rect 1023 435 1085 451
rect 1551 451 1567 485
rect 1601 451 1617 485
rect 1551 435 1617 451
rect 1839 485 1905 501
rect 1839 451 1855 485
rect 1889 451 1905 485
rect 2079 485 2145 501
rect 2079 452 2095 485
rect 1839 435 1905 451
rect 2083 451 2095 452
rect 2129 451 2145 485
rect 2083 435 2145 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 559 231 593 352
rect 847 231 881 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 184 609 215
rect 831 215 897 231
rect 593 181 605 184
rect 543 165 605 181
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 184 1185 215
rect 1407 215 1473 231
rect 1169 181 1181 184
rect 1119 165 1181 181
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1567 215 1601 435
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 1999 231 2033 352
rect 1567 150 1601 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 639 134 705 150
rect 639 100 655 134
rect 689 100 705 134
rect 639 84 705 100
rect 1023 134 1085 150
rect 1023 100 1039 134
rect 1073 131 1085 134
rect 1215 134 1281 150
rect 1073 100 1089 131
rect 1023 84 1089 100
rect 1215 100 1231 134
rect 1265 100 1281 134
rect 1215 84 1281 100
rect 1551 134 1617 150
rect 1551 100 1567 134
rect 1601 100 1617 134
rect 1551 84 1617 100
rect 1839 134 1905 150
rect 1839 100 1855 134
rect 1889 100 1905 134
rect 2083 134 2145 150
rect 2083 131 2095 134
rect 1839 84 1905 100
rect 2079 100 2095 131
rect 2129 100 2145 134
rect 2079 84 2145 100
rect 1231 48 1265 84
rect 31 17 2273 48
rect 0 -17 655 17
rect 689 -17 2304 17
<< viali >>
rect 1231 649 1265 683
rect 655 559 689 593
rect 1231 559 1265 593
rect 127 451 161 485
rect 1039 451 1073 485
rect 1855 451 1889 485
rect 2095 451 2129 485
rect 271 368 305 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1567 181 1601 215
rect 1999 181 2033 215
rect 127 100 161 134
rect 655 100 689 134
rect 1039 100 1073 134
rect 1855 100 1889 134
rect 2095 100 2129 134
rect 655 -17 689 17
<< metal1 >>
rect 0 683 2304 714
rect 0 649 1231 683
rect 1265 649 2304 683
rect 0 618 2304 649
rect 643 593 701 618
rect 643 559 655 593
rect 689 559 701 593
rect 643 547 701 559
rect 1219 593 1277 618
rect 1219 559 1231 593
rect 1265 559 1277 593
rect 1219 547 1277 559
rect 115 485 173 497
rect 115 451 127 485
rect 161 451 173 485
rect 115 439 173 451
rect 1027 485 1085 497
rect 1027 451 1039 485
rect 1073 482 1085 485
rect 1843 485 1901 497
rect 1843 482 1855 485
rect 1073 454 1855 482
rect 1073 451 1085 454
rect 1027 439 1085 451
rect 1843 451 1855 454
rect 1889 451 1901 485
rect 1843 439 1901 451
rect 2083 485 2141 497
rect 2083 451 2095 485
rect 2129 451 2141 485
rect 2083 439 2141 451
rect 130 146 158 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 399 317 402
rect 1123 402 1181 414
rect 1123 399 1135 402
rect 305 371 1135 399
rect 305 368 317 371
rect 259 356 317 368
rect 1123 368 1135 371
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 1411 402 1469 414
rect 1411 368 1423 402
rect 1457 399 1469 402
rect 2098 399 2126 439
rect 1457 371 2126 399
rect 1457 368 1469 371
rect 1411 356 1469 368
rect 274 227 302 356
rect 1138 227 1166 356
rect 1426 227 1454 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 212 605 215
rect 835 215 893 227
rect 835 212 847 215
rect 593 184 847 212
rect 593 181 605 184
rect 547 169 605 181
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 1411 215 1469 227
rect 1411 181 1423 215
rect 1457 181 1469 215
rect 1411 169 1469 181
rect 1555 215 1613 227
rect 1555 181 1567 215
rect 1601 212 1613 215
rect 1987 215 2045 227
rect 1987 212 1999 215
rect 1601 184 1999 212
rect 1601 181 1613 184
rect 1555 169 1613 181
rect 1987 181 1999 184
rect 2033 181 2045 215
rect 1987 169 2045 181
rect 2098 146 2126 371
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 643 134 701 146
rect 643 100 655 134
rect 689 100 701 134
rect 643 88 701 100
rect 1027 134 1085 146
rect 1027 100 1039 134
rect 1073 131 1085 134
rect 1843 134 1901 146
rect 1843 131 1855 134
rect 1073 103 1855 131
rect 1073 100 1085 103
rect 1027 88 1085 100
rect 1843 100 1855 103
rect 1889 100 1901 134
rect 1843 88 1901 100
rect 2083 134 2141 146
rect 2083 100 2095 134
rect 2129 100 2141 134
rect 2083 88 2141 100
rect 658 48 686 88
rect 0 17 2304 48
rect 0 -17 655 17
rect 689 -17 2304 17
rect 0 -48 2304 -17
<< labels >>
rlabel metal1 0 618 2304 714 0 VPWR
port 4 se
rlabel metal1 0 618 2304 714 0 VPWR
port 4 se
rlabel metal1 0 -48 2304 48 0 VGND
port 3 se
rlabel metal1 0 -48 2304 48 0 VGND
port 3 se
rlabel metal1 1555 169 1613 184 0 C
port 2 se
rlabel metal1 1987 169 2045 184 0 C
port 2 se
rlabel metal1 1555 184 2045 212 0 C
port 2 se
rlabel metal1 1555 212 1613 227 0 C
port 2 se
rlabel metal1 1987 212 2045 227 0 C
port 2 se
rlabel metal1 259 169 317 227 0 B
port 1 se
rlabel metal1 1123 169 1181 227 0 B
port 1 se
rlabel metal1 274 227 302 356 0 B
port 1 se
rlabel metal1 1138 227 1166 356 0 B
port 1 se
rlabel metal1 259 356 317 371 0 B
port 1 se
rlabel metal1 1123 356 1181 371 0 B
port 1 se
rlabel metal1 259 371 1181 399 0 B
port 1 se
rlabel metal1 259 399 317 414 0 B
port 1 se
rlabel metal1 1123 399 1181 414 0 B
port 1 se
rlabel metal1 547 169 605 184 0 A
port 0 se
rlabel metal1 835 169 893 184 0 A
port 0 se
rlabel metal1 547 184 893 212 0 A
port 0 se
rlabel metal1 547 212 605 227 0 A
port 0 se
rlabel metal1 835 212 893 227 0 A
port 0 se
rlabel locali 0 -17 2304 17 4 VGND
port 3 se ground default abutment
rlabel locali 31 17 2273 48 4 VGND
port 3 se ground default abutment
rlabel locali 0 649 2304 683 4 VPWR
port 4 se power default abutment
rlabel metal1 31 618 2273 649 4 VGND
port 3 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 2304 666
<< end >>
