magic
tech sky130A
timestamp 1621277170
<< end >>
