VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.840 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 15.840 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.840 0.240 ;
    END
  END gnd
  PIN YS
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 14.740 2.150 15.030 2.440 ;
        RECT 14.810 0.690 14.950 2.150 ;
        RECT 14.740 0.400 15.030 0.690 ;
    END
  END YS
  PIN YC
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.150 0.870 2.440 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 0.580 0.400 0.870 0.690 ;
    END
  END YC
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.750 5.910 2.040 ;
        RECT 5.690 1.090 5.830 1.750 ;
        RECT 5.620 0.800 5.910 1.090 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.750 4.470 2.040 ;
        RECT 9.940 1.750 10.230 2.040 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 10.010 1.090 10.150 1.750 ;
        RECT 4.180 0.800 4.470 1.090 ;
        RECT 9.940 0.800 10.230 1.090 ;
        RECT 4.250 0.610 4.390 0.800 ;
        RECT 10.010 0.610 10.150 0.800 ;
        RECT 4.250 0.470 10.150 0.610 ;
    END
  END B
END HAX1
END LIBRARY

