magic
tech sky130A
timestamp 1624065832
<< nwell >>
rect 0 179 1584 333
<< nmos >>
rect 137 24 152 66
rect 425 24 440 66
rect 569 24 584 66
rect 857 24 872 66
rect 1001 24 1016 66
rect 1145 24 1160 66
rect 1433 24 1448 66
<< pmos >>
rect 137 225 152 309
rect 425 225 440 309
rect 569 225 584 309
rect 857 225 872 309
rect 1001 225 1016 309
rect 1145 225 1160 309
rect 1433 225 1448 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 346 67 375 73
rect 81 50 137 66
rect 58 24 137 50
rect 152 49 231 66
rect 152 32 184 49
rect 201 32 231 49
rect 152 24 231 32
rect 346 50 352 67
rect 369 66 375 67
rect 946 67 975 73
rect 946 66 952 67
rect 369 50 425 66
rect 346 24 425 50
rect 440 24 569 66
rect 584 49 663 66
rect 584 32 616 49
rect 633 32 663 49
rect 584 24 663 32
rect 778 49 857 66
rect 778 32 784 49
rect 801 32 857 49
rect 778 24 857 32
rect 872 50 952 66
rect 969 66 975 67
rect 1042 67 1071 73
rect 1042 66 1048 67
rect 969 50 1001 66
rect 872 24 1001 50
rect 1016 50 1048 66
rect 1065 66 1071 67
rect 1186 67 1215 73
rect 1186 66 1192 67
rect 1065 50 1145 66
rect 1016 24 1145 50
rect 1160 50 1192 66
rect 1209 66 1215 67
rect 1474 67 1503 73
rect 1474 66 1480 67
rect 1209 50 1239 66
rect 1160 24 1239 50
rect 1354 49 1433 66
rect 1354 32 1360 49
rect 1377 32 1433 49
rect 1354 24 1433 32
rect 1448 50 1480 66
rect 1497 66 1503 67
rect 1497 50 1527 66
rect 1448 24 1527 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 301 231 309
rect 152 284 184 301
rect 201 284 231 301
rect 152 225 231 284
rect 346 243 425 309
rect 346 226 352 243
rect 369 226 425 243
rect 346 225 425 226
rect 440 301 569 309
rect 440 284 472 301
rect 489 284 569 301
rect 440 225 569 284
rect 584 243 663 309
rect 584 226 616 243
rect 633 226 663 243
rect 584 225 663 226
rect 778 301 857 309
rect 778 284 784 301
rect 801 284 857 301
rect 778 225 857 284
rect 872 243 1001 309
rect 872 226 952 243
rect 969 226 1001 243
rect 872 225 1001 226
rect 1016 225 1145 309
rect 1160 301 1239 309
rect 1160 284 1192 301
rect 1209 284 1239 301
rect 1160 225 1239 284
rect 1354 301 1433 309
rect 1354 284 1360 301
rect 1377 284 1433 301
rect 1354 225 1433 284
rect 1448 243 1527 309
rect 1448 226 1480 243
rect 1497 226 1527 243
rect 1448 225 1527 226
rect 58 220 87 225
rect 346 220 375 225
rect 610 220 639 225
rect 946 220 975 225
rect 1474 220 1503 225
<< ndiffc >>
rect 64 50 81 67
rect 184 32 201 49
rect 352 50 369 67
rect 616 32 633 49
rect 784 32 801 49
rect 952 50 969 67
rect 1048 50 1065 67
rect 1192 50 1209 67
rect 1360 32 1377 49
rect 1480 50 1497 67
<< pdiffc >>
rect 64 226 81 243
rect 184 284 201 301
rect 352 226 369 243
rect 472 284 489 301
rect 616 226 633 243
rect 784 284 801 301
rect 952 226 969 243
rect 1192 284 1209 301
rect 1360 284 1377 301
rect 1480 226 1497 243
<< poly >>
rect 137 309 152 322
rect 425 309 440 322
rect 569 309 584 322
rect 857 309 872 322
rect 1001 309 1016 322
rect 1145 309 1160 322
rect 1433 309 1448 322
rect 137 209 152 225
rect 425 209 440 225
rect 569 209 584 225
rect 857 209 872 225
rect 1001 209 1016 225
rect 1145 209 1160 225
rect 1433 209 1448 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 848 201 881 209
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 992 201 1025 209
rect 992 184 1000 201
rect 1017 184 1025 201
rect 992 176 1025 184
rect 1136 201 1169 209
rect 1136 184 1144 201
rect 1161 184 1169 201
rect 1136 176 1169 184
rect 1424 201 1457 209
rect 1424 184 1432 201
rect 1449 184 1457 201
rect 1424 176 1457 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 848 108 881 116
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 992 108 1025 116
rect 992 91 1000 108
rect 1017 91 1025 108
rect 992 83 1025 91
rect 1136 108 1169 116
rect 1136 91 1144 108
rect 1161 91 1169 108
rect 1136 83 1169 91
rect 1424 108 1457 116
rect 1424 91 1432 108
rect 1449 91 1457 108
rect 1424 83 1457 91
rect 137 66 152 83
rect 425 66 440 83
rect 569 66 584 83
rect 857 66 872 83
rect 1001 66 1016 83
rect 1145 66 1160 83
rect 1433 66 1448 83
rect 137 11 152 24
rect 425 11 440 24
rect 569 11 584 24
rect 857 11 872 24
rect 1001 11 1016 24
rect 1145 11 1160 24
rect 1433 11 1448 24
<< polycont >>
rect 136 184 153 201
rect 424 184 441 201
rect 568 184 585 201
rect 856 184 873 201
rect 1000 184 1017 201
rect 1144 184 1161 201
rect 1432 184 1449 201
rect 136 91 153 108
rect 424 91 441 108
rect 568 91 585 108
rect 856 91 873 108
rect 1000 91 1017 108
rect 1144 91 1161 108
rect 1432 91 1449 108
<< locali >>
rect 176 301 209 309
rect 176 284 184 301
rect 201 284 209 301
rect 176 276 209 284
rect 464 301 497 309
rect 464 284 472 301
rect 489 284 497 301
rect 464 276 497 284
rect 776 301 809 309
rect 776 284 784 301
rect 801 284 809 301
rect 776 276 809 284
rect 1184 301 1217 309
rect 1184 284 1192 301
rect 1209 284 1217 301
rect 1184 276 1217 284
rect 1352 301 1385 309
rect 1352 284 1360 301
rect 1377 284 1385 301
rect 1352 276 1385 284
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 344 243 377 251
rect 344 226 352 243
rect 369 226 377 243
rect 344 218 377 226
rect 608 243 641 251
rect 608 226 616 243
rect 633 226 641 243
rect 608 218 641 226
rect 944 243 977 251
rect 944 226 952 243
rect 969 226 977 243
rect 1472 243 1505 251
rect 1472 226 1480 243
rect 1497 226 1505 243
rect 944 218 975 226
rect 1474 218 1505 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 591 209
rect 848 201 881 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 992 201 1025 209
rect 992 176 1000 201
rect 856 116 873 176
rect 1017 176 1025 201
rect 1136 201 1169 209
rect 1000 116 1017 172
rect 1136 184 1144 201
rect 1161 184 1169 201
rect 1136 176 1169 184
rect 1424 201 1457 209
rect 1424 184 1432 201
rect 1449 184 1457 201
rect 1424 176 1457 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 848 108 881 116
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 992 108 1025 116
rect 992 91 1000 108
rect 1017 92 1025 108
rect 1017 91 1023 92
rect 992 83 1023 91
rect 1048 75 1065 172
rect 1136 108 1169 116
rect 1136 91 1144 108
rect 1161 91 1169 108
rect 1136 83 1169 91
rect 1424 108 1457 116
rect 1424 91 1432 108
rect 1449 92 1457 108
rect 1449 91 1455 92
rect 1424 83 1455 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 344 67 377 75
rect 56 42 89 50
rect 176 49 209 57
rect 176 32 184 49
rect 201 32 209 49
rect 344 50 352 67
rect 369 50 377 67
rect 944 67 975 75
rect 344 42 377 50
rect 608 49 641 57
rect 176 24 209 32
rect 608 32 616 49
rect 633 32 641 49
rect 608 27 641 32
rect 608 24 616 27
rect 633 24 641 27
rect 776 49 809 57
rect 776 32 784 49
rect 801 32 809 49
rect 944 50 952 67
rect 969 66 975 67
rect 1040 67 1073 75
rect 969 50 977 66
rect 944 42 977 50
rect 1040 50 1048 67
rect 1065 50 1073 67
rect 1186 67 1217 75
rect 1186 66 1192 67
rect 1040 42 1073 50
rect 1184 50 1192 66
rect 1209 50 1217 67
rect 1472 67 1505 75
rect 1184 42 1217 50
rect 1352 49 1385 57
rect 776 27 809 32
rect 776 24 784 27
rect 801 24 809 27
rect 1352 32 1360 49
rect 1377 32 1385 49
rect 1472 50 1480 67
rect 1497 50 1505 67
rect 1472 42 1505 50
rect 1352 24 1385 32
<< viali >>
rect 184 284 201 301
rect 472 284 489 301
rect 784 284 801 301
rect 1192 284 1209 301
rect 1360 284 1377 301
rect 64 226 81 243
rect 352 226 369 243
rect 616 226 633 243
rect 952 226 969 243
rect 1480 226 1497 243
rect 136 184 153 201
rect 424 184 441 201
rect 568 184 585 201
rect 856 184 873 201
rect 1000 184 1017 201
rect 1000 172 1017 184
rect 1048 172 1065 189
rect 1144 184 1161 201
rect 1432 184 1449 201
rect 136 91 153 108
rect 424 91 441 108
rect 568 91 585 108
rect 1000 91 1017 108
rect 1144 91 1161 108
rect 1432 91 1449 108
rect 64 50 81 67
rect 184 32 201 49
rect 352 50 369 67
rect 616 10 633 27
rect 952 50 969 67
rect 1192 50 1209 67
rect 784 10 801 27
rect 1360 32 1377 49
rect 1480 50 1497 67
<< metal1 >>
rect 0 309 1584 357
rect 178 301 207 309
rect 178 284 184 301
rect 201 284 207 301
rect 178 278 207 284
rect 466 301 495 309
rect 466 284 472 301
rect 489 284 495 301
rect 466 278 495 284
rect 778 301 807 309
rect 778 284 784 301
rect 801 284 807 301
rect 778 278 807 284
rect 1186 301 1215 309
rect 1186 284 1192 301
rect 1209 284 1215 301
rect 1186 278 1215 284
rect 1354 301 1383 309
rect 1354 284 1360 301
rect 1377 284 1383 301
rect 1354 278 1383 284
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 58 220 87 226
rect 346 243 375 249
rect 346 226 352 243
rect 369 241 375 243
rect 610 243 639 249
rect 610 241 616 243
rect 369 227 616 241
rect 369 226 375 227
rect 346 220 375 226
rect 610 226 616 227
rect 633 241 639 243
rect 946 243 975 249
rect 633 227 871 241
rect 633 226 639 227
rect 610 220 639 226
rect 65 73 79 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 200 159 201
rect 353 200 367 220
rect 857 207 871 227
rect 946 226 952 243
rect 969 241 975 243
rect 1474 243 1503 249
rect 969 227 1447 241
rect 969 226 975 227
rect 946 220 975 226
rect 153 186 367 200
rect 153 184 159 186
rect 130 178 159 184
rect 137 114 151 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 353 73 367 186
rect 418 201 447 207
rect 418 184 424 201
rect 441 184 447 201
rect 418 178 447 184
rect 562 201 591 207
rect 562 184 568 201
rect 585 184 591 201
rect 562 178 591 184
rect 850 201 879 207
rect 850 184 856 201
rect 873 184 879 201
rect 850 178 879 184
rect 994 201 1023 207
rect 425 114 439 178
rect 569 147 583 178
rect 994 172 1000 201
rect 1017 172 1023 201
rect 1049 195 1063 227
rect 1433 207 1447 227
rect 1474 226 1480 243
rect 1497 226 1503 243
rect 1474 220 1503 226
rect 1138 201 1167 207
rect 994 166 1023 172
rect 1042 189 1071 195
rect 1042 172 1048 189
rect 1065 172 1071 189
rect 1138 184 1144 201
rect 1161 184 1167 201
rect 1138 178 1167 184
rect 1426 201 1455 207
rect 1426 184 1432 201
rect 1449 184 1455 201
rect 1426 178 1455 184
rect 1042 166 1071 172
rect 1145 147 1159 178
rect 569 133 1159 147
rect 569 114 583 133
rect 1145 114 1159 133
rect 1433 114 1447 178
rect 418 108 447 114
rect 418 91 424 108
rect 441 91 447 108
rect 418 85 447 91
rect 562 108 591 114
rect 562 91 568 108
rect 585 91 591 108
rect 994 108 1023 114
rect 994 106 1000 108
rect 562 85 591 91
rect 617 92 1000 106
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 346 67 375 73
rect 58 44 87 50
rect 178 49 207 55
rect 178 32 184 49
rect 201 32 207 49
rect 346 50 352 67
rect 369 50 375 67
rect 425 66 439 85
rect 617 66 631 92
rect 994 91 1000 92
rect 1017 91 1023 108
rect 994 85 1023 91
rect 1138 108 1167 114
rect 1138 91 1144 108
rect 1161 91 1167 108
rect 1138 85 1167 91
rect 1426 108 1455 114
rect 1426 91 1432 108
rect 1449 91 1455 108
rect 1426 85 1455 91
rect 1481 73 1495 220
rect 425 52 631 66
rect 946 67 975 73
rect 346 44 375 50
rect 946 50 952 67
rect 969 66 975 67
rect 1186 67 1215 73
rect 1186 66 1192 67
rect 969 52 1192 66
rect 969 50 975 52
rect 946 44 975 50
rect 1186 50 1192 52
rect 1209 50 1215 67
rect 1474 67 1503 73
rect 1186 44 1215 50
rect 1354 49 1383 55
rect 178 24 207 32
rect 610 27 639 33
rect 610 24 616 27
rect 0 10 616 24
rect 633 24 639 27
rect 778 27 807 33
rect 778 24 784 27
rect 633 10 784 24
rect 801 24 807 27
rect 1354 32 1360 49
rect 1377 32 1383 49
rect 1474 50 1480 67
rect 1497 50 1503 67
rect 1474 44 1503 50
rect 1354 24 1383 32
rect 801 10 1584 24
rect 0 -24 1584 10
<< labels >>
rlabel metal1 0 309 1584 357 0 VDD
port 1 se
rlabel metal1 0 -24 1584 24 0 GND
port 2 se
rlabel metal1 58 44 87 73 0 YC
port 3 se
rlabel metal1 65 73 79 220 0 YC
port 4 se
rlabel metal1 58 220 87 249 0 YC
port 5 se
rlabel metal1 1474 44 1503 73 0 YS
port 6 se
rlabel metal1 1481 73 1495 220 0 YS
port 7 se
rlabel metal1 1474 220 1503 249 0 YS
port 8 se
rlabel metal1 425 52 631 66 0 B
port 9 se
rlabel metal1 425 66 439 85 0 B
port 10 se
rlabel metal1 617 66 631 92 0 B
port 11 se
rlabel metal1 994 85 1023 92 0 B
port 12 se
rlabel metal1 617 92 1023 106 0 B
port 13 se
rlabel metal1 418 85 447 114 0 B
port 14 se
rlabel metal1 994 106 1023 114 0 B
port 15 se
rlabel metal1 425 114 439 178 0 B
port 16 se
rlabel metal1 418 178 447 207 0 B
port 17 se
rlabel metal1 562 85 591 114 0 A
port 18 se
rlabel metal1 1138 85 1167 114 0 A
port 19 se
rlabel metal1 569 114 583 133 0 A
port 20 se
rlabel metal1 1145 114 1159 133 0 A
port 21 se
rlabel metal1 569 133 1159 147 0 A
port 22 se
rlabel metal1 569 147 583 178 0 A
port 23 se
rlabel metal1 1145 147 1159 178 0 A
port 24 se
rlabel metal1 562 178 591 207 0 A
port 25 se
rlabel metal1 1138 178 1167 207 0 A
port 26 se
<< properties >>
string FIXED_BBOX 0 0 1584 333
<< end >>
