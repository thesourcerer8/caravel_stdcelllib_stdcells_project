VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 4.175 1.995 4.465 2.070 ;
        RECT 4.175 1.855 5.830 1.995 ;
        RECT 4.175 1.780 4.465 1.855 ;
        RECT 5.690 1.135 5.830 1.855 ;
        RECT 8.495 1.780 8.785 2.070 ;
        RECT 8.570 1.135 8.710 1.780 ;
        RECT 5.615 1.060 5.905 1.135 ;
        RECT 8.495 1.060 8.785 1.135 ;
        RECT 5.615 0.920 8.785 1.060 ;
        RECT 5.615 0.845 5.905 0.920 ;
        RECT 8.495 0.845 8.785 0.920 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.995 1.585 2.070 ;
        RECT 2.735 1.995 3.025 2.070 ;
        RECT 1.295 1.855 3.025 1.995 ;
        RECT 1.295 1.780 1.585 1.855 ;
        RECT 2.735 1.780 3.025 1.855 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 2.810 1.135 2.950 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
        RECT 2.735 0.845 3.025 1.135 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA 1.124200 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 7.535 0.440 7.825 0.730 ;
        RECT 1.850 0.240 1.990 0.440 ;
        RECT 7.610 0.240 7.750 0.440 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 7.535 2.735 7.825 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 2.167200 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.155 3.090 9.925 3.245 ;
        RECT 1.755 2.715 2.085 3.090 ;
        RECT 7.515 2.715 7.845 3.090 ;
      LAYER mcon ;
        RECT 7.595 3.245 7.765 3.415 ;
        RECT 7.595 2.795 7.765 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 4.655 0.440 4.945 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 10.080 3.330 ;
      LAYER li1 ;
        RECT 0.555 2.175 0.885 2.505 ;
        RECT 4.635 2.260 4.965 2.505 ;
        RECT 4.655 2.175 4.965 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 4.155 0.825 4.465 0.920 ;
        RECT 4.715 0.750 4.885 2.175 ;
        RECT 5.675 2.090 5.845 2.425 ;
        RECT 7.115 2.090 7.285 2.830 ;
        RECT 8.955 2.175 9.285 2.505 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 8.475 2.005 8.785 2.090 ;
        RECT 8.475 1.760 8.805 2.005 ;
        RECT 7.115 1.155 7.285 1.760 ;
        RECT 5.595 0.825 5.925 1.155 ;
        RECT 7.035 0.920 7.365 1.155 ;
        RECT 7.035 0.825 7.345 0.920 ;
        RECT 8.475 0.825 8.805 1.155 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.775 0.655 2.085 0.750 ;
        RECT 1.755 0.420 2.085 0.655 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 7.515 0.420 7.845 0.750 ;
        RECT 8.975 0.655 9.285 0.750 ;
        RECT 8.955 0.420 9.285 0.655 ;
        RECT 0.155 0.085 9.925 0.240 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 7.115 2.660 7.285 2.830 ;
        RECT 0.635 2.255 0.805 2.425 ;
        RECT 5.675 2.255 5.845 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 9.035 2.255 9.205 2.425 ;
        RECT 8.555 1.840 8.725 2.010 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 8.555 0.905 8.725 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 7.595 0.500 7.765 0.670 ;
        RECT 9.035 0.500 9.205 0.670 ;
        RECT 7.595 -0.085 7.765 0.085 ;
      LAYER met1 ;
        RECT 7.055 2.815 7.345 2.890 ;
        RECT 0.650 2.675 7.345 2.815 ;
        RECT 0.650 2.485 0.790 2.675 ;
        RECT 7.055 2.600 7.345 2.675 ;
        RECT 0.575 2.195 0.865 2.485 ;
        RECT 5.615 2.410 5.905 2.485 ;
        RECT 8.975 2.410 9.265 2.485 ;
        RECT 3.770 2.270 9.265 2.410 ;
        RECT 0.650 0.730 0.790 2.195 ;
        RECT 3.770 1.060 3.910 2.270 ;
        RECT 5.615 2.195 5.905 2.270 ;
        RECT 8.975 2.195 9.265 2.270 ;
        RECT 4.175 1.060 4.465 1.135 ;
        RECT 3.770 0.920 4.465 1.060 ;
        RECT 4.175 0.845 4.465 0.920 ;
        RECT 9.050 0.730 9.190 2.195 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 8.975 0.440 9.265 0.730 ;
  END
END XNOR2X1
END LIBRARY

