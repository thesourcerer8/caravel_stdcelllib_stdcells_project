magic
tech sky130A
timestamp 1624702806
<< nwell >>
rect 0 179 576 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 370 67 399 73
rect 370 66 376 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 51 281 66
rect 152 34 184 51
rect 201 34 281 51
rect 152 24 281 34
rect 296 50 376 66
rect 393 66 399 67
rect 393 50 425 66
rect 296 24 425 50
rect 440 51 519 66
rect 440 34 472 51
rect 489 34 519 51
rect 440 24 519 34
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 299 281 309
rect 152 282 184 299
rect 201 282 281 299
rect 152 225 281 282
rect 296 243 425 309
rect 296 226 376 243
rect 393 226 425 243
rect 296 225 425 226
rect 440 299 519 309
rect 440 282 472 299
rect 489 282 519 299
rect 440 225 519 282
rect 58 220 87 225
rect 370 220 399 225
<< ndiffc >>
rect 64 50 81 67
rect 184 34 201 51
rect 376 50 393 67
rect 472 34 489 51
<< pdiffc >>
rect 64 226 81 243
rect 184 282 201 299
rect 376 226 393 243
rect 472 282 489 299
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
<< locali >>
rect 0 342 576 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 576 342
rect 0 309 576 325
rect 176 299 209 309
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 464 299 497 309
rect 464 282 472 299
rect 489 282 497 299
rect 464 274 497 282
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 368 243 401 251
rect 368 226 376 243
rect 393 226 401 243
rect 368 218 401 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 418 201 449 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 136 116 153 131
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 416 108 449 116
rect 416 92 424 108
rect 272 83 305 91
rect 418 91 424 92
rect 441 91 449 108
rect 418 83 449 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 368 67 401 75
rect 56 42 89 50
rect 176 51 209 59
rect 176 34 184 51
rect 201 34 209 51
rect 368 50 376 67
rect 393 50 401 67
rect 368 42 401 50
rect 464 51 497 59
rect 176 24 209 34
rect 464 34 472 51
rect 489 34 497 51
rect 464 24 497 34
rect 0 9 576 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 576 9
rect 0 -24 576 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 304 325 321 342
rect 352 325 369 342
rect 400 325 417 342
rect 448 325 465 342
rect 496 325 513 342
rect 544 325 561 342
rect 184 282 201 299
rect 472 282 489 299
rect 64 226 81 243
rect 376 226 393 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 136 131 153 148
rect 280 91 297 108
rect 424 91 441 108
rect 64 50 81 67
rect 184 34 201 51
rect 376 50 393 67
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
rect 304 -9 321 9
rect 352 -9 369 9
rect 400 -9 417 9
rect 448 -9 465 9
rect 496 -9 513 9
rect 544 -9 561 9
<< metal1 >>
rect 0 342 576 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 576 342
rect 0 309 576 325
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 466 299 495 309
rect 466 282 472 299
rect 489 282 495 299
rect 466 276 495 282
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 58 220 87 226
rect 370 243 399 249
rect 370 226 376 243
rect 393 241 399 243
rect 393 227 487 241
rect 393 226 399 227
rect 370 220 399 226
rect 65 106 79 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 418 201 447 207
rect 418 184 424 201
rect 441 184 447 201
rect 418 178 447 184
rect 137 154 151 178
rect 130 148 159 154
rect 130 131 136 148
rect 153 131 159 148
rect 130 125 159 131
rect 281 114 295 178
rect 425 114 439 178
rect 274 108 303 114
rect 274 106 280 108
rect 65 92 280 106
rect 65 73 79 92
rect 274 91 280 92
rect 297 106 303 108
rect 418 108 447 114
rect 418 106 424 108
rect 297 92 424 106
rect 297 91 303 92
rect 274 85 303 91
rect 418 91 424 92
rect 441 91 447 108
rect 418 85 447 91
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 370 67 399 73
rect 58 44 87 50
rect 178 51 207 57
rect 178 34 184 51
rect 201 34 207 51
rect 370 50 376 67
rect 393 66 399 67
rect 473 66 487 227
rect 393 52 487 66
rect 393 50 399 52
rect 370 44 399 50
rect 178 24 207 34
rect 0 9 576 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 576 9
rect 0 -24 576 -9
<< labels >>
rlabel locali 0 309 576 357 0 VDD
port 1 se
rlabel metal1 0 309 576 357 0 VDD
port 2 se
rlabel locali 0 -24 576 24 0 GND
port 3 se
rlabel metal1 0 -24 576 24 0 GND
port 4 se
rlabel metal1 370 44 399 52 0 Y
port 5 se
rlabel metal1 370 52 487 66 0 Y
port 6 se
rlabel metal1 370 66 399 73 0 Y
port 7 se
rlabel metal1 370 220 399 227 0 Y
port 8 se
rlabel metal1 473 66 487 227 0 Y
port 9 se
rlabel metal1 370 227 487 241 0 Y
port 10 se
rlabel metal1 370 241 399 249 0 Y
port 11 se
rlabel metal1 130 125 159 154 0 A
port 12 se
rlabel metal1 137 154 151 178 0 A
port 13 se
rlabel metal1 130 178 159 207 0 A
port 14 se
<< properties >>
string FIXED_BBOX 0 0 576 333
<< end >>
