magic
tech sky130A
timestamp 1623602813
<< nwell >>
rect 0 179 576 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
<< ndiff >>
rect 82 66 111 69
rect 466 66 495 69
rect 58 63 137 66
rect 58 46 88 63
rect 105 46 137 63
rect 58 24 137 46
rect 152 24 281 66
rect 296 36 425 66
rect 296 24 328 36
rect 322 19 328 24
rect 345 24 425 36
rect 440 63 519 66
rect 440 46 472 63
rect 489 46 519 63
rect 440 24 519 46
rect 345 19 351 24
rect 322 13 351 19
<< pdiff >>
rect 58 309 87 312
rect 322 309 351 312
rect 58 306 137 309
rect 58 289 64 306
rect 81 289 137 306
rect 58 225 137 289
rect 152 238 281 309
rect 152 225 184 238
rect 178 221 184 225
rect 201 225 281 238
rect 296 306 425 309
rect 296 289 328 306
rect 345 289 425 306
rect 296 225 425 289
rect 440 238 519 309
rect 440 225 472 238
rect 201 221 207 225
rect 178 215 207 221
rect 466 221 472 225
rect 489 225 519 238
rect 489 221 495 225
rect 466 215 495 221
<< ndiffc >>
rect 88 46 105 63
rect 328 19 345 36
rect 472 46 489 63
<< pdiffc >>
rect 64 289 81 306
rect 184 221 201 238
rect 328 289 345 306
rect 472 221 489 238
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 425 309 440 330
rect 137 206 152 225
rect 281 206 296 225
rect 425 206 440 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 137 66 152 78
rect 281 66 296 78
rect 425 66 440 78
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
<< locali >>
rect 56 306 89 314
rect 56 289 64 306
rect 81 289 89 306
rect 56 281 89 289
rect 320 306 353 314
rect 320 289 328 306
rect 345 289 353 306
rect 320 281 353 289
rect 176 238 209 246
rect 176 223 184 238
rect 178 221 184 223
rect 201 221 209 238
rect 464 238 497 246
rect 464 223 472 238
rect 178 213 209 221
rect 466 221 472 223
rect 489 221 497 238
rect 466 213 497 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 128 103 161 111
rect 128 88 136 103
rect 130 86 136 88
rect 153 86 161 103
rect 130 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 80 63 113 71
rect 80 46 88 63
rect 105 46 113 63
rect 466 63 497 71
rect 466 61 472 63
rect 80 38 113 46
rect 464 46 472 61
rect 489 46 497 63
rect 320 36 353 44
rect 464 38 497 46
rect 320 19 328 36
rect 345 19 353 36
rect 320 11 353 19
<< viali >>
rect 64 289 81 306
rect 328 289 345 306
rect 184 221 201 238
rect 472 221 489 238
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 88 46 105 63
rect 472 46 489 63
rect 328 19 345 36
<< metal1 >>
rect 0 309 576 357
rect 58 306 87 309
rect 58 289 64 306
rect 81 289 87 306
rect 58 283 87 289
rect 322 306 351 309
rect 322 289 328 306
rect 345 289 351 306
rect 322 283 351 289
rect 178 238 207 244
rect 178 237 184 238
rect 89 223 184 237
rect 89 69 103 223
rect 178 221 184 223
rect 201 237 207 238
rect 466 238 495 244
rect 201 223 439 237
rect 201 221 207 223
rect 178 215 207 221
rect 425 204 439 223
rect 466 221 472 238
rect 489 221 495 238
rect 466 215 495 221
rect 130 198 159 204
rect 130 181 136 198
rect 153 181 159 198
rect 130 175 159 181
rect 274 198 303 204
rect 274 181 280 198
rect 297 181 303 198
rect 274 175 303 181
rect 418 198 447 204
rect 418 181 424 198
rect 441 181 447 198
rect 418 175 447 181
rect 137 109 151 175
rect 281 109 295 175
rect 425 109 439 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 86 159 103
rect 130 80 159 86
rect 274 103 303 109
rect 274 86 280 103
rect 297 86 303 103
rect 274 80 303 86
rect 418 103 447 109
rect 418 86 424 103
rect 441 86 447 103
rect 418 80 447 86
rect 473 69 487 215
rect 82 63 111 69
rect 82 46 88 63
rect 105 46 111 63
rect 82 40 111 46
rect 466 63 495 69
rect 466 46 472 63
rect 489 46 495 63
rect 322 36 351 42
rect 466 40 495 46
rect 322 24 328 36
rect 0 19 328 24
rect 345 24 351 36
rect 345 19 576 24
rect 0 -24 576 19
<< labels >>
rlabel metal1 0 309 576 357 0 VDD
port 1 se
rlabel metal1 0 -24 576 24 0 GND
port 2 se
rlabel metal1 466 40 495 69 0 Y
port 3 se
rlabel metal1 473 69 487 215 0 Y
port 4 se
rlabel metal1 466 215 495 244 0 Y
port 5 se
rlabel metal1 130 80 159 109 0 A
port 6 se
rlabel metal1 137 109 151 175 0 A
port 7 se
rlabel metal1 130 175 159 204 0 A
port 8 se
rlabel metal1 274 80 303 109 0 B
port 9 se
rlabel metal1 281 109 295 175 0 B
port 10 se
rlabel metal1 274 175 303 204 0 B
port 11 se
<< properties >>
string FIXED_BBOX 0 0 576 333
<< end >>
