VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BUFX4
  CLASS CORE ;
  FOREIGN BUFX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 0.914200 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 4.655 0.440 4.945 0.730 ;
        RECT 1.850 0.240 1.990 0.440 ;
        RECT 4.730 0.240 4.870 0.440 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 1.775 2.735 2.065 3.090 ;
        RECT 4.655 2.735 4.945 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.155 3.215 5.605 3.245 ;
        RECT 0.155 3.090 4.465 3.215 ;
        RECT 5.135 3.090 5.605 3.215 ;
        RECT 1.755 2.715 2.085 3.090 ;
      LAYER mcon ;
        RECT 4.715 3.245 4.885 3.415 ;
        RECT 1.835 2.795 2.005 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 3.215 0.440 3.505 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 5.760 3.330 ;
      LAYER li1 ;
        RECT 4.635 2.715 4.965 3.045 ;
        RECT 0.555 2.175 0.885 2.505 ;
        RECT 3.195 2.175 3.525 2.505 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 2.005 3.025 2.090 ;
        RECT 2.715 1.760 3.045 2.005 ;
        RECT 1.355 1.155 1.525 1.760 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 3.275 0.750 3.445 2.175 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 4.155 0.825 4.465 0.920 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.215 0.655 3.525 0.750 ;
        RECT 3.195 0.420 3.525 0.655 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 0.155 0.085 5.605 0.240 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 4.715 2.795 4.885 2.965 ;
        RECT 0.635 2.255 0.805 2.425 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 4.715 -0.085 4.885 0.085 ;
      LAYER met1 ;
        RECT 0.575 2.195 0.865 2.485 ;
        RECT 0.650 1.995 0.790 2.195 ;
        RECT 2.735 1.995 3.025 2.070 ;
        RECT 4.175 1.995 4.465 2.070 ;
        RECT 0.650 1.855 4.465 1.995 ;
        RECT 0.650 0.730 0.790 1.855 ;
        RECT 2.735 1.780 3.025 1.855 ;
        RECT 4.175 1.780 4.465 1.855 ;
        RECT 2.810 1.135 2.950 1.780 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 2.735 0.845 3.025 1.135 ;
        RECT 4.175 0.845 4.465 1.135 ;
        RECT 0.575 0.440 0.865 0.730 ;
  END
END BUFX4
END LIBRARY

