magic
tech sky130A
timestamp 1621277891
<< end >>
