VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF2
  CLASS CORE ;
  FOREIGN CLKBUF2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.370 2.675 2.950 2.815 ;
        RECT 1.370 2.070 1.510 2.675 ;
        RECT 2.810 2.070 2.950 2.675 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 2.735 1.780 3.025 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 3.514700 ;
    PORT
      LAYER met1 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 3.215 0.440 3.505 0.730 ;
        RECT 6.095 0.440 6.385 0.730 ;
        RECT 8.975 0.440 9.265 0.730 ;
        RECT 11.855 0.440 12.145 0.730 ;
        RECT 14.735 0.440 15.025 0.730 ;
        RECT 17.615 0.440 17.905 0.730 ;
        RECT 0.650 0.240 0.790 0.440 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 6.170 0.240 6.310 0.440 ;
        RECT 9.050 0.240 9.190 0.440 ;
        RECT 11.930 0.240 12.070 0.440 ;
        RECT 14.810 0.240 14.950 0.440 ;
        RECT 17.690 0.240 17.830 0.440 ;
        RECT 0.000 -0.240 18.720 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 18.720 3.570 ;
        RECT 0.575 2.735 0.865 3.090 ;
        RECT 3.215 2.735 3.505 3.090 ;
        RECT 6.095 2.735 6.385 3.090 ;
        RECT 8.975 2.735 9.265 3.090 ;
        RECT 11.855 2.735 12.145 3.090 ;
        RECT 14.735 2.735 15.025 3.090 ;
        RECT 17.615 2.735 17.905 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 5.661600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 18.720 3.415 ;
        RECT 0.155 3.215 18.565 3.245 ;
        RECT 0.155 3.090 3.025 3.215 ;
        RECT 3.695 3.090 18.565 3.215 ;
        RECT 0.555 2.715 0.885 3.090 ;
        RECT 6.075 2.715 6.405 3.090 ;
        RECT 8.955 2.715 9.285 3.090 ;
        RECT 11.835 2.715 12.165 3.090 ;
        RECT 14.715 2.715 15.045 3.090 ;
        RECT 17.595 2.715 17.925 3.090 ;
      LAYER mcon ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 16.475 3.245 16.645 3.415 ;
        RECT 16.955 3.245 17.125 3.415 ;
        RECT 17.435 3.245 17.605 3.415 ;
        RECT 17.915 3.245 18.085 3.415 ;
        RECT 0.635 2.795 0.805 2.965 ;
        RECT 6.155 2.795 6.325 2.965 ;
        RECT 9.035 2.795 9.205 2.965 ;
        RECT 11.915 2.795 12.085 2.965 ;
        RECT 14.795 2.795 14.965 2.965 ;
        RECT 17.675 2.795 17.845 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 16.175 0.440 16.465 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 18.720 3.330 ;
      LAYER li1 ;
        RECT 3.195 2.715 3.525 3.045 ;
        RECT 1.755 2.260 2.085 2.505 ;
        RECT 1.775 2.175 2.085 2.260 ;
        RECT 4.635 2.175 4.965 2.505 ;
        RECT 5.675 2.090 5.845 2.830 ;
        RECT 7.515 2.260 7.845 2.505 ;
        RECT 7.535 2.175 7.845 2.260 ;
        RECT 8.555 2.090 8.725 2.830 ;
        RECT 10.395 2.260 10.725 2.505 ;
        RECT 10.415 2.175 10.725 2.260 ;
        RECT 11.435 2.090 11.605 2.830 ;
        RECT 13.275 2.260 13.605 2.505 ;
        RECT 13.295 2.175 13.605 2.260 ;
        RECT 14.315 2.090 14.485 2.830 ;
        RECT 16.155 2.175 16.485 2.505 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 2.005 4.465 2.090 ;
        RECT 4.155 1.760 4.485 2.005 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 9.915 1.760 10.245 2.090 ;
        RECT 11.355 1.760 11.685 2.090 ;
        RECT 12.795 1.760 13.125 2.090 ;
        RECT 14.235 1.760 14.565 2.090 ;
        RECT 15.675 2.005 15.985 2.090 ;
        RECT 15.675 1.760 16.005 2.005 ;
        RECT 2.795 1.155 2.965 1.760 ;
        RECT 5.675 1.445 5.845 1.760 ;
        RECT 8.555 1.445 8.725 1.760 ;
        RECT 11.435 1.445 11.605 1.760 ;
        RECT 14.315 1.445 14.485 1.760 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 4.155 0.825 4.465 0.920 ;
        RECT 5.595 0.825 5.925 1.155 ;
        RECT 7.035 0.920 7.365 1.155 ;
        RECT 8.475 0.920 8.805 1.155 ;
        RECT 9.915 0.920 10.245 1.155 ;
        RECT 7.035 0.825 7.345 0.920 ;
        RECT 8.475 0.825 8.785 0.920 ;
        RECT 9.915 0.825 10.225 0.920 ;
        RECT 11.355 0.825 11.685 1.155 ;
        RECT 12.795 0.920 13.125 1.155 ;
        RECT 14.235 0.920 14.565 1.155 ;
        RECT 15.675 0.920 16.005 1.155 ;
        RECT 12.795 0.825 13.105 0.920 ;
        RECT 14.235 0.825 14.545 0.920 ;
        RECT 15.675 0.825 15.985 0.920 ;
        RECT 16.235 0.750 16.405 2.175 ;
        RECT 17.115 1.760 17.445 2.090 ;
        RECT 17.115 0.825 17.445 1.155 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.215 0.655 3.525 0.750 ;
        RECT 3.195 0.420 3.525 0.655 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 6.095 0.655 6.405 0.750 ;
        RECT 6.075 0.420 6.405 0.655 ;
        RECT 7.515 0.420 7.845 0.750 ;
        RECT 8.955 0.420 9.285 0.750 ;
        RECT 10.395 0.420 10.725 0.750 ;
        RECT 11.855 0.655 12.165 0.750 ;
        RECT 11.835 0.420 12.165 0.655 ;
        RECT 13.275 0.420 13.605 0.750 ;
        RECT 14.715 0.420 15.045 0.750 ;
        RECT 16.155 0.420 16.485 0.750 ;
        RECT 17.615 0.655 17.925 0.750 ;
        RECT 17.595 0.420 17.925 0.655 ;
        RECT 0.155 0.085 18.565 0.240 ;
        RECT 0.000 -0.085 18.720 0.085 ;
      LAYER mcon ;
        RECT 3.275 2.795 3.445 2.965 ;
        RECT 5.675 2.660 5.845 2.830 ;
        RECT 1.835 2.255 2.005 2.425 ;
        RECT 4.715 2.255 4.885 2.425 ;
        RECT 8.555 2.660 8.725 2.830 ;
        RECT 7.595 2.255 7.765 2.425 ;
        RECT 11.435 2.660 11.605 2.830 ;
        RECT 10.475 2.255 10.645 2.425 ;
        RECT 14.315 2.660 14.485 2.830 ;
        RECT 13.355 2.255 13.525 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 7.115 1.840 7.285 2.010 ;
        RECT 9.995 1.840 10.165 2.010 ;
        RECT 12.875 1.840 13.045 2.010 ;
        RECT 15.755 1.840 15.925 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 7.115 0.905 7.285 1.075 ;
        RECT 8.555 0.905 8.725 1.075 ;
        RECT 9.995 0.905 10.165 1.075 ;
        RECT 11.435 0.905 11.605 1.075 ;
        RECT 12.875 0.905 13.045 1.075 ;
        RECT 14.315 0.905 14.485 1.075 ;
        RECT 15.755 0.905 15.925 1.075 ;
        RECT 17.195 1.840 17.365 2.010 ;
        RECT 17.195 0.905 17.365 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 6.155 0.500 6.325 0.670 ;
        RECT 7.595 0.500 7.765 0.670 ;
        RECT 9.035 0.500 9.205 0.670 ;
        RECT 10.475 0.500 10.645 0.670 ;
        RECT 11.915 0.500 12.085 0.670 ;
        RECT 13.355 0.500 13.525 0.670 ;
        RECT 14.795 0.500 14.965 0.670 ;
        RECT 16.235 0.500 16.405 0.670 ;
        RECT 17.675 0.500 17.845 0.670 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
        RECT 16.955 -0.085 17.125 0.085 ;
        RECT 17.435 -0.085 17.605 0.085 ;
        RECT 17.915 -0.085 18.085 0.085 ;
      LAYER met1 ;
        RECT 5.615 2.815 5.905 2.890 ;
        RECT 8.495 2.815 8.785 2.890 ;
        RECT 11.375 2.815 11.665 2.890 ;
        RECT 14.255 2.815 14.545 2.890 ;
        RECT 4.250 2.675 5.905 2.815 ;
        RECT 1.775 2.195 2.065 2.485 ;
        RECT 1.850 1.060 1.990 2.195 ;
        RECT 4.250 2.070 4.390 2.675 ;
        RECT 5.615 2.600 5.905 2.675 ;
        RECT 7.130 2.675 8.785 2.815 ;
        RECT 4.655 2.195 4.945 2.485 ;
        RECT 4.175 1.780 4.465 2.070 ;
        RECT 4.730 1.995 4.870 2.195 ;
        RECT 7.130 2.070 7.270 2.675 ;
        RECT 8.495 2.600 8.785 2.675 ;
        RECT 10.010 2.675 11.665 2.815 ;
        RECT 7.535 2.195 7.825 2.485 ;
        RECT 7.055 1.995 7.345 2.070 ;
        RECT 4.730 1.855 7.345 1.995 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 4.175 1.060 4.465 1.135 ;
        RECT 1.850 0.920 4.465 1.060 ;
        RECT 1.850 0.730 1.990 0.920 ;
        RECT 4.175 0.845 4.465 0.920 ;
        RECT 4.730 0.730 4.870 1.855 ;
        RECT 7.055 1.780 7.345 1.855 ;
        RECT 7.610 1.995 7.750 2.195 ;
        RECT 10.010 2.070 10.150 2.675 ;
        RECT 11.375 2.600 11.665 2.675 ;
        RECT 12.890 2.675 14.545 2.815 ;
        RECT 10.415 2.195 10.705 2.485 ;
        RECT 9.935 1.995 10.225 2.070 ;
        RECT 7.610 1.855 10.225 1.995 ;
        RECT 5.615 1.385 5.905 1.675 ;
        RECT 5.690 1.135 5.830 1.385 ;
        RECT 7.130 1.135 7.270 1.780 ;
        RECT 5.615 0.845 5.905 1.135 ;
        RECT 7.055 0.845 7.345 1.135 ;
        RECT 7.610 0.730 7.750 1.855 ;
        RECT 9.935 1.780 10.225 1.855 ;
        RECT 10.490 1.995 10.630 2.195 ;
        RECT 12.890 2.070 13.030 2.675 ;
        RECT 14.255 2.600 14.545 2.675 ;
        RECT 13.295 2.195 13.585 2.485 ;
        RECT 12.815 1.995 13.105 2.070 ;
        RECT 10.490 1.855 13.105 1.995 ;
        RECT 8.495 1.385 8.785 1.675 ;
        RECT 8.570 1.135 8.710 1.385 ;
        RECT 10.010 1.135 10.150 1.780 ;
        RECT 8.495 0.845 8.785 1.135 ;
        RECT 9.935 0.845 10.225 1.135 ;
        RECT 10.490 0.730 10.630 1.855 ;
        RECT 12.815 1.780 13.105 1.855 ;
        RECT 13.370 1.995 13.510 2.195 ;
        RECT 15.695 1.995 15.985 2.070 ;
        RECT 17.135 1.995 17.425 2.070 ;
        RECT 13.370 1.855 17.425 1.995 ;
        RECT 11.375 1.385 11.665 1.675 ;
        RECT 11.450 1.135 11.590 1.385 ;
        RECT 12.890 1.135 13.030 1.780 ;
        RECT 11.375 0.845 11.665 1.135 ;
        RECT 12.815 0.845 13.105 1.135 ;
        RECT 13.370 0.730 13.510 1.855 ;
        RECT 15.695 1.780 15.985 1.855 ;
        RECT 17.135 1.780 17.425 1.855 ;
        RECT 14.255 1.385 14.545 1.675 ;
        RECT 14.330 1.135 14.470 1.385 ;
        RECT 15.770 1.135 15.910 1.780 ;
        RECT 17.210 1.135 17.350 1.780 ;
        RECT 14.255 0.845 14.545 1.135 ;
        RECT 15.695 0.845 15.985 1.135 ;
        RECT 17.135 0.845 17.425 1.135 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 4.655 0.440 4.945 0.730 ;
        RECT 7.535 0.440 7.825 0.730 ;
        RECT 10.415 0.440 10.705 0.730 ;
        RECT 13.295 0.440 13.585 0.730 ;
  END
END CLKBUF2
END LIBRARY

