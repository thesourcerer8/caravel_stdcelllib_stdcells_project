`default_nettype none

/*
 *-------------------------------------------------------------
 *
 * user_proj_cells  (LibreSilicon Testwafer #1)
 *
 */

module AND2X1(
  inout B, // input
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module AND2X2(
  inout B, // input
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module AOI21X1(
  inout C, // input
  inout B, // input
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module AOI22X1(
  inout D, // input
  inout C, // input
  inout B, // input
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module BUFX2(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module BUFX4(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module CLKBUF1(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module HAX1(
  inout B, // input
  inout A, // input
  inout YS, // output
  inout YC, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module INV(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module INVX1(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module INVX2(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module INVX4(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

module INVX8(
  inout A, // input
  inout Y, // output
	inout vdd, // cell power supply
	inout gnd  // cell ground supply
);
endmodule

