VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 1.780 3.025 2.070 ;
        RECT 2.810 1.135 2.950 1.780 ;
        RECT 2.735 0.845 3.025 1.135 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA 0.562100 ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 0.575 2.735 0.865 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 0.663600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.155 3.090 4.165 3.245 ;
        RECT 0.555 2.715 0.885 3.090 ;
      LAYER mcon ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 0.635 2.795 0.805 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.383750 ;
    PORT
      LAYER met1 ;
        RECT 3.215 2.195 3.505 2.485 ;
        RECT 3.290 0.730 3.430 2.195 ;
        RECT 0.815 0.655 1.105 0.730 ;
        RECT 3.215 0.655 3.505 0.730 ;
        RECT 0.815 0.515 3.505 0.655 ;
        RECT 0.815 0.440 1.105 0.515 ;
        RECT 3.215 0.440 3.505 0.515 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 4.320 3.330 ;
      LAYER li1 ;
        RECT 3.195 2.260 3.525 2.505 ;
        RECT 3.215 2.175 3.525 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 2.715 0.920 3.045 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 2.715 0.825 3.025 0.920 ;
        RECT 0.795 0.655 1.105 0.750 ;
        RECT 0.795 0.420 1.125 0.655 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.195 0.420 3.525 0.750 ;
        RECT 1.835 0.240 2.005 0.420 ;
        RECT 0.155 0.085 4.165 0.240 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 3.275 2.255 3.445 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 0.875 0.500 1.045 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 1.835 -0.085 2.005 0.085 ;
  END
END NOR2X1
END LIBRARY

