MACRO XOR2X1
 CLASS CORE ;
 FOREIGN XOR2X1 0 0 ;
 SIZE 10.08 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 3.09000000 10.08000000 3.57000000 ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 10.08000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 -0.24000000 10.08000000 0.24000000 ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 10.08000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 5.13500000 0.44000000 5.42500000 0.51500000 ;
        RECT 6.09500000 0.44000000 6.38500000 0.51500000 ;
        RECT 5.13500000 0.51500000 6.38500000 0.65500000 ;
        RECT 5.13500000 0.65500000 5.42500000 0.73000000 ;
        RECT 6.09500000 0.65500000 6.38500000 0.73000000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 8.49500000 0.84500000 8.78500000 1.13500000 ;
        RECT 2.73500000 1.25000000 3.02500000 1.32500000 ;
        RECT 8.57000000 1.13500000 8.71000000 1.32500000 ;
        RECT 2.73500000 1.32500000 8.71000000 1.46500000 ;
        RECT 2.73500000 1.46500000 3.02500000 1.54000000 ;
        RECT 8.57000000 1.46500000 8.71000000 1.78000000 ;
        RECT 8.49500000 1.78000000 8.78500000 2.07000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 4.17500000 0.44000000 4.46500000 0.51500000 ;
        RECT 2.09000000 0.51500000 4.46500000 0.65500000 ;
        RECT 4.17500000 0.65500000 4.46500000 0.73000000 ;
        RECT 2.09000000 0.65500000 2.23000000 0.78500000 ;
        RECT 1.37000000 0.78500000 2.23000000 0.84500000 ;
        RECT 1.29500000 0.84500000 2.23000000 0.92500000 ;
        RECT 1.29500000 0.92500000 1.58500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.38500000 ;
        RECT 1.29500000 1.38500000 1.58500000 1.67500000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 5.67500000 0.90500000 5.84500000 1.07500000 ;
     RECT 7.11500000 0.90500000 7.28500000 1.07500000 ;
     RECT 8.55500000 0.90500000 8.72500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;
     RECT 7.11500000 1.84000000 7.28500000 2.01000000 ;
     RECT 8.55500000 1.84000000 8.72500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 9.03500000 2.25500000 9.20500000 2.42500000 ;
     RECT 5.19500000 2.79500000 5.36500000 2.96500000 ;
     RECT 1.83500000 2.82000000 2.00500000 2.99000000 ;
     RECT 7.59500000 2.82000000 7.76500000 2.99000000 ;

    LAYER ndiffc ;
     RECT 1.83500000 0.34000000 2.00500000 0.51000000 ;
     RECT 7.59500000 0.34000000 7.76500000 0.51000000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 5.19500000 0.50000000 5.36500000 0.67000000 ;
     RECT 9.03500000 0.50000000 9.20500000 0.67000000 ;

    LAYER li1 ;
     RECT 1.75500000 0.26000000 2.08500000 0.59000000 ;
     RECT 0.00000000 -0.24000000 10.08000000 0.24000000 ;
     RECT 7.51500000 0.24000000 7.84500000 0.59000000 ;
     RECT 0.55500000 0.42000000 0.88500000 0.75000000 ;
     RECT 5.11500000 0.42000000 5.44500000 0.75000000 ;
     RECT 8.95500000 0.42000000 9.28500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 4.23500000 0.50000000 4.40500000 0.82500000 ;
     RECT 4.15500000 0.82500000 4.48500000 1.15500000 ;
     RECT 5.59500000 0.82500000 5.92500000 1.15500000 ;
     RECT 7.03500000 0.82500000 7.36500000 1.15500000 ;
     RECT 8.47500000 0.82500000 8.80500000 1.15500000 ;
     RECT 6.15500000 0.50000000 6.32500000 1.88500000 ;
     RECT 2.71500000 0.82500000 3.04500000 1.15500000 ;
     RECT 2.79500000 1.15500000 2.96500000 1.76000000 ;
     RECT 2.71500000 1.76000000 3.04500000 2.09000000 ;
     RECT 4.15500000 1.76000000 4.48500000 2.09000000 ;
     RECT 5.59500000 1.76000000 5.92500000 2.09000000 ;
     RECT 7.03500000 1.76000000 7.36500000 2.09000000 ;
     RECT 8.47500000 1.76000000 8.80500000 2.09000000 ;
     RECT 1.35500000 1.44500000 1.52500000 1.76000000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 1.35500000 2.09000000 1.52500000 2.42500000 ;
     RECT 0.55500000 2.17500000 0.88500000 2.50500000 ;
     RECT 8.95500000 2.17500000 9.28500000 2.50500000 ;
     RECT 5.11500000 2.71500000 5.44500000 3.04500000 ;
     RECT 1.75500000 2.74000000 2.08500000 3.07000000 ;
     RECT 7.51500000 2.74000000 7.84500000 3.07000000 ;
     RECT 0.00000000 3.09000000 10.08000000 3.57000000 ;

    LAYER viali ;
     RECT 0.15500000 -0.08500000 0.32500000 0.08500000 ;
     RECT 0.63500000 -0.08500000 0.80500000 0.08500000 ;
     RECT 1.11500000 -0.08500000 1.28500000 0.08500000 ;
     RECT 1.59500000 -0.08500000 1.76500000 0.08500000 ;
     RECT 2.07500000 -0.08500000 2.24500000 0.08500000 ;
     RECT 2.55500000 -0.08500000 2.72500000 0.08500000 ;
     RECT 3.03500000 -0.08500000 3.20500000 0.08500000 ;
     RECT 3.51500000 -0.08500000 3.68500000 0.08500000 ;
     RECT 3.99500000 -0.08500000 4.16500000 0.08500000 ;
     RECT 4.47500000 -0.08500000 4.64500000 0.08500000 ;
     RECT 4.95500000 -0.08500000 5.12500000 0.08500000 ;
     RECT 5.43500000 -0.08500000 5.60500000 0.08500000 ;
     RECT 5.91500000 -0.08500000 6.08500000 0.08500000 ;
     RECT 6.39500000 -0.08500000 6.56500000 0.08500000 ;
     RECT 6.87500000 -0.08500000 7.04500000 0.08500000 ;
     RECT 7.35500000 -0.08500000 7.52500000 0.08500000 ;
     RECT 7.83500000 -0.08500000 8.00500000 0.08500000 ;
     RECT 8.31500000 -0.08500000 8.48500000 0.08500000 ;
     RECT 8.79500000 -0.08500000 8.96500000 0.08500000 ;
     RECT 9.27500000 -0.08500000 9.44500000 0.08500000 ;
     RECT 9.75500000 -0.08500000 9.92500000 0.08500000 ;
     RECT 1.83500000 0.34000000 2.00500000 0.51000000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 4.23500000 0.50000000 4.40500000 0.67000000 ;
     RECT 5.19500000 0.50000000 5.36500000 0.67000000 ;
     RECT 6.15500000 0.50000000 6.32500000 0.67000000 ;
     RECT 9.03500000 0.50000000 9.20500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 5.67500000 0.90500000 5.84500000 1.07500000 ;
     RECT 7.11500000 0.90500000 7.28500000 1.07500000 ;
     RECT 8.55500000 0.90500000 8.72500000 1.07500000 ;
     RECT 2.79500000 1.31000000 2.96500000 1.48000000 ;
     RECT 1.35500000 1.44500000 1.52500000 1.61500000 ;
     RECT 6.15500000 1.71500000 6.32500000 1.88500000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;
     RECT 7.11500000 1.84000000 7.28500000 2.01000000 ;
     RECT 8.55500000 1.84000000 8.72500000 2.01000000 ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 1.35500000 2.25500000 1.52500000 2.42500000 ;
     RECT 9.03500000 2.25500000 9.20500000 2.42500000 ;
     RECT 5.19500000 2.79500000 5.36500000 2.96500000 ;
     RECT 1.83500000 2.82000000 2.00500000 2.99000000 ;
     RECT 7.59500000 2.82000000 7.76500000 2.99000000 ;
     RECT 0.15500000 3.24500000 0.32500000 3.41500000 ;
     RECT 0.63500000 3.24500000 0.80500000 3.41500000 ;
     RECT 1.11500000 3.24500000 1.28500000 3.41500000 ;
     RECT 1.59500000 3.24500000 1.76500000 3.41500000 ;
     RECT 2.07500000 3.24500000 2.24500000 3.41500000 ;
     RECT 2.55500000 3.24500000 2.72500000 3.41500000 ;
     RECT 3.03500000 3.24500000 3.20500000 3.41500000 ;
     RECT 3.51500000 3.24500000 3.68500000 3.41500000 ;
     RECT 3.99500000 3.24500000 4.16500000 3.41500000 ;
     RECT 4.47500000 3.24500000 4.64500000 3.41500000 ;
     RECT 4.95500000 3.24500000 5.12500000 3.41500000 ;
     RECT 5.43500000 3.24500000 5.60500000 3.41500000 ;
     RECT 5.91500000 3.24500000 6.08500000 3.41500000 ;
     RECT 6.39500000 3.24500000 6.56500000 3.41500000 ;
     RECT 6.87500000 3.24500000 7.04500000 3.41500000 ;
     RECT 7.35500000 3.24500000 7.52500000 3.41500000 ;
     RECT 7.83500000 3.24500000 8.00500000 3.41500000 ;
     RECT 8.31500000 3.24500000 8.48500000 3.41500000 ;
     RECT 8.79500000 3.24500000 8.96500000 3.41500000 ;
     RECT 9.27500000 3.24500000 9.44500000 3.41500000 ;
     RECT 9.75500000 3.24500000 9.92500000 3.41500000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 10.08000000 0.24000000 ;
     RECT 1.77500000 0.24000000 2.06500000 0.57000000 ;
     RECT 5.13500000 0.44000000 5.42500000 0.51500000 ;
     RECT 6.09500000 0.44000000 6.38500000 0.51500000 ;
     RECT 5.13500000 0.51500000 6.38500000 0.65500000 ;
     RECT 5.13500000 0.65500000 5.42500000 0.73000000 ;
     RECT 6.09500000 0.65500000 6.38500000 0.73000000 ;
     RECT 4.17500000 0.44000000 4.46500000 0.51500000 ;
     RECT 2.09000000 0.51500000 4.46500000 0.65500000 ;
     RECT 4.17500000 0.65500000 4.46500000 0.73000000 ;
     RECT 2.09000000 0.65500000 2.23000000 0.78500000 ;
     RECT 1.37000000 0.78500000 2.23000000 0.84500000 ;
     RECT 1.29500000 0.84500000 2.23000000 0.92500000 ;
     RECT 1.29500000 0.92500000 1.58500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.38500000 ;
     RECT 1.29500000 1.38500000 1.58500000 1.67500000 ;
     RECT 8.49500000 0.84500000 8.78500000 1.13500000 ;
     RECT 2.73500000 1.25000000 3.02500000 1.32500000 ;
     RECT 8.57000000 1.13500000 8.71000000 1.32500000 ;
     RECT 2.73500000 1.32500000 8.71000000 1.46500000 ;
     RECT 2.73500000 1.46500000 3.02500000 1.54000000 ;
     RECT 8.57000000 1.46500000 8.71000000 1.78000000 ;
     RECT 8.49500000 1.78000000 8.78500000 2.07000000 ;
     RECT 0.57500000 0.44000000 0.86500000 0.73000000 ;
     RECT 5.61500000 0.84500000 5.90500000 0.92000000 ;
     RECT 2.33000000 0.92000000 5.90500000 1.06000000 ;
     RECT 5.61500000 1.06000000 5.90500000 1.13500000 ;
     RECT 0.65000000 0.73000000 0.79000000 1.85500000 ;
     RECT 2.33000000 1.06000000 2.47000000 1.85500000 ;
     RECT 4.17500000 1.78000000 4.46500000 1.85500000 ;
     RECT 0.65000000 1.85500000 4.46500000 1.99500000 ;
     RECT 4.17500000 1.99500000 4.46500000 2.07000000 ;
     RECT 0.65000000 1.99500000 0.79000000 2.19500000 ;
     RECT 0.57500000 2.19500000 0.86500000 2.48500000 ;
     RECT 5.61500000 1.78000000 5.90500000 2.07000000 ;
     RECT 1.29500000 2.19500000 1.58500000 2.27000000 ;
     RECT 5.69000000 2.07000000 5.83000000 2.27000000 ;
     RECT 1.29500000 2.27000000 5.83000000 2.41000000 ;
     RECT 1.29500000 2.41000000 1.58500000 2.48500000 ;
     RECT 8.97500000 0.44000000 9.26500000 0.51500000 ;
     RECT 7.13000000 0.51500000 9.26500000 0.65500000 ;
     RECT 8.97500000 0.65500000 9.26500000 0.73000000 ;
     RECT 7.13000000 0.65500000 7.27000000 0.84500000 ;
     RECT 7.05500000 0.84500000 7.34500000 1.13500000 ;
     RECT 7.05500000 1.78000000 7.34500000 2.07000000 ;
     RECT 9.05000000 0.73000000 9.19000000 2.19500000 ;
     RECT 7.13000000 2.07000000 7.27000000 2.27000000 ;
     RECT 8.97500000 2.19500000 9.26500000 2.27000000 ;
     RECT 7.13000000 2.27000000 9.26500000 2.41000000 ;
     RECT 8.97500000 2.41000000 9.26500000 2.48500000 ;
     RECT 6.09500000 1.65500000 6.38500000 1.94500000 ;
     RECT 5.13500000 2.73500000 5.42500000 2.81000000 ;
     RECT 6.17000000 1.94500000 6.31000000 2.81000000 ;
     RECT 5.13500000 2.81000000 6.31000000 2.95000000 ;
     RECT 5.13500000 2.95000000 5.42500000 3.02500000 ;
     RECT 1.77500000 2.76000000 2.06500000 3.09000000 ;
     RECT 7.53500000 2.76000000 7.82500000 3.09000000 ;
     RECT 0.00000000 3.09000000 10.08000000 3.57000000 ;

 END
END XOR2X1
