magic
tech sky130A
timestamp 1624575530
<< nwell >>
rect 0 179 864 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
rect 713 24 728 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
rect 713 225 728 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 466 67 495 73
rect 466 66 472 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 51 281 66
rect 152 34 184 51
rect 201 34 281 51
rect 152 24 281 34
rect 296 24 425 66
rect 440 50 472 66
rect 489 66 495 67
rect 489 50 569 66
rect 440 24 569 50
rect 584 24 713 66
rect 728 51 807 66
rect 728 34 760 51
rect 777 34 807 51
rect 728 24 807 34
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 299 281 309
rect 152 282 184 299
rect 201 282 281 299
rect 152 225 281 282
rect 296 225 425 309
rect 440 243 569 309
rect 440 226 472 243
rect 489 226 569 243
rect 440 225 569 226
rect 584 225 713 309
rect 728 299 807 309
rect 728 282 760 299
rect 777 282 807 299
rect 728 225 807 282
rect 58 220 87 225
rect 466 220 495 225
<< ndiffc >>
rect 64 50 81 67
rect 184 34 201 51
rect 472 50 489 67
rect 760 34 777 51
<< pdiffc >>
rect 64 226 81 243
rect 184 282 201 299
rect 472 226 489 243
rect 760 282 777 299
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 713 309 728 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 713 209 728 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 713 66 728 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
rect 713 11 728 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 712 184 729 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
rect 712 91 729 108
<< locali >>
rect 0 342 864 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 736 342
rect 753 325 784 342
rect 801 325 832 342
rect 849 325 864 342
rect 0 309 864 325
rect 159 307 226 309
rect 735 307 802 309
rect 176 299 209 307
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 752 299 785 307
rect 752 282 760 299
rect 777 282 785 299
rect 752 274 785 282
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 464 243 497 251
rect 464 226 472 243
rect 489 226 497 243
rect 464 218 497 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 447 209
rect 560 201 593 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 136 162 153 176
rect 280 148 297 176
rect 280 116 297 131
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 92 449 108
rect 441 91 447 92
rect 416 83 447 91
rect 472 75 489 184
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 464 67 497 75
rect 56 42 89 50
rect 176 51 209 59
rect 176 34 184 51
rect 201 34 209 51
rect 464 50 472 67
rect 489 50 497 67
rect 464 42 497 50
rect 752 51 785 59
rect 176 24 209 34
rect 752 34 760 51
rect 777 34 785 51
rect 752 26 785 34
rect 735 24 802 26
rect 0 9 864 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 736 9
rect 753 -9 784 9
rect 801 -9 832 9
rect 849 -9 864 9
rect 0 -24 864 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 304 325 321 342
rect 352 325 369 342
rect 400 325 417 342
rect 448 325 465 342
rect 496 325 513 342
rect 544 325 561 342
rect 592 325 609 342
rect 640 325 657 342
rect 688 325 705 342
rect 736 325 753 342
rect 784 325 801 342
rect 832 325 849 342
rect 184 282 201 299
rect 760 282 777 299
rect 64 226 81 243
rect 472 226 489 243
rect 424 184 441 201
rect 472 184 489 201
rect 136 145 153 162
rect 280 131 297 148
rect 136 91 153 108
rect 424 91 441 108
rect 568 184 585 201
rect 712 184 729 201
rect 568 91 585 108
rect 712 91 729 108
rect 64 50 81 67
rect 184 34 201 51
rect 760 34 777 51
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
rect 304 -9 321 9
rect 352 -9 369 9
rect 400 -9 417 9
rect 448 -9 465 9
rect 496 -9 513 9
rect 544 -9 561 9
rect 592 -9 609 9
rect 640 -9 657 9
rect 688 -9 705 9
rect 736 -9 753 9
rect 784 -9 801 9
rect 832 -9 849 9
<< metal1 >>
rect 0 342 864 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 736 342
rect 753 325 784 342
rect 801 325 832 342
rect 849 325 864 342
rect 0 309 864 325
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 754 299 783 309
rect 754 282 760 299
rect 777 282 783 299
rect 754 276 783 282
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 58 220 87 226
rect 466 243 495 249
rect 466 226 472 243
rect 489 226 495 243
rect 65 200 79 220
rect 418 201 447 207
rect 418 200 424 201
rect 65 186 424 200
rect 65 73 79 186
rect 418 184 424 186
rect 441 184 447 201
rect 418 178 447 184
rect 466 201 495 226
rect 466 184 472 201
rect 489 184 495 201
rect 466 178 495 184
rect 562 201 591 207
rect 562 184 568 201
rect 585 200 591 201
rect 706 201 735 207
rect 585 186 631 200
rect 585 184 591 186
rect 562 178 591 184
rect 130 162 159 168
rect 130 145 136 162
rect 153 145 159 162
rect 425 160 439 178
rect 130 139 159 145
rect 274 148 303 154
rect 137 114 151 139
rect 274 131 280 148
rect 297 131 303 148
rect 425 146 583 160
rect 274 125 303 131
rect 569 114 583 146
rect 130 108 159 114
rect 130 91 136 108
rect 153 106 159 108
rect 418 108 447 114
rect 418 106 424 108
rect 153 92 424 106
rect 153 91 159 92
rect 130 85 159 91
rect 418 91 424 92
rect 441 91 447 108
rect 418 85 447 91
rect 562 108 591 114
rect 562 91 568 108
rect 585 91 591 108
rect 562 85 591 91
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 425 66 439 85
rect 617 66 631 186
rect 706 184 712 201
rect 729 184 735 201
rect 706 178 735 184
rect 713 114 727 178
rect 706 108 735 114
rect 706 91 712 108
rect 729 91 735 108
rect 706 85 735 91
rect 58 44 87 50
rect 178 51 207 57
rect 425 52 631 66
rect 178 34 184 51
rect 201 34 207 51
rect 178 24 207 34
rect 754 51 783 57
rect 754 34 760 51
rect 777 34 783 51
rect 754 24 783 34
rect 0 9 864 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 736 9
rect 753 -9 784 9
rect 801 -9 832 9
rect 849 -9 864 9
rect 0 -24 864 -9
<< labels >>
rlabel metal1 425 52 631 66 0 S
port 6 se
rlabel metal1 425 66 439 85 0 S
port 7 se
rlabel metal1 137 114 151 139 0 S
port 13 se
rlabel metal1 617 66 631 186 0 S
port 16 se
rlabel metal1 713 114 727 178 0 B
port 21 se
rlabel locali 0 309 864 357 0 VDD
port 1 se
rlabel metal1 0 309 864 357 0 VDD
port 2 se
rlabel locali 0 -24 864 24 0 GND
port 3 se
rlabel metal1 0 -24 864 24 0 GND
port 4 se
rlabel metal1 466 178 495 249 0 Y
port 5 se
rlabel metal1 130 85 159 92 0 S
port 8 se
rlabel metal1 418 85 447 92 0 S
port 9 se
rlabel metal1 130 92 447 106 0 S
port 10 se
rlabel metal1 130 106 159 114 0 S
port 11 se
rlabel metal1 418 106 447 114 0 S
port 12 se
rlabel metal1 130 139 159 168 0 S
port 14 se
rlabel metal1 562 178 591 186 0 S
port 15 se
rlabel metal1 562 186 631 200 0 S
port 17 se
rlabel metal1 562 200 591 207 0 S
port 18 se
rlabel metal1 274 125 303 154 0 A
port 19 se
rlabel metal1 706 85 735 114 0 B
port 20 se
rlabel metal1 706 178 735 207 0 B
port 22 se
<< properties >>
string FIXED_BBOX 0 0 864 333
<< end >>
