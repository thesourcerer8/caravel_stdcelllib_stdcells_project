VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 1.780 3.060 2.070 3.090 ;
        RECT 1.780 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.070 3.060 ;
        RECT 1.780 2.830 2.070 2.890 ;
        RECT 7.540 3.060 7.830 3.090 ;
        RECT 7.540 2.890 7.600 3.060 ;
        RECT 7.770 2.890 7.830 3.060 ;
        RECT 7.540 2.830 7.830 2.890 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.360 2.070 0.420 ;
        RECT 1.780 0.240 1.840 0.360 ;
        RECT 2.010 0.240 2.070 0.360 ;
        RECT 7.540 0.240 7.830 0.280 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.150 4.950 2.440 ;
        RECT 4.730 2.040 4.870 2.150 ;
        RECT 4.660 1.750 4.950 2.040 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 8.500 1.750 8.790 2.040 ;
        RECT 8.570 1.090 8.710 1.750 ;
        RECT 8.500 0.800 8.790 1.090 ;
        RECT 3.700 0.610 3.990 0.690 ;
        RECT 5.620 0.610 5.910 0.690 ;
        RECT 8.570 0.610 8.710 0.800 ;
        RECT 3.700 0.470 8.710 0.610 ;
        RECT 3.700 0.400 3.990 0.470 ;
        RECT 5.620 0.400 5.910 0.470 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.960 1.590 2.040 ;
        RECT 2.740 1.960 3.030 2.040 ;
        RECT 1.300 1.820 3.030 1.960 ;
        RECT 1.300 1.750 1.590 1.820 ;
        RECT 2.740 1.750 3.030 1.820 ;
        RECT 1.370 1.500 1.510 1.750 ;
        RECT 1.300 1.210 1.590 1.500 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 1.760 3.060 2.090 3.140 ;
        RECT 1.760 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.090 3.060 ;
        RECT 1.760 2.810 2.090 2.890 ;
        RECT 7.520 3.060 7.850 3.140 ;
        RECT 7.520 2.890 7.600 3.060 ;
        RECT 7.770 2.890 7.850 3.060 ;
        RECT 7.520 2.810 7.850 2.890 ;
        RECT 0.560 2.380 0.890 2.460 ;
        RECT 0.560 2.210 0.640 2.380 ;
        RECT 0.810 2.210 0.890 2.380 ;
        RECT 0.560 2.130 0.890 2.210 ;
        RECT 4.640 2.380 4.970 2.460 ;
        RECT 4.640 2.210 4.720 2.380 ;
        RECT 4.890 2.210 4.970 2.380 ;
        RECT 8.960 2.380 9.290 2.460 ;
        RECT 8.960 2.230 9.040 2.380 ;
        RECT 4.640 2.180 4.970 2.210 ;
        RECT 4.730 2.150 4.970 2.180 ;
        RECT 8.980 2.210 9.040 2.230 ;
        RECT 9.210 2.210 9.290 2.380 ;
        RECT 8.980 2.130 9.290 2.210 ;
        RECT 1.280 1.980 1.610 2.060 ;
        RECT 1.280 1.810 1.360 1.980 ;
        RECT 1.530 1.810 1.610 1.980 ;
        RECT 1.280 1.730 1.610 1.810 ;
        RECT 2.720 1.980 3.050 2.060 ;
        RECT 2.720 1.810 2.800 1.980 ;
        RECT 2.970 1.810 3.050 1.980 ;
        RECT 2.720 1.730 3.050 1.810 ;
        RECT 4.160 2.010 4.470 2.060 ;
        RECT 4.160 1.980 4.490 2.010 ;
        RECT 4.160 1.810 4.240 1.980 ;
        RECT 4.410 1.810 4.490 1.980 ;
        RECT 5.600 1.980 5.930 2.060 ;
        RECT 5.600 1.810 5.680 1.980 ;
        RECT 5.850 1.810 5.930 1.980 ;
        RECT 4.160 1.740 4.490 1.810 ;
        RECT 1.360 1.110 1.530 1.270 ;
        RECT 2.800 1.110 2.970 1.730 ;
        RECT 1.280 1.030 1.610 1.110 ;
        RECT 1.280 0.860 1.360 1.030 ;
        RECT 1.530 0.860 1.610 1.030 ;
        RECT 1.280 0.780 1.610 0.860 ;
        RECT 2.720 1.030 3.050 1.110 ;
        RECT 2.720 0.860 2.800 1.030 ;
        RECT 2.970 0.860 3.050 1.030 ;
        RECT 2.720 0.780 3.050 0.860 ;
        RECT 0.560 0.630 0.890 0.710 ;
        RECT 3.760 0.630 3.930 1.270 ;
        RECT 4.240 1.110 4.410 1.400 ;
        RECT 4.160 1.030 4.490 1.110 ;
        RECT 4.160 0.860 4.240 1.030 ;
        RECT 4.410 0.880 4.490 1.030 ;
        RECT 4.410 0.860 4.470 0.880 ;
        RECT 4.160 0.780 4.470 0.860 ;
        RECT 4.720 0.710 4.890 1.810 ;
        RECT 5.600 1.730 5.930 1.810 ;
        RECT 7.040 1.980 7.370 2.060 ;
        RECT 7.040 1.810 7.120 1.980 ;
        RECT 7.290 1.810 7.370 1.980 ;
        RECT 7.040 1.730 7.370 1.810 ;
        RECT 8.480 1.980 8.810 2.060 ;
        RECT 8.480 1.810 8.560 1.980 ;
        RECT 8.730 1.810 8.810 1.980 ;
        RECT 8.480 1.730 8.810 1.810 ;
        RECT 5.600 1.030 5.930 1.110 ;
        RECT 5.600 0.860 5.680 1.030 ;
        RECT 5.850 0.860 5.930 1.030 ;
        RECT 5.600 0.780 5.930 0.860 ;
        RECT 7.040 1.030 7.370 1.110 ;
        RECT 7.040 0.860 7.120 1.030 ;
        RECT 7.290 0.860 7.370 1.030 ;
        RECT 7.040 0.780 7.370 0.860 ;
        RECT 8.480 1.030 8.810 1.110 ;
        RECT 8.480 0.860 8.560 1.030 ;
        RECT 8.730 0.860 8.810 1.030 ;
        RECT 8.480 0.780 8.810 0.860 ;
        RECT 4.640 0.630 4.970 0.710 ;
        RECT 5.680 0.630 5.850 0.780 ;
        RECT 8.980 0.630 9.290 0.710 ;
        RECT 0.560 0.460 0.640 0.630 ;
        RECT 0.810 0.460 0.890 0.630 ;
        RECT 0.560 0.380 0.890 0.460 ;
        RECT 4.640 0.460 4.720 0.630 ;
        RECT 4.890 0.460 4.970 0.630 ;
        RECT 8.980 0.610 9.040 0.630 ;
        RECT 1.760 0.360 2.090 0.440 ;
        RECT 4.640 0.380 4.970 0.460 ;
        RECT 8.960 0.460 9.040 0.610 ;
        RECT 9.210 0.460 9.290 0.630 ;
        RECT 1.760 0.190 1.840 0.360 ;
        RECT 2.010 0.190 2.090 0.360 ;
        RECT 1.760 0.110 2.090 0.190 ;
        RECT 7.520 0.360 7.850 0.440 ;
        RECT 8.960 0.380 9.290 0.460 ;
        RECT 7.520 0.110 7.600 0.360 ;
        RECT 7.770 0.110 7.850 0.360 ;
      LAYER met1 ;
        RECT 0.580 2.380 0.870 2.440 ;
        RECT 0.580 2.210 0.640 2.380 ;
        RECT 0.810 2.210 0.870 2.380 ;
        RECT 8.980 2.380 9.270 2.440 ;
        RECT 8.980 2.370 9.040 2.380 ;
        RECT 0.580 2.150 0.870 2.210 ;
        RECT 5.690 2.230 9.040 2.370 ;
        RECT 0.650 1.020 0.790 2.150 ;
        RECT 5.690 2.040 5.830 2.230 ;
        RECT 8.980 2.210 9.040 2.230 ;
        RECT 9.210 2.210 9.270 2.380 ;
        RECT 8.980 2.150 9.270 2.210 ;
        RECT 4.180 1.980 4.470 2.040 ;
        RECT 4.180 1.960 4.240 1.980 ;
        RECT 3.770 1.820 4.240 1.960 ;
        RECT 3.770 1.500 3.910 1.820 ;
        RECT 4.180 1.810 4.240 1.820 ;
        RECT 4.410 1.810 4.470 1.980 ;
        RECT 4.180 1.770 4.470 1.810 ;
        RECT 5.620 1.980 5.910 2.040 ;
        RECT 5.620 1.810 5.680 1.980 ;
        RECT 5.850 1.810 5.910 1.980 ;
        RECT 5.620 1.750 5.910 1.810 ;
        RECT 7.060 1.980 7.350 2.040 ;
        RECT 7.060 1.810 7.120 1.980 ;
        RECT 7.290 1.810 7.350 1.980 ;
        RECT 7.060 1.750 7.350 1.810 ;
        RECT 4.180 1.570 4.470 1.630 ;
        RECT 3.700 1.440 3.990 1.500 ;
        RECT 3.700 1.270 3.760 1.440 ;
        RECT 3.930 1.270 3.990 1.440 ;
        RECT 4.180 1.400 4.240 1.570 ;
        RECT 4.410 1.560 4.470 1.570 ;
        RECT 5.690 1.560 5.830 1.750 ;
        RECT 4.410 1.420 5.830 1.560 ;
        RECT 4.410 1.400 4.470 1.420 ;
        RECT 4.180 1.340 4.470 1.400 ;
        RECT 3.700 1.210 3.990 1.270 ;
        RECT 7.130 1.090 7.270 1.750 ;
        RECT 7.060 1.030 7.350 1.090 ;
        RECT 7.060 1.020 7.120 1.030 ;
        RECT 0.650 0.880 7.120 1.020 ;
        RECT 0.650 0.690 0.790 0.880 ;
        RECT 7.060 0.860 7.120 0.880 ;
        RECT 7.290 0.860 7.350 1.030 ;
        RECT 7.060 0.800 7.350 0.860 ;
        RECT 9.050 0.690 9.190 2.150 ;
        RECT 0.580 0.630 0.870 0.690 ;
        RECT 0.580 0.460 0.640 0.630 ;
        RECT 0.810 0.460 0.870 0.630 ;
        RECT 0.580 0.400 0.870 0.460 ;
        RECT 8.980 0.630 9.270 0.690 ;
        RECT 8.980 0.460 9.040 0.630 ;
        RECT 9.210 0.460 9.270 0.630 ;
        RECT 8.980 0.400 9.270 0.460 ;
  END
END XNOR2X1
END LIBRARY

