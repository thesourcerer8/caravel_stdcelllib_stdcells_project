MACRO INVX8
 CLASS CORE ;
 FOREIGN INVX8 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 7.20000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 7.20000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.57500000 0.39500000 0.86500000 0.47000000 ;
        RECT 3.21500000 0.39500000 3.50500000 0.47000000 ;
        RECT 6.09500000 0.39500000 6.38500000 0.47000000 ;
        RECT 0.57500000 0.47000000 6.38500000 0.61000000 ;
        RECT 0.57500000 0.61000000 0.86500000 0.68500000 ;
        RECT 3.21500000 0.61000000 3.50500000 0.68500000 ;
        RECT 6.09500000 0.61000000 6.38500000 0.68500000 ;
        RECT 0.65000000 0.68500000 0.79000000 2.15000000 ;
        RECT 6.17000000 0.68500000 6.31000000 2.15000000 ;
        RECT 0.57500000 2.15000000 0.86500000 2.22500000 ;
        RECT 3.21500000 2.15000000 3.50500000 2.22500000 ;
        RECT 0.57500000 2.22500000 3.50500000 2.36500000 ;
        RECT 0.57500000 2.36500000 0.86500000 2.44000000 ;
        RECT 3.21500000 2.36500000 3.50500000 2.44000000 ;
        RECT 6.09500000 2.15000000 6.38500000 2.44000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.29500000 0.80000000 1.58500000 1.09000000 ;
        RECT 2.73500000 0.80000000 3.02500000 1.09000000 ;
        RECT 4.17500000 0.80000000 4.46500000 1.09000000 ;
        RECT 5.61500000 0.80000000 5.90500000 1.09000000 ;
        RECT 1.37000000 1.09000000 1.51000000 1.74500000 ;
        RECT 2.81000000 1.09000000 2.95000000 1.74500000 ;
        RECT 4.25000000 1.09000000 4.39000000 1.74500000 ;
        RECT 5.69000000 1.09000000 5.83000000 1.74500000 ;
        RECT 1.29500000 1.74500000 1.58500000 1.82000000 ;
        RECT 2.73500000 1.74500000 3.02500000 1.82000000 ;
        RECT 4.17500000 1.74500000 4.46500000 1.82000000 ;
        RECT 5.61500000 1.74500000 5.90500000 1.82000000 ;
        RECT 1.29500000 1.82000000 5.90500000 1.96000000 ;
        RECT 1.29500000 1.96000000 1.58500000 2.03500000 ;
        RECT 2.73500000 1.96000000 3.02500000 2.03500000 ;
        RECT 4.17500000 1.96000000 4.46500000 2.03500000 ;
        RECT 5.61500000 1.96000000 5.90500000 2.03500000 ;
    END
  END A


END INVX8
