VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO VANBERKEL1991
  CLASS CORE ;
  FOREIGN VANBERKEL1991 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
        RECT 1.370 0.655 1.510 0.845 ;
        RECT 3.215 0.655 3.505 0.730 ;
        RECT 1.370 0.515 3.505 0.655 ;
        RECT 3.215 0.440 3.505 0.515 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 1.060 3.025 1.135 ;
        RECT 8.495 1.060 8.785 1.135 ;
        RECT 2.735 0.920 8.785 1.060 ;
        RECT 2.735 0.845 3.025 0.920 ;
        RECT 8.495 0.845 8.785 0.920 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.189000 ;
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 7.055 2.410 7.345 2.485 ;
        RECT 10.415 2.410 10.705 2.485 ;
        RECT 7.055 2.270 10.705 2.410 ;
        RECT 7.055 2.195 7.345 2.270 ;
        RECT 10.415 2.195 10.705 2.270 ;
        RECT 10.490 0.730 10.630 2.195 ;
        RECT 10.415 0.440 10.705 0.730 ;
    END
  END C
  PIN VGND
    ANTENNADIFFAREA 0.914200 ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.520 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 11.520 3.570 ;
        RECT 8.975 2.735 9.265 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.747200 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 11.520 3.415 ;
        RECT 0.155 3.090 11.365 3.245 ;
        RECT 4.635 2.715 4.965 3.090 ;
        RECT 8.955 2.715 9.285 3.090 ;
      LAYER mcon ;
        RECT 4.715 3.245 4.885 3.415 ;
        RECT 9.035 2.795 9.205 2.965 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 11.520 3.330 ;
      LAYER li1 ;
        RECT 0.795 2.580 1.125 2.910 ;
        RECT 7.515 2.580 7.845 2.910 ;
        RECT 1.755 2.260 2.085 2.505 ;
        RECT 1.775 2.175 2.085 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 1.835 0.750 2.005 2.175 ;
        RECT 2.315 1.310 2.485 2.290 ;
        RECT 3.675 2.260 4.005 2.505 ;
        RECT 3.675 2.175 3.985 2.260 ;
        RECT 6.315 2.175 6.645 2.505 ;
        RECT 7.115 2.090 7.285 2.425 ;
        RECT 10.395 2.260 10.725 2.505 ;
        RECT 10.415 2.175 10.725 2.260 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 9.915 1.760 10.245 2.090 ;
        RECT 2.795 1.155 2.965 1.760 ;
        RECT 4.235 1.210 4.405 1.760 ;
        RECT 3.275 1.155 4.405 1.210 ;
        RECT 7.115 1.155 7.285 1.760 ;
        RECT 8.555 1.155 8.725 1.760 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 3.275 1.040 4.485 1.155 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.275 0.500 3.445 1.040 ;
        RECT 4.155 0.920 4.485 1.040 ;
        RECT 4.155 0.825 4.465 0.920 ;
        RECT 7.035 0.825 7.365 1.155 ;
        RECT 8.475 0.920 8.805 1.155 ;
        RECT 9.915 0.920 10.245 1.155 ;
        RECT 8.495 0.825 8.785 0.920 ;
        RECT 9.915 0.825 10.225 0.920 ;
        RECT 3.675 0.655 3.985 0.750 ;
        RECT 3.675 0.420 4.005 0.655 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 6.315 0.420 6.645 0.750 ;
        RECT 7.995 0.420 8.325 0.750 ;
        RECT 8.955 0.420 9.285 0.750 ;
        RECT 10.395 0.420 10.725 0.750 ;
        RECT 4.715 0.240 4.885 0.420 ;
        RECT 9.035 0.240 9.205 0.420 ;
        RECT 0.155 0.085 11.365 0.240 ;
        RECT 0.000 -0.085 11.520 0.085 ;
      LAYER mcon ;
        RECT 0.875 2.660 1.045 2.830 ;
        RECT 7.595 2.660 7.765 2.830 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 1.835 1.715 2.005 1.885 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.315 2.120 2.485 2.290 ;
        RECT 3.755 2.255 3.925 2.425 ;
        RECT 6.395 2.255 6.565 2.425 ;
        RECT 7.115 2.255 7.285 2.425 ;
        RECT 10.475 2.255 10.645 2.425 ;
        RECT 9.995 1.840 10.165 2.010 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 8.555 0.905 8.725 1.075 ;
        RECT 9.995 0.905 10.165 1.075 ;
        RECT 3.755 0.500 3.925 0.670 ;
        RECT 6.395 0.500 6.565 0.670 ;
        RECT 8.075 0.500 8.245 0.670 ;
        RECT 10.475 0.500 10.645 0.670 ;
        RECT 9.035 -0.085 9.205 0.085 ;
      LAYER met1 ;
        RECT 0.815 2.815 1.105 2.890 ;
        RECT 7.535 2.815 7.825 2.890 ;
        RECT 0.815 2.675 7.825 2.815 ;
        RECT 0.815 2.600 1.105 2.675 ;
        RECT 7.535 2.600 7.825 2.675 ;
        RECT 3.695 2.410 3.985 2.485 ;
        RECT 6.335 2.410 6.625 2.485 ;
        RECT 0.650 2.350 2.470 2.410 ;
        RECT 0.650 2.270 2.545 2.350 ;
        RECT 0.650 0.730 0.790 2.270 ;
        RECT 2.255 2.060 2.545 2.270 ;
        RECT 3.695 2.270 6.625 2.410 ;
        RECT 3.695 2.195 3.985 2.270 ;
        RECT 6.335 2.195 6.625 2.270 ;
        RECT 1.775 1.870 2.065 1.945 ;
        RECT 9.935 1.870 10.225 2.070 ;
        RECT 1.775 1.780 10.225 1.870 ;
        RECT 1.775 1.730 10.150 1.780 ;
        RECT 1.775 1.655 2.065 1.730 ;
        RECT 2.255 1.465 2.545 1.540 ;
        RECT 2.255 1.325 9.190 1.465 ;
        RECT 2.255 1.250 2.545 1.325 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 3.695 0.655 3.985 0.730 ;
        RECT 6.335 0.655 6.625 0.730 ;
        RECT 3.695 0.515 6.625 0.655 ;
        RECT 3.695 0.440 3.985 0.515 ;
        RECT 6.335 0.440 6.625 0.515 ;
        RECT 8.015 0.655 8.305 0.730 ;
        RECT 9.050 0.655 9.190 1.325 ;
        RECT 10.010 1.135 10.150 1.730 ;
        RECT 9.935 0.845 10.225 1.135 ;
        RECT 8.015 0.515 9.190 0.655 ;
        RECT 8.015 0.440 8.305 0.515 ;
  END
END VANBERKEL1991
END LIBRARY

