magic
tech sky130A
magscale 1 2
timestamp 1636809583
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 2304 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1425 48 1455 132
rect 1713 48 1743 132
rect 2001 48 2031 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1425 450 1455 618
rect 1713 450 1743 618
rect 2001 450 2031 618
<< ndiff >>
rect 163 134 221 146
rect 163 132 175 134
rect 115 100 175 132
rect 209 132 221 134
rect 355 134 413 146
rect 355 132 367 134
rect 209 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 739 134 797 146
rect 739 132 751 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 100 751 132
rect 785 132 797 134
rect 931 134 989 146
rect 931 132 943 134
rect 785 100 849 132
rect 591 48 849 100
rect 879 100 943 132
rect 977 132 989 134
rect 1267 134 1325 146
rect 977 100 1037 132
rect 879 48 1037 100
rect 1267 100 1279 134
rect 1313 132 1325 134
rect 1507 134 1565 146
rect 1507 132 1519 134
rect 1313 100 1425 132
rect 1267 48 1425 100
rect 1455 100 1519 132
rect 1553 132 1565 134
rect 1795 134 1853 146
rect 1795 132 1807 134
rect 1553 100 1713 132
rect 1455 48 1713 100
rect 1743 100 1807 132
rect 1841 132 1853 134
rect 2083 134 2141 146
rect 2083 132 2095 134
rect 1841 100 2001 132
rect 1743 48 2001 100
rect 2031 100 2095 132
rect 2129 132 2141 134
rect 2129 100 2189 132
rect 2031 48 2189 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 175 485
rect 209 451 273 485
rect 115 450 273 451
rect 303 485 561 618
rect 303 451 367 485
rect 401 451 561 485
rect 303 450 561 451
rect 591 566 849 618
rect 591 532 751 566
rect 785 532 849 566
rect 591 450 849 532
rect 879 593 1037 618
rect 879 559 943 593
rect 977 559 1037 593
rect 879 450 1037 559
rect 1267 566 1425 618
rect 1267 532 1279 566
rect 1313 532 1425 566
rect 1267 450 1425 532
rect 1455 485 1713 618
rect 1455 451 1519 485
rect 1553 451 1713 485
rect 1455 450 1713 451
rect 1743 593 2001 618
rect 1743 559 1807 593
rect 1841 559 2001 593
rect 1743 450 2001 559
rect 2031 485 2189 618
rect 2031 451 2095 485
rect 2129 451 2189 485
rect 2031 450 2189 451
rect 163 439 221 450
rect 355 439 413 450
rect 1507 439 1565 450
rect 2083 439 2141 450
<< ndiffc >>
rect 175 100 209 134
rect 367 100 401 134
rect 751 100 785 134
rect 943 100 977 134
rect 1279 100 1313 134
rect 1519 100 1553 134
rect 1807 100 1841 134
rect 2095 100 2129 134
<< pdiffc >>
rect 175 451 209 485
rect 367 451 401 485
rect 751 532 785 566
rect 943 559 977 593
rect 1279 532 1313 566
rect 1519 451 1553 485
rect 1807 559 1841 593
rect 2095 451 2129 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1425 618 1455 644
rect 1713 618 1743 644
rect 2001 618 2031 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1425 418 1455 450
rect 1713 418 1743 450
rect 2001 418 2031 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1425 132 1455 165
rect 1713 132 1743 165
rect 2001 132 2031 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1425 22 1455 48
rect 1713 22 1743 48
rect 2001 22 2031 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 1999 181 2033 215
<< locali >>
rect 0 649 943 683
rect 977 649 2304 683
rect 31 618 2273 649
rect 927 593 993 618
rect 735 566 801 582
rect 735 532 751 566
rect 785 532 801 566
rect 927 559 943 593
rect 977 559 993 593
rect 1791 593 1857 618
rect 927 543 993 559
rect 1263 566 1329 582
rect 735 516 801 532
rect 1263 532 1279 566
rect 1313 532 1329 566
rect 1791 559 1807 593
rect 1841 559 1857 593
rect 1791 543 1857 559
rect 1263 516 1329 532
rect 159 485 225 501
rect 159 451 175 485
rect 209 452 225 485
rect 351 485 417 501
rect 209 451 221 452
rect 159 435 221 451
rect 351 451 367 485
rect 401 451 417 485
rect 1503 485 1569 501
rect 1503 452 1519 485
rect 351 435 417 451
rect 1507 451 1519 452
rect 1553 451 1569 485
rect 2079 485 2145 501
rect 2079 452 2095 485
rect 1507 435 1569 451
rect 2083 451 2095 452
rect 2129 451 2145 485
rect 2083 435 2145 451
rect 255 402 317 418
rect 255 368 271 402
rect 305 401 317 402
rect 367 402 401 435
rect 305 368 321 401
rect 255 352 321 368
rect 271 231 305 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 184 321 215
rect 305 181 317 184
rect 255 165 317 181
rect 367 150 401 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 559 231 593 352
rect 847 242 881 352
rect 655 231 881 242
rect 1423 231 1457 352
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 655 215 897 231
rect 655 208 847 215
rect 159 134 221 150
rect 159 100 175 134
rect 209 131 221 134
rect 351 134 417 150
rect 209 100 225 131
rect 159 84 225 100
rect 351 100 367 134
rect 401 100 417 134
rect 655 134 689 208
rect 831 184 847 208
rect 835 181 847 184
rect 881 184 897 215
rect 1407 215 1473 231
rect 881 181 893 184
rect 835 165 893 181
rect 1407 181 1423 215
rect 1457 184 1473 215
rect 1457 181 1469 184
rect 1407 165 1469 181
rect 735 134 801 150
rect 735 100 751 134
rect 785 100 801 134
rect 351 84 417 100
rect 735 84 801 100
rect 927 134 993 150
rect 927 100 943 134
rect 977 100 993 134
rect 927 84 993 100
rect 1263 134 1329 150
rect 1263 100 1279 134
rect 1313 100 1329 134
rect 1423 134 1457 165
rect 1519 150 1553 289
rect 1711 231 1745 352
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 184 1761 215
rect 1983 215 2049 231
rect 1745 181 1757 184
rect 1695 165 1757 181
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 1503 134 1569 150
rect 1503 100 1519 134
rect 1553 100 1569 134
rect 1263 84 1329 100
rect 1503 84 1569 100
rect 1791 134 1857 150
rect 1791 100 1807 134
rect 1841 100 1857 134
rect 2083 134 2145 150
rect 2083 131 2095 134
rect 1791 84 1857 100
rect 2079 100 2095 131
rect 2129 100 2145 134
rect 2079 84 2145 100
rect 943 48 977 84
rect 1807 48 1841 84
rect 31 17 2273 48
rect 0 -17 1807 17
rect 1841 -17 2304 17
<< viali >>
rect 943 649 977 683
rect 751 532 785 566
rect 1279 532 1313 566
rect 1807 559 1841 593
rect 175 451 209 485
rect 1519 451 1553 485
rect 2095 451 2129 485
rect 367 368 401 402
rect 271 181 305 215
rect 1999 368 2033 402
rect 1519 289 1553 323
rect 559 181 593 215
rect 175 100 209 134
rect 655 100 689 134
rect 751 100 785 134
rect 1279 100 1313 134
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 1423 100 1457 134
rect 2095 100 2129 134
rect 1807 -17 1841 17
<< metal1 >>
rect 0 683 2304 714
rect 0 649 943 683
rect 977 649 2304 683
rect 0 618 2304 649
rect 1795 593 1853 618
rect 739 566 797 578
rect 739 532 751 566
rect 785 563 797 566
rect 1267 566 1325 578
rect 1267 563 1279 566
rect 785 535 1279 563
rect 785 532 797 535
rect 739 520 797 532
rect 1267 532 1279 535
rect 1313 532 1325 566
rect 1795 559 1807 593
rect 1841 559 1853 593
rect 1795 547 1853 559
rect 1267 520 1325 532
rect 163 485 221 497
rect 163 451 175 485
rect 209 482 221 485
rect 1507 485 1565 497
rect 1507 482 1519 485
rect 209 454 1519 482
rect 209 451 221 454
rect 163 439 221 451
rect 1507 451 1519 454
rect 1553 451 1565 485
rect 1507 439 1565 451
rect 2083 485 2141 497
rect 2083 451 2095 485
rect 2129 451 2141 485
rect 2083 439 2141 451
rect 355 402 413 414
rect 355 368 367 402
rect 401 399 413 402
rect 1987 402 2045 414
rect 1987 399 1999 402
rect 401 371 1999 399
rect 401 368 413 371
rect 355 356 413 368
rect 1987 368 1999 371
rect 2033 368 2045 402
rect 1987 356 2045 368
rect 1507 323 1565 335
rect 1507 320 1519 323
rect 178 292 1519 320
rect 178 146 206 292
rect 1507 289 1519 292
rect 1553 289 1565 323
rect 1507 277 1565 289
rect 2002 227 2030 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 212 605 215
rect 1699 215 1757 227
rect 1699 212 1711 215
rect 593 184 1711 212
rect 593 181 605 184
rect 547 169 605 181
rect 1699 181 1711 184
rect 1745 181 1757 215
rect 1699 169 1757 181
rect 1987 215 2045 227
rect 1987 181 1999 215
rect 2033 181 2045 215
rect 1987 169 2045 181
rect 163 134 221 146
rect 163 100 175 134
rect 209 100 221 134
rect 274 131 302 169
rect 2098 146 2126 439
rect 643 134 701 146
rect 643 131 655 134
rect 274 103 655 131
rect 163 88 221 100
rect 643 100 655 103
rect 689 100 701 134
rect 643 88 701 100
rect 739 134 797 146
rect 739 100 751 134
rect 785 131 797 134
rect 1267 134 1325 146
rect 1267 131 1279 134
rect 785 103 1279 131
rect 785 100 797 103
rect 739 88 797 100
rect 1267 100 1279 103
rect 1313 100 1325 134
rect 1267 88 1325 100
rect 1411 134 1469 146
rect 1411 100 1423 134
rect 1457 131 1469 134
rect 2083 134 2141 146
rect 2083 131 2095 134
rect 1457 103 2095 131
rect 1457 100 1469 103
rect 1411 88 1469 100
rect 2083 100 2095 103
rect 2129 100 2141 134
rect 2083 88 2141 100
rect 0 17 2304 48
rect 0 -17 1807 17
rect 1841 -17 2304 17
rect 0 -48 2304 -17
<< labels >>
rlabel metal1 0 618 2304 714 0 VPWR
port 5 se
rlabel metal1 0 618 2304 714 0 VPWR
port 5 se
rlabel metal1 0 -48 2304 48 0 VGND
port 4 se
rlabel metal1 0 -48 2304 48 0 VGND
port 4 se
rlabel metal1 1987 169 2045 227 0 CN
port 3 se
rlabel metal1 2002 227 2030 356 0 CN
port 3 se
rlabel metal1 355 356 413 371 0 CN
port 3 se
rlabel metal1 1987 356 2045 371 0 CN
port 3 se
rlabel metal1 355 371 2045 399 0 CN
port 3 se
rlabel metal1 355 399 413 414 0 CN
port 3 se
rlabel metal1 1987 399 2045 414 0 CN
port 3 se
rlabel metal1 1411 88 1469 103 0 C
port 2 se
rlabel metal1 2083 88 2141 103 0 C
port 2 se
rlabel metal1 1411 103 2141 131 0 C
port 2 se
rlabel metal1 1411 131 1469 146 0 C
port 2 se
rlabel metal1 2083 131 2141 146 0 C
port 2 se
rlabel metal1 2098 146 2126 439 0 C
port 2 se
rlabel metal1 2083 439 2141 497 0 C
port 2 se
rlabel metal1 643 88 701 103 0 A
port 0 se
rlabel metal1 274 103 701 131 0 A
port 0 se
rlabel metal1 643 131 701 146 0 A
port 0 se
rlabel metal1 274 131 302 169 0 A
port 0 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 547 169 605 184 0 B
port 1 se
rlabel metal1 1699 169 1757 184 0 B
port 1 se
rlabel metal1 547 184 1757 212 0 B
port 1 se
rlabel metal1 547 212 605 227 0 B
port 1 se
rlabel metal1 1699 212 1757 227 0 B
port 1 se
rlabel locali 0 -17 2304 17 4 VGND
port 4 se ground default abutment
rlabel locali 31 17 2273 48 4 VGND
port 4 se ground default abutment
rlabel locali 0 649 2304 683 4 VPWR
port 5 se power default abutment
rlabel locali 31 618 2273 649 4 VGND
port 4 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 2304 666
<< end >>
