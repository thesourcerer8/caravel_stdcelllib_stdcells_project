magic
tech sky130A
timestamp 1624064557
<< nwell >>
rect 0 179 432 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 322 67 351 73
rect 322 66 328 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 49 281 66
rect 152 32 184 49
rect 201 32 281 49
rect 152 24 281 32
rect 296 50 328 66
rect 345 66 351 67
rect 345 50 375 66
rect 296 24 375 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 301 281 309
rect 152 284 184 301
rect 201 284 281 301
rect 152 225 281 284
rect 296 243 375 309
rect 296 226 328 243
rect 345 226 375 243
rect 296 225 375 226
rect 58 220 87 225
rect 322 220 351 225
<< ndiffc >>
rect 64 50 81 67
rect 184 32 201 49
rect 328 50 345 67
<< pdiffc >>
rect 64 226 81 243
rect 184 284 201 301
rect 328 226 345 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 137 209 152 225
rect 281 209 296 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 137 66 152 83
rect 281 66 296 83
rect 137 11 152 24
rect 281 11 296 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 136 91 153 108
rect 280 91 297 108
<< locali >>
rect 176 301 209 309
rect 176 284 184 301
rect 201 284 209 301
rect 176 276 209 284
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 320 243 353 251
rect 320 226 328 243
rect 345 226 353 243
rect 320 218 353 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 303 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 136 116 153 176
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 92 305 108
rect 297 91 303 92
rect 272 83 303 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 320 67 353 75
rect 56 42 89 50
rect 176 49 209 57
rect 176 32 184 49
rect 201 32 209 49
rect 320 50 328 67
rect 345 50 353 67
rect 320 42 353 50
rect 176 24 209 32
<< viali >>
rect 184 284 201 301
rect 64 226 81 243
rect 328 226 345 243
rect 136 184 153 201
rect 280 184 297 201
rect 280 91 297 108
rect 64 50 81 67
rect 184 32 201 49
rect 328 50 345 67
<< metal1 >>
rect 0 309 432 357
rect 178 301 207 309
rect 178 284 184 301
rect 201 284 207 301
rect 178 278 207 284
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 58 220 87 226
rect 322 243 351 249
rect 322 226 328 243
rect 345 226 351 243
rect 322 220 351 226
rect 65 106 79 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 281 114 295 178
rect 274 108 303 114
rect 274 106 280 108
rect 65 92 280 106
rect 65 73 79 92
rect 274 91 280 92
rect 297 91 303 108
rect 274 85 303 91
rect 329 73 343 220
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 322 67 351 73
rect 58 44 87 50
rect 178 49 207 55
rect 178 32 184 49
rect 201 32 207 49
rect 322 50 328 67
rect 345 50 351 67
rect 322 44 351 50
rect 178 24 207 32
rect 0 -24 432 24
<< labels >>
rlabel metal1 0 309 432 357 0 VDD
port 1 se
rlabel metal1 0 -24 432 24 0 GND
port 2 se
rlabel metal1 322 44 351 73 0 Y
port 3 se
rlabel metal1 329 73 343 220 0 Y
port 4 se
rlabel metal1 322 220 351 249 0 Y
port 5 se
rlabel metal1 130 178 159 207 0 A
port 6 se
<< properties >>
string FIXED_BBOX 0 0 432 333
<< end >>
