magic
tech sky130A
magscale 1 2
timestamp 1624892581
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 576 666
<< nmos >>
rect 273 48 303 132
<< pmos >>
rect 273 450 303 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 102 461 132
rect 303 68 367 102
rect 401 68 461 102
rect 303 48 461 68
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 598 461 618
rect 303 564 367 598
rect 401 564 461 598
rect 303 450 461 564
rect 115 439 173 450
<< ndiffc >>
rect 127 100 161 134
rect 367 68 401 102
<< pdiffc >>
rect 127 451 161 485
rect 367 564 401 598
<< poly >>
rect 273 618 303 644
rect 273 418 303 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 273 132 303 165
rect 273 22 303 48
<< polycont >>
rect 271 368 305 402
rect 271 181 305 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 31 618 545 649
rect 351 598 417 618
rect 351 564 367 598
rect 401 564 417 598
rect 351 548 417 564
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 351 102 417 118
rect 351 68 367 102
rect 401 68 417 102
rect 351 48 417 68
rect 31 17 545 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 367 564 401 598
rect 127 451 161 485
rect 271 368 305 402
rect 271 181 305 215
rect 127 100 161 134
rect 367 68 401 102
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 714
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 618 576 649
rect 355 598 413 618
rect 355 564 367 598
rect 401 564 413 598
rect 355 552 413 564
rect 115 485 173 497
rect 115 451 127 485
rect 161 451 173 485
rect 115 439 173 451
rect 130 146 158 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 274 227 302 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 355 102 413 114
rect 355 68 367 102
rect 401 68 413 102
rect 355 48 413 68
rect 0 17 576 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -48 576 -17
<< labels >>
rlabel metal1 0 618 576 714 0 VDD
port 2 se
rlabel metal1 0 618 576 714 0 VDD
port 2 se
rlabel metal1 0 -48 576 48 0 GND
port 1 se
rlabel metal1 0 -48 576 48 0 GND
port 1 se
rlabel metal1 115 88 173 146 0 Y
port 3 se
rlabel metal1 130 146 158 439 0 Y
port 3 se
rlabel metal1 115 439 173 497 0 Y
port 3 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel locali 0 -17 576 17 4 GND
port 1 se ground default abutment
rlabel locali 31 17 545 48 4 GND
port 1 se ground default abutment
rlabel locali 0 649 576 683 4 VDD
port 2 se power default abutment
rlabel locali 31 618 545 649 4 VDD
port 2 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 576 666
<< end >>
