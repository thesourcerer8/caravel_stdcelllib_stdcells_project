VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 1.780 2.970 2.070 3.090 ;
        RECT 1.780 2.800 1.840 2.970 ;
        RECT 2.010 2.800 2.070 2.970 ;
        RECT 1.780 2.740 2.070 2.800 ;
        RECT 7.540 2.970 7.830 3.090 ;
        RECT 7.540 2.800 7.600 2.970 ;
        RECT 7.770 2.800 7.830 2.970 ;
        RECT 7.540 2.740 7.830 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 1.760 2.970 2.090 3.090 ;
        RECT 1.760 2.800 1.840 2.970 ;
        RECT 2.010 2.800 2.090 2.970 ;
        RECT 1.760 2.720 2.090 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.780 0.670 2.090 0.750 ;
        RECT 1.780 0.660 1.840 0.670 ;
        RECT 1.760 0.500 1.840 0.660 ;
        RECT 2.010 0.500 2.090 0.670 ;
        RECT 7.540 0.670 7.850 0.750 ;
        RECT 7.540 0.660 7.600 0.670 ;
        RECT 1.760 0.420 2.090 0.500 ;
        RECT 7.520 0.500 7.600 0.660 ;
        RECT 7.770 0.500 7.850 0.670 ;
        RECT 7.520 0.420 7.850 0.500 ;
        RECT 1.840 0.240 2.010 0.420 ;
        RECT 7.600 0.240 7.770 0.420 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.600 4.950 2.890 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 5.620 2.000 5.910 2.070 ;
        RECT 4.250 1.860 5.910 2.000 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 4.250 1.140 4.390 1.860 ;
        RECT 5.620 1.780 5.910 1.860 ;
        RECT 1.300 1.060 1.590 1.140 ;
        RECT 4.180 1.060 4.470 1.140 ;
        RECT 1.300 0.920 4.470 1.060 ;
        RECT 1.300 0.850 1.590 0.920 ;
        RECT 4.180 0.850 4.470 0.920 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.810 2.270 8.710 2.410 ;
        RECT 2.810 2.070 2.950 2.270 ;
        RECT 8.570 2.070 8.710 2.270 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 8.500 1.780 8.790 2.070 ;
        RECT 8.570 1.140 8.710 1.780 ;
        RECT 8.500 0.850 8.790 1.140 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 7.520 2.970 7.850 3.050 ;
        RECT 4.640 2.830 4.970 2.910 ;
        RECT 4.640 2.660 4.720 2.830 ;
        RECT 4.890 2.660 4.970 2.830 ;
        RECT 7.520 2.800 7.600 2.970 ;
        RECT 7.770 2.800 7.850 2.970 ;
        RECT 7.520 2.720 7.850 2.800 ;
        RECT 4.640 2.580 4.970 2.660 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 5.140 2.430 5.450 2.510 ;
        RECT 5.140 2.410 5.200 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 5.120 2.260 5.200 2.410 ;
        RECT 5.370 2.260 5.450 2.430 ;
        RECT 8.960 2.430 9.290 2.510 ;
        RECT 8.960 2.260 9.040 2.430 ;
        RECT 9.210 2.260 9.290 2.430 ;
        RECT 5.120 2.180 5.450 2.260 ;
        RECT 8.980 2.180 9.290 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.890 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 2.800 1.160 2.970 1.760 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 4.720 0.670 4.890 1.840 ;
        RECT 5.200 0.750 5.370 2.180 ;
        RECT 5.620 2.010 5.930 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 7.040 2.010 7.370 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 8.480 2.010 8.810 2.090 ;
        RECT 8.480 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.810 2.010 ;
        RECT 8.480 1.760 8.810 1.840 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.920 5.680 1.080 ;
        RECT 5.620 0.910 5.680 0.920 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.620 0.830 5.930 0.910 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.370 1.080 ;
        RECT 7.040 0.830 7.370 0.910 ;
        RECT 8.480 1.080 8.810 1.160 ;
        RECT 8.480 0.910 8.560 1.080 ;
        RECT 8.730 0.920 8.810 1.080 ;
        RECT 8.730 0.910 8.790 0.920 ;
        RECT 8.480 0.830 8.790 0.910 ;
        RECT 5.120 0.670 5.450 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 5.120 0.500 5.200 0.670 ;
        RECT 5.370 0.500 5.450 0.670 ;
        RECT 5.120 0.420 5.450 0.500 ;
        RECT 8.960 0.670 9.290 0.750 ;
        RECT 8.960 0.500 9.040 0.670 ;
        RECT 9.210 0.500 9.290 0.670 ;
        RECT 8.960 0.420 9.290 0.500 ;
      LAYER met1 ;
        RECT 0.580 2.430 0.870 2.490 ;
        RECT 0.580 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.870 2.430 ;
        RECT 0.580 2.200 0.870 2.260 ;
        RECT 8.980 2.430 9.270 2.490 ;
        RECT 8.980 2.260 9.040 2.430 ;
        RECT 9.210 2.260 9.270 2.430 ;
        RECT 8.980 2.200 9.270 2.260 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 7.060 2.010 7.350 2.070 ;
        RECT 7.060 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.350 2.010 ;
        RECT 7.060 1.780 7.350 1.840 ;
        RECT 7.130 1.140 7.270 1.780 ;
        RECT 5.620 1.080 5.910 1.140 ;
        RECT 5.620 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.910 1.080 ;
        RECT 5.620 0.850 5.910 0.910 ;
        RECT 7.060 1.080 7.350 1.140 ;
        RECT 7.060 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.350 1.080 ;
        RECT 7.060 0.850 7.350 0.910 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.660 0.870 0.670 ;
        RECT 4.660 0.670 4.950 0.730 ;
        RECT 4.660 0.660 4.720 0.670 ;
        RECT 0.810 0.520 4.720 0.660 ;
        RECT 0.810 0.500 0.870 0.520 ;
        RECT 0.580 0.440 0.870 0.500 ;
        RECT 4.660 0.500 4.720 0.520 ;
        RECT 4.890 0.660 4.950 0.670 ;
        RECT 5.690 0.660 5.830 0.850 ;
        RECT 4.890 0.520 5.830 0.660 ;
        RECT 7.130 0.660 7.270 0.850 ;
        RECT 9.050 0.730 9.190 2.200 ;
        RECT 8.980 0.670 9.270 0.730 ;
        RECT 8.980 0.660 9.040 0.670 ;
        RECT 7.130 0.520 9.040 0.660 ;
        RECT 4.890 0.500 4.950 0.520 ;
        RECT 4.660 0.440 4.950 0.500 ;
        RECT 8.980 0.500 9.040 0.520 ;
        RECT 9.210 0.500 9.270 0.670 ;
        RECT 8.980 0.440 9.270 0.500 ;
  END
END XOR2X1
END LIBRARY

