VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SUTHERLAND1989
  CLASS CORE ;
  FOREIGN SUTHERLAND1989 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 1.060 3.025 1.135 ;
        RECT 4.175 1.060 4.465 1.135 ;
        RECT 2.735 0.920 4.465 1.060 ;
        RECT 2.735 0.845 3.025 0.920 ;
        RECT 4.175 0.845 4.465 0.920 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.995 1.585 2.070 ;
        RECT 5.615 1.995 5.905 2.070 ;
        RECT 1.295 1.855 5.905 1.995 ;
        RECT 1.295 1.780 1.585 1.855 ;
        RECT 5.615 1.780 5.905 1.855 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 5.690 1.135 5.830 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
        RECT 5.615 0.845 5.905 1.135 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.189000 ;
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.060 8.065 1.135 ;
        RECT 9.935 1.060 10.225 1.135 ;
        RECT 7.775 0.920 10.225 1.060 ;
        RECT 7.775 0.845 8.065 0.920 ;
        RECT 9.935 0.845 10.225 0.920 ;
    END
  END C
  PIN VGND
    ANTENNADIFFAREA 1.124200 ;
    PORT
      LAYER met1 ;
        RECT 3.215 0.440 3.505 0.730 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 0.000 -0.240 11.520 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 11.520 3.570 ;
        RECT 3.215 2.735 3.505 3.090 ;
        RECT 6.095 2.735 6.385 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 11.520 3.415 ;
        RECT 0.155 3.215 11.365 3.245 ;
        RECT 0.155 3.090 5.905 3.215 ;
        RECT 6.575 3.090 11.365 3.215 ;
        RECT 3.195 2.715 3.525 3.090 ;
      LAYER mcon ;
        RECT 6.155 3.245 6.325 3.415 ;
        RECT 3.275 2.795 3.445 2.965 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 11.520 3.330 ;
      LAYER li1 ;
        RECT 6.075 2.715 6.405 3.045 ;
        RECT 0.555 2.175 0.885 2.505 ;
        RECT 5.115 2.260 5.445 2.505 ;
        RECT 5.115 2.175 5.425 2.260 ;
        RECT 7.755 2.175 8.085 2.505 ;
        RECT 9.195 2.175 9.525 2.505 ;
        RECT 10.395 2.260 10.725 2.505 ;
        RECT 10.415 2.175 10.725 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 2.795 1.155 2.965 1.760 ;
        RECT 4.235 1.155 4.405 1.760 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 2.715 0.920 3.045 1.155 ;
        RECT 2.715 0.825 3.025 0.920 ;
        RECT 4.155 0.825 4.485 1.155 ;
        RECT 5.595 0.920 5.925 1.155 ;
        RECT 5.595 0.825 5.905 0.920 ;
        RECT 7.035 0.825 7.365 1.155 ;
        RECT 7.835 0.750 8.005 2.175 ;
        RECT 9.915 1.760 10.245 2.090 ;
        RECT 9.995 1.155 10.165 1.760 ;
        RECT 9.915 0.825 10.245 1.155 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 3.195 0.420 3.525 0.750 ;
        RECT 5.115 0.655 5.425 0.750 ;
        RECT 5.115 0.420 5.445 0.655 ;
        RECT 6.075 0.420 6.405 0.750 ;
        RECT 7.755 0.420 8.085 0.750 ;
        RECT 9.195 0.420 9.525 0.750 ;
        RECT 10.415 0.655 10.725 0.750 ;
        RECT 10.395 0.420 10.725 0.655 ;
        RECT 6.155 0.240 6.325 0.420 ;
        RECT 0.155 0.085 11.365 0.240 ;
        RECT 0.000 -0.085 11.520 0.085 ;
      LAYER mcon ;
        RECT 6.155 2.795 6.325 2.965 ;
        RECT 0.635 2.255 0.805 2.425 ;
        RECT 5.195 2.255 5.365 2.425 ;
        RECT 9.275 2.255 9.445 2.425 ;
        RECT 10.475 2.255 10.645 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 5.675 1.840 5.845 2.010 ;
        RECT 7.115 1.840 7.285 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 7.115 0.905 7.285 1.075 ;
        RECT 7.835 0.905 8.005 1.075 ;
        RECT 9.995 0.905 10.165 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 5.195 0.500 5.365 0.670 ;
        RECT 9.275 0.500 9.445 0.670 ;
        RECT 10.475 0.500 10.645 0.670 ;
        RECT 3.275 -0.085 3.445 0.085 ;
      LAYER met1 ;
        RECT 0.575 2.195 0.865 2.485 ;
        RECT 5.135 2.410 5.425 2.485 ;
        RECT 9.215 2.410 9.505 2.485 ;
        RECT 5.135 2.270 9.505 2.410 ;
        RECT 5.135 2.195 5.425 2.270 ;
        RECT 9.215 2.195 9.505 2.270 ;
        RECT 10.415 2.195 10.705 2.485 ;
        RECT 0.650 0.730 0.790 2.195 ;
        RECT 7.055 1.995 7.345 2.070 ;
        RECT 10.490 1.995 10.630 2.195 ;
        RECT 7.055 1.855 10.630 1.995 ;
        RECT 7.055 1.780 7.345 1.855 ;
        RECT 7.130 1.135 7.270 1.780 ;
        RECT 7.055 0.845 7.345 1.135 ;
        RECT 10.490 0.730 10.630 1.855 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 5.135 0.655 5.425 0.730 ;
        RECT 9.215 0.655 9.505 0.730 ;
        RECT 5.135 0.515 9.505 0.655 ;
        RECT 5.135 0.440 5.425 0.515 ;
        RECT 9.215 0.440 9.505 0.515 ;
        RECT 10.415 0.440 10.705 0.730 ;
  END
END SUTHERLAND1989
END LIBRARY

