VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 1.780 3.060 2.070 3.090 ;
        RECT 1.780 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.070 3.060 ;
        RECT 1.780 2.830 2.070 2.890 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.360 2.070 0.420 ;
        RECT 1.780 0.240 1.840 0.360 ;
        RECT 2.010 0.240 2.070 0.360 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.370 0.870 2.440 ;
        RECT 3.220 2.370 3.510 2.440 ;
        RECT 0.580 2.230 3.510 2.370 ;
        RECT 0.580 2.150 0.870 2.230 ;
        RECT 3.220 2.150 3.510 2.230 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 3.290 0.690 3.430 2.150 ;
        RECT 0.580 0.400 0.870 0.690 ;
        RECT 3.220 0.400 3.510 0.690 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 2.740 1.750 3.030 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 1.300 1.020 1.590 1.090 ;
        RECT 2.740 1.020 3.030 1.090 ;
        RECT 1.300 0.880 3.030 1.020 ;
        RECT 1.300 0.800 1.590 0.880 ;
        RECT 2.740 0.800 3.030 0.880 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 3.060 2.090 3.140 ;
        RECT 1.760 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.090 3.060 ;
        RECT 1.760 2.810 2.090 2.890 ;
        RECT 0.560 2.380 0.890 2.460 ;
        RECT 0.560 2.210 0.640 2.380 ;
        RECT 0.810 2.210 0.890 2.380 ;
        RECT 0.560 2.130 0.890 2.210 ;
        RECT 3.200 2.380 3.530 2.460 ;
        RECT 3.200 2.210 3.280 2.380 ;
        RECT 3.450 2.210 3.530 2.380 ;
        RECT 3.200 2.130 3.530 2.210 ;
        RECT 1.280 1.980 1.610 2.060 ;
        RECT 1.280 1.810 1.360 1.980 ;
        RECT 1.530 1.810 1.610 1.980 ;
        RECT 1.280 1.730 1.610 1.810 ;
        RECT 2.720 1.980 3.030 2.060 ;
        RECT 2.720 1.810 2.800 1.980 ;
        RECT 2.970 1.960 3.030 1.980 ;
        RECT 2.970 1.810 3.050 1.960 ;
        RECT 2.720 1.730 3.050 1.810 ;
        RECT 1.280 1.030 1.610 1.110 ;
        RECT 1.280 0.860 1.360 1.030 ;
        RECT 1.530 0.860 1.610 1.030 ;
        RECT 1.280 0.780 1.610 0.860 ;
        RECT 2.720 1.030 3.050 1.110 ;
        RECT 2.720 0.860 2.800 1.030 ;
        RECT 2.970 0.880 3.050 1.030 ;
        RECT 2.970 0.860 3.030 0.880 ;
        RECT 2.720 0.780 3.030 0.860 ;
        RECT 0.560 0.630 0.890 0.710 ;
        RECT 0.560 0.460 0.640 0.630 ;
        RECT 0.810 0.460 0.890 0.630 ;
        RECT 0.560 0.380 0.890 0.460 ;
        RECT 3.200 0.630 3.530 0.710 ;
        RECT 3.200 0.460 3.280 0.630 ;
        RECT 3.450 0.460 3.530 0.630 ;
        RECT 1.760 0.360 2.090 0.440 ;
        RECT 3.200 0.380 3.530 0.460 ;
        RECT 1.760 0.190 1.840 0.360 ;
        RECT 2.010 0.190 2.090 0.360 ;
        RECT 1.760 0.110 2.090 0.190 ;
  END
END INVX4
END LIBRARY

