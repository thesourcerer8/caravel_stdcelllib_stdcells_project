VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 12.960 3.570 ;
        RECT 0.580 2.990 0.870 3.090 ;
        RECT 0.580 2.820 0.640 2.990 ;
        RECT 0.810 2.820 0.870 2.990 ;
        RECT 0.580 2.760 0.870 2.820 ;
        RECT 3.220 2.990 3.510 3.090 ;
        RECT 3.220 2.820 3.280 2.990 ;
        RECT 3.450 2.820 3.510 2.990 ;
        RECT 3.220 2.760 3.510 2.820 ;
        RECT 6.100 2.990 6.390 3.090 ;
        RECT 6.100 2.820 6.160 2.990 ;
        RECT 6.330 2.820 6.390 2.990 ;
        RECT 6.100 2.760 6.390 2.820 ;
        RECT 8.980 2.990 9.270 3.090 ;
        RECT 8.980 2.820 9.040 2.990 ;
        RECT 9.210 2.820 9.270 2.990 ;
        RECT 8.980 2.760 9.270 2.820 ;
        RECT 11.860 2.990 12.150 3.090 ;
        RECT 11.860 2.820 11.920 2.990 ;
        RECT 12.090 2.820 12.150 2.990 ;
        RECT 11.860 2.760 12.150 2.820 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 12.960 3.570 ;
        RECT 0.560 2.990 0.890 3.090 ;
        RECT 0.560 2.820 0.640 2.990 ;
        RECT 0.810 2.820 0.890 2.990 ;
        RECT 0.560 2.740 0.890 2.820 ;
        RECT 3.200 2.990 3.530 3.090 ;
        RECT 3.200 2.820 3.280 2.990 ;
        RECT 3.450 2.820 3.530 2.990 ;
        RECT 3.200 2.740 3.530 2.820 ;
        RECT 6.080 2.990 6.410 3.090 ;
        RECT 6.080 2.820 6.160 2.990 ;
        RECT 6.330 2.820 6.410 2.990 ;
        RECT 6.080 2.740 6.410 2.820 ;
        RECT 8.960 2.990 9.290 3.090 ;
        RECT 8.960 2.820 9.040 2.990 ;
        RECT 9.210 2.820 9.290 2.990 ;
        RECT 8.960 2.740 9.290 2.820 ;
        RECT 11.840 2.990 12.170 3.090 ;
        RECT 11.840 2.820 11.920 2.990 ;
        RECT 12.090 2.820 12.170 2.990 ;
        RECT 11.840 2.740 12.170 2.820 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 0.510 0.870 0.570 ;
        RECT 0.580 0.340 0.640 0.510 ;
        RECT 0.810 0.340 0.870 0.510 ;
        RECT 0.580 0.240 0.870 0.340 ;
        RECT 3.220 0.510 3.510 0.570 ;
        RECT 3.220 0.340 3.280 0.510 ;
        RECT 3.450 0.340 3.510 0.510 ;
        RECT 3.220 0.240 3.510 0.340 ;
        RECT 6.100 0.510 6.390 0.570 ;
        RECT 6.100 0.340 6.160 0.510 ;
        RECT 6.330 0.340 6.390 0.510 ;
        RECT 6.100 0.240 6.390 0.340 ;
        RECT 8.980 0.510 9.270 0.570 ;
        RECT 8.980 0.340 9.040 0.510 ;
        RECT 9.210 0.340 9.270 0.510 ;
        RECT 8.980 0.240 9.270 0.340 ;
        RECT 11.860 0.510 12.150 0.570 ;
        RECT 11.860 0.340 11.920 0.510 ;
        RECT 12.090 0.340 12.150 0.510 ;
        RECT 11.860 0.240 12.150 0.340 ;
        RECT 0.000 -0.240 12.960 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.560 0.510 0.890 0.590 ;
        RECT 0.560 0.340 0.640 0.510 ;
        RECT 0.810 0.340 0.890 0.510 ;
        RECT 0.560 0.240 0.890 0.340 ;
        RECT 3.200 0.510 3.530 0.590 ;
        RECT 3.200 0.340 3.280 0.510 ;
        RECT 3.450 0.340 3.530 0.510 ;
        RECT 3.200 0.240 3.530 0.340 ;
        RECT 6.080 0.510 6.410 0.590 ;
        RECT 6.080 0.340 6.160 0.510 ;
        RECT 6.330 0.340 6.410 0.510 ;
        RECT 6.080 0.240 6.410 0.340 ;
        RECT 8.960 0.510 9.290 0.590 ;
        RECT 8.960 0.340 9.040 0.510 ;
        RECT 9.210 0.340 9.290 0.510 ;
        RECT 8.960 0.240 9.290 0.340 ;
        RECT 11.840 0.510 12.170 0.590 ;
        RECT 11.840 0.340 11.920 0.510 ;
        RECT 12.090 0.340 12.170 0.510 ;
        RECT 11.840 0.240 12.170 0.340 ;
        RECT 0.000 -0.240 12.960 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 10.420 0.440 10.710 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.370 2.680 2.950 2.820 ;
        RECT 1.370 2.070 1.510 2.680 ;
        RECT 2.810 2.070 2.950 2.680 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 2.810 1.540 2.950 1.780 ;
        RECT 2.740 1.250 3.030 1.540 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 2.430 2.090 2.510 ;
        RECT 1.760 2.260 1.840 2.430 ;
        RECT 2.010 2.260 2.090 2.430 ;
        RECT 4.640 2.430 4.970 2.510 ;
        RECT 4.640 2.260 4.720 2.430 ;
        RECT 4.890 2.260 4.970 2.430 ;
        RECT 1.780 2.180 2.090 2.260 ;
        RECT 4.660 2.180 4.970 2.260 ;
        RECT 5.680 2.090 5.850 2.660 ;
        RECT 7.520 2.430 7.850 2.510 ;
        RECT 7.520 2.260 7.600 2.430 ;
        RECT 7.770 2.260 7.850 2.430 ;
        RECT 7.520 2.180 7.850 2.260 ;
        RECT 8.560 2.090 8.730 2.660 ;
        RECT 10.400 2.430 10.730 2.510 ;
        RECT 10.400 2.260 10.480 2.430 ;
        RECT 10.650 2.260 10.730 2.430 ;
        RECT 10.420 2.180 10.730 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 2.010 5.930 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 7.040 2.010 7.350 2.090 ;
        RECT 8.480 2.010 8.810 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 8.480 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.810 2.010 ;
        RECT 8.480 1.760 8.810 1.840 ;
        RECT 9.920 2.010 10.250 2.090 ;
        RECT 9.920 1.840 10.000 2.010 ;
        RECT 10.170 1.840 10.250 2.010 ;
        RECT 9.920 1.760 10.250 1.840 ;
        RECT 5.680 1.620 5.850 1.760 ;
        RECT 8.560 1.620 8.730 1.760 ;
        RECT 2.800 1.160 2.970 1.310 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.920 4.490 1.080 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 4.410 0.910 4.470 0.920 ;
        RECT 4.160 0.830 4.470 0.910 ;
        RECT 5.600 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.600 0.830 5.930 0.910 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.920 7.370 1.080 ;
        RECT 8.480 1.080 8.810 1.160 ;
        RECT 7.290 0.910 7.350 0.920 ;
        RECT 7.040 0.830 7.350 0.910 ;
        RECT 8.480 0.910 8.560 1.080 ;
        RECT 8.730 0.910 8.810 1.080 ;
        RECT 8.480 0.830 8.810 0.910 ;
        RECT 9.920 1.080 10.250 1.160 ;
        RECT 9.920 0.910 10.000 1.080 ;
        RECT 10.170 0.920 10.250 1.080 ;
        RECT 10.170 0.910 10.230 0.920 ;
        RECT 9.920 0.830 10.230 0.910 ;
        RECT 10.480 0.750 10.650 2.180 ;
        RECT 11.360 2.010 11.690 2.090 ;
        RECT 11.360 1.840 11.440 2.010 ;
        RECT 11.610 1.840 11.690 2.010 ;
        RECT 11.360 1.760 11.690 1.840 ;
        RECT 11.360 1.080 11.690 1.160 ;
        RECT 11.360 0.910 11.440 1.080 ;
        RECT 11.610 0.910 11.690 1.080 ;
        RECT 11.360 0.830 11.690 0.910 ;
        RECT 1.780 0.670 2.090 0.750 ;
        RECT 1.780 0.660 1.840 0.670 ;
        RECT 1.760 0.500 1.840 0.660 ;
        RECT 2.010 0.500 2.090 0.670 ;
        RECT 1.760 0.420 2.090 0.500 ;
        RECT 4.640 0.670 4.970 0.750 ;
        RECT 4.640 0.500 4.720 0.670 ;
        RECT 4.890 0.500 4.970 0.670 ;
        RECT 4.640 0.420 4.970 0.500 ;
        RECT 7.520 0.670 7.850 0.750 ;
        RECT 7.520 0.500 7.600 0.670 ;
        RECT 7.770 0.500 7.850 0.670 ;
        RECT 7.520 0.420 7.850 0.500 ;
        RECT 10.400 0.670 10.730 0.750 ;
        RECT 10.400 0.500 10.480 0.670 ;
        RECT 10.650 0.500 10.730 0.670 ;
        RECT 10.400 0.420 10.730 0.500 ;
      LAYER met1 ;
        RECT 5.620 2.830 5.910 2.890 ;
        RECT 5.620 2.820 5.680 2.830 ;
        RECT 4.250 2.680 5.680 2.820 ;
        RECT 1.780 2.430 2.070 2.490 ;
        RECT 1.780 2.260 1.840 2.430 ;
        RECT 2.010 2.260 2.070 2.430 ;
        RECT 1.780 2.200 2.070 2.260 ;
        RECT 1.850 1.060 1.990 2.200 ;
        RECT 4.250 2.070 4.390 2.680 ;
        RECT 5.620 2.660 5.680 2.680 ;
        RECT 5.850 2.660 5.910 2.830 ;
        RECT 8.500 2.830 8.790 2.890 ;
        RECT 8.500 2.820 8.560 2.830 ;
        RECT 5.620 2.600 5.910 2.660 ;
        RECT 7.130 2.680 8.560 2.820 ;
        RECT 4.660 2.430 4.950 2.490 ;
        RECT 4.660 2.260 4.720 2.430 ;
        RECT 4.890 2.260 4.950 2.430 ;
        RECT 4.660 2.200 4.950 2.260 ;
        RECT 4.180 2.010 4.470 2.070 ;
        RECT 4.180 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.470 2.010 ;
        RECT 4.180 1.780 4.470 1.840 ;
        RECT 4.730 2.000 4.870 2.200 ;
        RECT 7.130 2.070 7.270 2.680 ;
        RECT 8.500 2.660 8.560 2.680 ;
        RECT 8.730 2.660 8.790 2.830 ;
        RECT 8.500 2.600 8.790 2.660 ;
        RECT 7.540 2.430 7.830 2.490 ;
        RECT 7.540 2.260 7.600 2.430 ;
        RECT 7.770 2.260 7.830 2.430 ;
        RECT 7.540 2.200 7.830 2.260 ;
        RECT 7.060 2.010 7.350 2.070 ;
        RECT 7.060 2.000 7.120 2.010 ;
        RECT 4.730 1.860 7.120 2.000 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 4.180 1.080 4.470 1.140 ;
        RECT 4.180 1.060 4.240 1.080 ;
        RECT 1.850 0.920 4.240 1.060 ;
        RECT 1.850 0.730 1.990 0.920 ;
        RECT 4.180 0.910 4.240 0.920 ;
        RECT 4.410 0.910 4.470 1.080 ;
        RECT 4.180 0.850 4.470 0.910 ;
        RECT 4.730 0.730 4.870 1.860 ;
        RECT 7.060 1.840 7.120 1.860 ;
        RECT 7.290 1.840 7.350 2.010 ;
        RECT 7.060 1.780 7.350 1.840 ;
        RECT 7.610 2.000 7.750 2.200 ;
        RECT 9.940 2.010 10.230 2.070 ;
        RECT 9.940 2.000 10.000 2.010 ;
        RECT 7.610 1.860 10.000 2.000 ;
        RECT 5.620 1.620 5.910 1.680 ;
        RECT 5.620 1.450 5.680 1.620 ;
        RECT 5.850 1.450 5.910 1.620 ;
        RECT 5.620 1.390 5.910 1.450 ;
        RECT 5.690 1.140 5.830 1.390 ;
        RECT 7.130 1.140 7.270 1.780 ;
        RECT 5.620 1.080 5.910 1.140 ;
        RECT 5.620 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.910 1.080 ;
        RECT 5.620 0.850 5.910 0.910 ;
        RECT 7.060 1.080 7.350 1.140 ;
        RECT 7.060 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.350 1.080 ;
        RECT 7.060 0.850 7.350 0.910 ;
        RECT 7.610 0.730 7.750 1.860 ;
        RECT 9.940 1.840 10.000 1.860 ;
        RECT 10.170 2.000 10.230 2.010 ;
        RECT 11.380 2.010 11.670 2.070 ;
        RECT 11.380 2.000 11.440 2.010 ;
        RECT 10.170 1.860 11.440 2.000 ;
        RECT 10.170 1.840 10.230 1.860 ;
        RECT 9.940 1.780 10.230 1.840 ;
        RECT 11.380 1.840 11.440 1.860 ;
        RECT 11.610 1.840 11.670 2.010 ;
        RECT 11.380 1.780 11.670 1.840 ;
        RECT 8.500 1.620 8.790 1.680 ;
        RECT 8.500 1.450 8.560 1.620 ;
        RECT 8.730 1.450 8.790 1.620 ;
        RECT 8.500 1.390 8.790 1.450 ;
        RECT 8.570 1.140 8.710 1.390 ;
        RECT 10.010 1.140 10.150 1.780 ;
        RECT 11.450 1.140 11.590 1.780 ;
        RECT 8.500 1.080 8.790 1.140 ;
        RECT 8.500 0.910 8.560 1.080 ;
        RECT 8.730 0.910 8.790 1.080 ;
        RECT 8.500 0.850 8.790 0.910 ;
        RECT 9.940 1.080 10.230 1.140 ;
        RECT 9.940 0.910 10.000 1.080 ;
        RECT 10.170 0.910 10.230 1.080 ;
        RECT 9.940 0.850 10.230 0.910 ;
        RECT 11.380 1.080 11.670 1.140 ;
        RECT 11.380 0.910 11.440 1.080 ;
        RECT 11.610 0.910 11.670 1.080 ;
        RECT 11.380 0.850 11.670 0.910 ;
        RECT 1.780 0.670 2.070 0.730 ;
        RECT 1.780 0.500 1.840 0.670 ;
        RECT 2.010 0.500 2.070 0.670 ;
        RECT 1.780 0.440 2.070 0.500 ;
        RECT 4.660 0.670 4.950 0.730 ;
        RECT 4.660 0.500 4.720 0.670 ;
        RECT 4.890 0.500 4.950 0.670 ;
        RECT 4.660 0.440 4.950 0.500 ;
        RECT 7.540 0.670 7.830 0.730 ;
        RECT 7.540 0.500 7.600 0.670 ;
        RECT 7.770 0.500 7.830 0.670 ;
        RECT 7.540 0.440 7.830 0.500 ;
  END
END CLKBUF1
END LIBRARY

