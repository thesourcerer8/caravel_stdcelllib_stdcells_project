magic
tech sky130A
timestamp 1624575626
<< nwell >>
rect 0 179 1008 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
rect 713 24 728 66
rect 857 24 872 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
rect 713 225 728 309
rect 857 225 872 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 466 67 495 73
rect 466 66 472 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 51 281 66
rect 152 34 184 51
rect 201 34 281 51
rect 152 24 281 34
rect 296 24 425 66
rect 440 50 472 66
rect 489 66 495 67
rect 898 67 927 73
rect 898 66 904 67
rect 489 50 569 66
rect 440 24 569 50
rect 584 24 713 66
rect 728 51 857 66
rect 728 34 760 51
rect 777 34 857 51
rect 728 24 857 34
rect 872 50 904 66
rect 921 66 927 67
rect 921 50 951 66
rect 872 24 951 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 299 281 309
rect 152 282 184 299
rect 201 282 281 299
rect 152 225 281 282
rect 296 225 425 309
rect 440 243 569 309
rect 440 226 472 243
rect 489 226 569 243
rect 440 225 569 226
rect 584 225 713 309
rect 728 299 857 309
rect 728 282 760 299
rect 777 282 857 299
rect 728 225 857 282
rect 872 243 951 309
rect 872 226 904 243
rect 921 226 951 243
rect 872 225 951 226
rect 58 220 87 225
rect 466 220 495 225
rect 898 220 927 225
<< ndiffc >>
rect 64 50 81 67
rect 184 34 201 51
rect 472 50 489 67
rect 760 34 777 51
rect 904 50 921 67
<< pdiffc >>
rect 64 226 81 243
rect 184 282 201 299
rect 472 226 489 243
rect 760 282 777 299
rect 904 226 921 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 713 309 728 322
rect 857 309 872 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 713 209 728 225
rect 857 209 872 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 848 201 881 209
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 848 108 881 116
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 713 66 728 83
rect 857 66 872 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
rect 713 11 728 24
rect 857 11 872 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 712 184 729 201
rect 856 184 873 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
rect 712 91 729 108
rect 856 91 873 108
<< locali >>
rect 0 342 1008 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 736 342
rect 753 325 784 342
rect 801 325 832 342
rect 849 325 880 342
rect 897 325 928 342
rect 945 325 976 342
rect 993 325 1008 342
rect 0 309 1008 325
rect 176 299 209 309
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 752 299 785 309
rect 752 282 760 299
rect 777 282 785 299
rect 752 274 785 282
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 464 243 497 251
rect 464 226 472 243
rect 489 226 497 243
rect 896 243 929 251
rect 896 226 904 243
rect 921 226 929 243
rect 56 218 89 226
rect 466 218 497 226
rect 898 218 929 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 136 116 153 176
rect 280 116 297 176
rect 424 116 441 131
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 92 449 108
rect 441 91 447 92
rect 416 83 447 91
rect 472 75 489 218
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 848 201 881 209
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 520 108 537 172
rect 560 108 593 116
rect 520 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 848 108 881 116
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 464 67 497 75
rect 56 42 89 50
rect 176 51 209 59
rect 176 34 184 51
rect 201 34 209 51
rect 464 50 472 67
rect 489 50 497 67
rect 568 67 585 83
rect 898 67 929 75
rect 898 66 904 67
rect 752 51 785 59
rect 464 42 497 50
rect 176 26 209 34
rect 752 34 760 51
rect 777 34 785 51
rect 896 50 904 66
rect 921 50 929 67
rect 896 42 929 50
rect 159 24 226 26
rect 752 24 785 34
rect 0 9 1008 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 736 9
rect 753 -9 784 9
rect 801 -9 832 9
rect 849 -9 880 9
rect 897 -9 928 9
rect 945 -9 976 9
rect 993 -9 1008 9
rect 0 -24 1008 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 304 325 321 342
rect 352 325 369 342
rect 400 325 417 342
rect 448 325 465 342
rect 496 325 513 342
rect 544 325 561 342
rect 592 325 609 342
rect 640 325 657 342
rect 688 325 705 342
rect 736 325 753 342
rect 784 325 801 342
rect 832 325 849 342
rect 880 325 897 342
rect 928 325 945 342
rect 976 325 993 342
rect 184 282 201 299
rect 760 282 777 299
rect 64 226 81 243
rect 904 226 921 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 424 131 441 148
rect 520 172 537 189
rect 568 184 585 201
rect 712 184 729 201
rect 856 184 873 201
rect 712 91 729 108
rect 856 91 873 108
rect 64 50 81 67
rect 184 34 201 51
rect 472 50 489 67
rect 568 50 585 67
rect 904 50 921 67
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
rect 304 -9 321 9
rect 352 -9 369 9
rect 400 -9 417 9
rect 448 -9 465 9
rect 496 -9 513 9
rect 544 -9 561 9
rect 592 -9 609 9
rect 640 -9 657 9
rect 688 -9 705 9
rect 736 -9 753 9
rect 784 -9 801 9
rect 832 -9 849 9
rect 880 -9 897 9
rect 928 -9 945 9
rect 976 -9 993 9
<< metal1 >>
rect 0 342 1008 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 736 342
rect 753 325 784 342
rect 801 325 832 342
rect 849 325 880 342
rect 897 325 928 342
rect 945 325 976 342
rect 993 325 1008 342
rect 0 309 1008 325
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 754 299 783 309
rect 754 282 760 299
rect 777 282 783 299
rect 754 276 783 282
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 898 243 927 249
rect 898 241 904 243
rect 58 220 87 226
rect 569 227 904 241
rect 65 106 79 220
rect 569 207 583 227
rect 898 226 904 227
rect 921 226 927 243
rect 898 220 927 226
rect 130 201 159 207
rect 130 184 136 201
rect 153 200 159 201
rect 274 201 303 207
rect 274 200 280 201
rect 153 186 280 200
rect 153 184 159 186
rect 130 178 159 184
rect 274 184 280 186
rect 297 184 303 201
rect 274 178 303 184
rect 418 201 447 207
rect 418 184 424 201
rect 441 187 447 201
rect 562 201 591 207
rect 514 189 543 195
rect 514 187 520 189
rect 441 184 520 187
rect 418 178 520 184
rect 425 173 520 178
rect 514 172 520 173
rect 537 172 543 189
rect 562 184 568 201
rect 585 184 591 201
rect 562 178 591 184
rect 706 201 735 207
rect 706 184 712 201
rect 729 184 735 201
rect 706 178 735 184
rect 850 201 879 207
rect 850 184 856 201
rect 873 184 879 201
rect 850 178 879 184
rect 514 166 543 172
rect 418 148 447 154
rect 418 131 424 148
rect 441 147 447 148
rect 569 147 583 178
rect 441 133 583 147
rect 441 131 447 133
rect 418 125 447 131
rect 713 114 727 178
rect 857 114 871 178
rect 706 108 735 114
rect 706 106 712 108
rect 65 92 712 106
rect 65 73 79 92
rect 706 91 712 92
rect 729 91 735 108
rect 706 85 735 91
rect 850 108 879 114
rect 850 91 856 108
rect 873 91 879 108
rect 850 85 879 91
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 466 67 495 73
rect 58 44 87 50
rect 178 51 207 57
rect 178 34 184 51
rect 201 34 207 51
rect 466 50 472 67
rect 489 50 495 67
rect 466 44 495 50
rect 562 67 591 73
rect 562 50 568 67
rect 585 66 591 67
rect 857 66 871 85
rect 905 73 919 220
rect 585 52 871 66
rect 898 67 927 73
rect 585 50 591 52
rect 562 44 591 50
rect 898 50 904 67
rect 921 50 927 67
rect 898 44 927 50
rect 178 24 207 34
rect 0 9 1008 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 736 9
rect 753 -9 784 9
rect 801 -9 832 9
rect 849 -9 880 9
rect 897 -9 928 9
rect 945 -9 976 9
rect 993 -9 1008 9
rect 0 -24 1008 -9
<< labels >>
rlabel locali 0 309 1008 357 0 VDD
port 1 se
rlabel metal1 0 309 1008 357 0 VDD
port 2 se
rlabel locali 0 -24 1008 24 0 GND
port 3 se
rlabel metal1 0 -24 1008 24 0 GND
port 4 se
rlabel metal1 466 44 495 73 0 Y
port 5 se
rlabel metal1 130 178 159 186 0 B
port 6 se
rlabel metal1 274 178 303 186 0 B
port 7 se
rlabel metal1 130 186 303 200 0 B
port 8 se
rlabel metal1 130 200 159 207 0 B
port 9 se
rlabel metal1 274 200 303 207 0 B
port 10 se
rlabel metal1 514 166 543 173 0 A
port 11 se
rlabel metal1 425 173 543 178 0 A
port 12 se
rlabel metal1 418 178 543 187 0 A
port 13 se
rlabel metal1 514 187 543 195 0 A
port 14 se
rlabel metal1 418 187 447 207 0 A
port 15 se
<< properties >>
string FIXED_BBOX 0 0 1008 333
<< end >>
