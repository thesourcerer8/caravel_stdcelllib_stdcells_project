VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.150 4.950 2.440 ;
        RECT 4.730 2.040 4.870 2.150 ;
        RECT 4.660 1.750 4.950 2.040 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 8.500 1.750 8.790 2.040 ;
        RECT 8.570 1.090 8.710 1.750 ;
        RECT 8.500 0.800 8.790 1.090 ;
        RECT 3.700 0.610 3.990 0.690 ;
        RECT 5.620 0.610 5.910 0.690 ;
        RECT 8.570 0.610 8.710 0.800 ;
        RECT 3.700 0.470 8.710 0.610 ;
        RECT 3.700 0.400 3.990 0.470 ;
        RECT 5.620 0.400 5.910 0.470 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.960 1.590 2.040 ;
        RECT 2.740 1.960 3.030 2.040 ;
        RECT 1.300 1.820 3.030 1.960 ;
        RECT 1.300 1.750 1.590 1.820 ;
        RECT 2.740 1.750 3.030 1.820 ;
        RECT 1.370 1.500 1.510 1.750 ;
        RECT 1.300 1.210 1.590 1.500 ;
    END
  END B
END XNOR2X1
END LIBRARY

