magic
tech sky130A
magscale 1 2
timestamp 1636963008
<< obsli1 >>
rect 1152 2647 59873 57293
<< obsm1 >>
rect 208 2083 59888 57325
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1268 0 1324 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2612 0 2668 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3092 0 3148 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 3956 0 4012 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4436 0 4492 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4820 0 4876 800
rect 4916 0 4972 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5300 0 5356 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5780 0 5836 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6164 0 6220 800
rect 6260 0 6316 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6644 0 6700 800
rect 6740 0 6796 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7124 0 7180 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7508 0 7564 800
rect 7604 0 7660 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 7988 0 8044 800
rect 8084 0 8140 800
rect 8276 0 8332 800
rect 8372 0 8428 800
rect 8468 0 8524 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8852 0 8908 800
rect 8948 0 9004 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9332 0 9388 800
rect 9428 0 9484 800
rect 9620 0 9676 800
rect 9716 0 9772 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10100 0 10156 800
rect 10196 0 10252 800
rect 10292 0 10348 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10676 0 10732 800
rect 10772 0 10828 800
rect 10964 0 11020 800
rect 11060 0 11116 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11444 0 11500 800
rect 11540 0 11596 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11924 0 11980 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12308 0 12364 800
rect 12404 0 12460 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12788 0 12844 800
rect 12884 0 12940 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13268 0 13324 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13748 0 13804 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14132 0 14188 800
rect 14228 0 14284 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14612 0 14668 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 15092 0 15148 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15476 0 15532 800
rect 15572 0 15628 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15956 0 16012 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16436 0 16492 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17300 0 17356 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17780 0 17836 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19124 0 19180 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20372 0 20428 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21716 0 21772 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22196 0 22252 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23060 0 23116 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23540 0 23596 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 23924 0 23980 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24404 0 24460 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24884 0 24940 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25268 0 25324 800
rect 25364 0 25420 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25748 0 25804 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26228 0 26284 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26612 0 26668 800
rect 26708 0 26764 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27092 0 27148 800
rect 27188 0 27244 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27572 0 27628 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 27956 0 28012 800
rect 28052 0 28108 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28436 0 28492 800
rect 28532 0 28588 800
rect 28724 0 28780 800
rect 28820 0 28876 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29204 0 29260 800
rect 29300 0 29356 800
rect 29396 0 29452 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29780 0 29836 800
rect 29876 0 29932 800
rect 30068 0 30124 800
rect 30164 0 30220 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30548 0 30604 800
rect 30644 0 30700 800
rect 30740 0 30796 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31124 0 31180 800
rect 31220 0 31276 800
rect 31412 0 31468 800
rect 31508 0 31564 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31892 0 31948 800
rect 31988 0 32044 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32372 0 32428 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32756 0 32812 800
rect 32852 0 32908 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33236 0 33292 800
rect 33332 0 33388 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33716 0 33772 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34196 0 34252 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34580 0 34636 800
rect 34676 0 34732 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 35060 0 35116 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35540 0 35596 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36404 0 36460 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36884 0 36940 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37748 0 37804 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38228 0 38284 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39572 0 39628 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40820 0 40876 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42164 0 42220 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42644 0 42700 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43508 0 43564 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 43988 0 44044 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44372 0 44428 800
rect 44468 0 44524 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44852 0 44908 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45332 0 45388 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45716 0 45772 800
rect 45812 0 45868 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46196 0 46252 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46676 0 46732 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47060 0 47116 800
rect 47156 0 47212 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47540 0 47596 800
rect 47636 0 47692 800
rect 47828 0 47884 800
rect 47924 0 47980 800
rect 48020 0 48076 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48404 0 48460 800
rect 48500 0 48556 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48884 0 48940 800
rect 48980 0 49036 800
rect 49172 0 49228 800
rect 49268 0 49324 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49652 0 49708 800
rect 49748 0 49804 800
rect 49844 0 49900 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50228 0 50284 800
rect 50324 0 50380 800
rect 50516 0 50572 800
rect 50612 0 50668 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50996 0 51052 800
rect 51092 0 51148 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51476 0 51532 800
rect 51572 0 51628 800
rect 51668 0 51724 800
rect 51860 0 51916 800
rect 51956 0 52012 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52340 0 52396 800
rect 52436 0 52492 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52820 0 52876 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53204 0 53260 800
rect 53300 0 53356 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53684 0 53740 800
rect 53780 0 53836 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54164 0 54220 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54644 0 54700 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 55028 0 55084 800
rect 55124 0 55180 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55508 0 55564 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55988 0 56044 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56852 0 56908 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57332 0 57388 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58676 0 58732 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< obsm2 >>
rect 324 59144 636 59288
rect 804 59144 1116 59288
rect 1284 59144 1692 59288
rect 1860 59144 2172 59288
rect 2340 59144 2748 59288
rect 2916 59144 3228 59288
rect 3396 59144 3804 59288
rect 3972 59144 4284 59288
rect 4452 59144 4860 59288
rect 5028 59144 5340 59288
rect 5508 59144 5916 59288
rect 6084 59144 6396 59288
rect 6564 59144 6972 59288
rect 7140 59144 7452 59288
rect 7620 59144 8028 59288
rect 8196 59144 8508 59288
rect 8676 59144 9084 59288
rect 9252 59144 9564 59288
rect 9732 59144 10140 59288
rect 10308 59144 10620 59288
rect 10788 59144 11196 59288
rect 11364 59144 11676 59288
rect 11844 59144 12252 59288
rect 12420 59144 12732 59288
rect 12900 59144 13308 59288
rect 13476 59144 13788 59288
rect 13956 59144 14364 59288
rect 14532 59144 14844 59288
rect 15012 59144 15324 59288
rect 15492 59144 15900 59288
rect 16068 59144 16380 59288
rect 16548 59144 16956 59288
rect 17124 59144 17436 59288
rect 17604 59144 18012 59288
rect 18180 59144 18492 59288
rect 18660 59144 19068 59288
rect 19236 59144 19548 59288
rect 19716 59144 20124 59288
rect 20292 59144 20604 59288
rect 20772 59144 21180 59288
rect 21348 59144 21660 59288
rect 21828 59144 22236 59288
rect 22404 59144 22716 59288
rect 22884 59144 23292 59288
rect 23460 59144 23772 59288
rect 23940 59144 24348 59288
rect 24516 59144 24828 59288
rect 24996 59144 25404 59288
rect 25572 59144 25884 59288
rect 26052 59144 26460 59288
rect 26628 59144 26940 59288
rect 27108 59144 27516 59288
rect 27684 59144 27996 59288
rect 28164 59144 28572 59288
rect 28740 59144 29052 59288
rect 29220 59144 29628 59288
rect 29796 59144 30108 59288
rect 30276 59144 30588 59288
rect 30756 59144 31164 59288
rect 31332 59144 31644 59288
rect 31812 59144 32220 59288
rect 32388 59144 32700 59288
rect 32868 59144 33276 59288
rect 33444 59144 33756 59288
rect 33924 59144 34332 59288
rect 34500 59144 34812 59288
rect 34980 59144 35388 59288
rect 35556 59144 35868 59288
rect 36036 59144 36444 59288
rect 36612 59144 36924 59288
rect 37092 59144 37500 59288
rect 37668 59144 37980 59288
rect 38148 59144 38556 59288
rect 38724 59144 39036 59288
rect 39204 59144 39612 59288
rect 39780 59144 40092 59288
rect 40260 59144 40668 59288
rect 40836 59144 41148 59288
rect 41316 59144 41724 59288
rect 41892 59144 42204 59288
rect 42372 59144 42780 59288
rect 42948 59144 43260 59288
rect 43428 59144 43836 59288
rect 44004 59144 44316 59288
rect 44484 59144 44892 59288
rect 45060 59144 45372 59288
rect 45540 59144 45852 59288
rect 46020 59144 46428 59288
rect 46596 59144 46908 59288
rect 47076 59144 47484 59288
rect 47652 59144 47964 59288
rect 48132 59144 48540 59288
rect 48708 59144 49020 59288
rect 49188 59144 49596 59288
rect 49764 59144 50076 59288
rect 50244 59144 50652 59288
rect 50820 59144 51132 59288
rect 51300 59144 51708 59288
rect 51876 59144 52188 59288
rect 52356 59144 52764 59288
rect 52932 59144 53244 59288
rect 53412 59144 53820 59288
rect 53988 59144 54300 59288
rect 54468 59144 54876 59288
rect 55044 59144 55356 59288
rect 55524 59144 55932 59288
rect 56100 59144 56412 59288
rect 56580 59144 56988 59288
rect 57156 59144 57468 59288
rect 57636 59144 58044 59288
rect 58212 59144 58524 59288
rect 58692 59144 59100 59288
rect 59268 59144 59580 59288
rect 59748 59144 59882 59288
rect 214 856 59882 59144
rect 420 800 444 856
rect 900 800 924 856
rect 1380 800 1404 856
rect 1764 800 1788 856
rect 2244 800 2268 856
rect 2724 800 2748 856
rect 3204 800 3228 856
rect 3588 800 3612 856
rect 4068 800 4092 856
rect 4548 800 4572 856
rect 5028 800 5052 856
rect 5412 800 5436 856
rect 5892 800 5916 856
rect 6372 800 6396 856
rect 6852 800 6876 856
rect 7236 800 7260 856
rect 7716 800 7740 856
rect 8196 800 8220 856
rect 8580 800 8604 856
rect 9060 800 9084 856
rect 9540 800 9564 856
rect 10020 800 10044 856
rect 10404 800 10428 856
rect 10884 800 10908 856
rect 11364 800 11388 856
rect 11844 800 11868 856
rect 12228 800 12252 856
rect 12708 800 12732 856
rect 13188 800 13212 856
rect 13668 800 13692 856
rect 14052 800 14076 856
rect 14532 800 14556 856
rect 15012 800 15036 856
rect 15396 800 15420 856
rect 15876 800 15900 856
rect 16356 800 16380 856
rect 16836 800 16860 856
rect 17220 800 17244 856
rect 17700 800 17724 856
rect 18180 800 18204 856
rect 18660 800 18684 856
rect 19044 800 19068 856
rect 19524 800 19548 856
rect 20004 800 20028 856
rect 20484 800 20508 856
rect 20868 800 20892 856
rect 21348 800 21372 856
rect 21828 800 21852 856
rect 22308 800 22332 856
rect 22692 800 22716 856
rect 23172 800 23196 856
rect 23652 800 23676 856
rect 24036 800 24060 856
rect 24516 800 24540 856
rect 24996 800 25020 856
rect 25476 800 25500 856
rect 25860 800 25884 856
rect 26340 800 26364 856
rect 26820 800 26844 856
rect 27300 800 27324 856
rect 27684 800 27708 856
rect 28164 800 28188 856
rect 28644 800 28668 856
rect 29124 800 29148 856
rect 29508 800 29532 856
rect 29988 800 30012 856
rect 30468 800 30492 856
rect 30852 800 30876 856
rect 31332 800 31356 856
rect 31812 800 31836 856
rect 32292 800 32316 856
rect 32676 800 32700 856
rect 33156 800 33180 856
rect 33636 800 33660 856
rect 34116 800 34140 856
rect 34500 800 34524 856
rect 34980 800 35004 856
rect 35460 800 35484 856
rect 35940 800 35964 856
rect 36324 800 36348 856
rect 36804 800 36828 856
rect 37284 800 37308 856
rect 37668 800 37692 856
rect 38148 800 38172 856
rect 38628 800 38652 856
rect 39108 800 39132 856
rect 39492 800 39516 856
rect 39972 800 39996 856
rect 40452 800 40476 856
rect 40932 800 40956 856
rect 41316 800 41340 856
rect 41796 800 41820 856
rect 42276 800 42300 856
rect 42756 800 42780 856
rect 43140 800 43164 856
rect 43620 800 43644 856
rect 44100 800 44124 856
rect 44580 800 44604 856
rect 44964 800 44988 856
rect 45444 800 45468 856
rect 45924 800 45948 856
rect 46308 800 46332 856
rect 46788 800 46812 856
rect 47268 800 47292 856
rect 47748 800 47772 856
rect 48132 800 48156 856
rect 48612 800 48636 856
rect 49092 800 49116 856
rect 49572 800 49596 856
rect 49956 800 49980 856
rect 50436 800 50460 856
rect 50916 800 50940 856
rect 51396 800 51420 856
rect 51780 800 51804 856
rect 52260 800 52284 856
rect 52740 800 52764 856
rect 53124 800 53148 856
rect 53604 800 53628 856
rect 54084 800 54108 856
rect 54564 800 54588 856
rect 54948 800 54972 856
rect 55428 800 55452 856
rect 55908 800 55932 856
rect 56388 800 56412 856
rect 56772 800 56796 856
rect 57252 800 57276 856
rect 57732 800 57756 856
rect 58212 800 58236 856
rect 58596 800 58620 856
rect 59076 800 59100 856
rect 59556 800 59580 856
<< obsm3 >>
rect 2799 2631 50656 57309
<< metal4 >>
rect 4256 2616 4576 57324
rect 19616 2616 19936 57324
rect 34976 2616 35296 57324
rect 50336 2616 50656 57324
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 59636 0 59692 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 59732 0 59788 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 59828 0 59884 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 12884 0 12940 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 49748 0 49804 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 50132 0 50188 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 50516 0 50572 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 51572 0 51628 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 51956 0 52012 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 52340 0 52396 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 53780 0 53836 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 54164 0 54220 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 55988 0 56044 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 17300 0 17356 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 19124 0 19180 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 13268 0 13324 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 23060 0 23116 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 24884 0 24940 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 25268 0 25324 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 26708 0 26764 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 27092 0 27148 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 28532 0 28588 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 28916 0 28972 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 29300 0 29356 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 30356 0 30412 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 30740 0 30796 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 31124 0 31180 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 31508 0 31564 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 32180 0 32236 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 32564 0 32620 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 32948 0 33004 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 33332 0 33388 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 33716 0 33772 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 34004 0 34060 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 34388 0 34444 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 34772 0 34828 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 35156 0 35212 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 35540 0 35596 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 35828 0 35884 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 36212 0 36268 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 36596 0 36652 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 36980 0 37036 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 37364 0 37420 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 37748 0 37804 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 38036 0 38092 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 15092 0 15148 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 38420 0 38476 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 38804 0 38860 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 39188 0 39244 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 39572 0 39628 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 39860 0 39916 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 40244 0 40300 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 40628 0 40684 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 41012 0 41068 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 41396 0 41452 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 41684 0 41740 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 42068 0 42124 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 42452 0 42508 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 42836 0 42892 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 43220 0 43276 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 43508 0 43564 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 43892 0 43948 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 44276 0 44332 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 44660 0 44716 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 45044 0 45100 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 45332 0 45388 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 45716 0 45772 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 46100 0 46156 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 46484 0 46540 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 46868 0 46924 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 47540 0 47596 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 47924 0 47980 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 48308 0 48364 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 48692 0 48748 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 12980 0 13036 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 49460 0 49516 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 49844 0 49900 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 50228 0 50284 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 50612 0 50668 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 50996 0 51052 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 51284 0 51340 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 51668 0 51724 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 52052 0 52108 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 52436 0 52492 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 52820 0 52876 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 16628 0 16684 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 53204 0 53260 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 53492 0 53548 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 53876 0 53932 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 54260 0 54316 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 54644 0 54700 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 55028 0 55084 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 55316 0 55372 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 55700 0 55756 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 56084 0 56140 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 56468 0 56524 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 17012 0 17068 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 56852 0 56908 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 57140 0 57196 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 57524 0 57580 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 57908 0 57964 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 58292 0 58348 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 58676 0 58732 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 58964 0 59020 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 59348 0 59404 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 17396 0 17452 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 17780 0 17836 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 18068 0 18124 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 18452 0 18508 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 18836 0 18892 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 19220 0 19276 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 19604 0 19660 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 19892 0 19948 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 13364 0 13420 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 20276 0 20332 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 20660 0 20716 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 21044 0 21100 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 21428 0 21484 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 21716 0 21772 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 22100 0 22156 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 22484 0 22540 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 22868 0 22924 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 23252 0 23308 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 23540 0 23596 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 13748 0 13804 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 23924 0 23980 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 24308 0 24364 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 24692 0 24748 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 25076 0 25132 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 25364 0 25420 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 25748 0 25804 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 26132 0 26188 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 26516 0 26572 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 26900 0 26956 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 27188 0 27244 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 27572 0 27628 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 27956 0 28012 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 28340 0 28396 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 28724 0 28780 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 29012 0 29068 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 29396 0 29452 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 29780 0 29836 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 30164 0 30220 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 30548 0 30604 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 30932 0 30988 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 14420 0 14476 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 31220 0 31276 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 31604 0 31660 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 31988 0 32044 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 32372 0 32428 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 32756 0 32812 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 33044 0 33100 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 33428 0 33484 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 33812 0 33868 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 34196 0 34252 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 34580 0 34636 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 14804 0 14860 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 34868 0 34924 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 35252 0 35308 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 35636 0 35692 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 36020 0 36076 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 36404 0 36460 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 36692 0 36748 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 37076 0 37132 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 37460 0 37516 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 37844 0 37900 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 38228 0 38284 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 15188 0 15244 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 38516 0 38572 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 38900 0 38956 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 39284 0 39340 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 39668 0 39724 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 40052 0 40108 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 40340 0 40396 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 40724 0 40780 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 41108 0 41164 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 41492 0 41548 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 41876 0 41932 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 15572 0 15628 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 42164 0 42220 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 42548 0 42604 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 42932 0 42988 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 43316 0 43372 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 43700 0 43756 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 43988 0 44044 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 44372 0 44428 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 44756 0 44812 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 45140 0 45196 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 45524 0 45580 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 15956 0 16012 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 45812 0 45868 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 46196 0 46252 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 46580 0 46636 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 46964 0 47020 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 47348 0 47404 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 47636 0 47692 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 48020 0 48076 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 48404 0 48460 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 48788 0 48844 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 49172 0 49228 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 16244 0 16300 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 13076 0 13132 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 51092 0 51148 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 16724 0 16780 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 53300 0 53356 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 55124 0 55180 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 55508 0 55564 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 17108 0 17164 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 57332 0 57388 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 17492 0 17548 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 17876 0 17932 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 18260 0 18316 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 18548 0 18604 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 18932 0 18988 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 19316 0 19372 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 19700 0 19756 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 20084 0 20140 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 13460 0 13516 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 20372 0 20428 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 20756 0 20812 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 21140 0 21196 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 21524 0 21580 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 21908 0 21964 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 22196 0 22252 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 22580 0 22636 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 22964 0 23020 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 23348 0 23404 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 23732 0 23788 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 13844 0 13900 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 24116 0 24172 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 24404 0 24460 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 24788 0 24844 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 25172 0 25228 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 25556 0 25612 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 25940 0 25996 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 26228 0 26284 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 26612 0 26668 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 26996 0 27052 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 27380 0 27436 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 14228 0 14284 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 27764 0 27820 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 28436 0 28492 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 28820 0 28876 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 29204 0 29260 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 29588 0 29644 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 30644 0 30700 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 31028 0 31084 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 14612 0 14668 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 31412 0 31468 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 32852 0 32908 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 33236 0 33292 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 34676 0 34732 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 14900 0 14956 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 35060 0 35116 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 36884 0 36940 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 15284 0 15340 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 40820 0 40876 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 15668 0 15724 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 42644 0 42700 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 44852 0 44908 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 16052 0 16108 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 46676 0 46732 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 47060 0 47116 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 48884 0 48940 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 49268 0 49324 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 16436 0 16492 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 502 nsew power input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 502 nsew power input
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 503 nsew ground input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 4820 0 4876 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 6260 0 6316 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 6644 0 6700 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 8084 0 8140 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 8468 0 8524 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 8852 0 8908 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 9908 0 9964 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 10292 0 10348 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 10676 0 10732 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 11060 0 11116 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 11732 0 11788 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 12116 0 12172 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 12500 0 12556 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 2612 0 2668 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 4436 0 4492 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 5300 0 5356 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 7124 0 7180 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 7508 0 7564 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 1268 0 1324 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 9332 0 9388 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 9716 0 9772 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 11540 0 11596 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 11924 0 11980 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 3092 0 3148 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 5780 0 5836 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 6164 0 6220 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 7988 0 8044 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 8372 0 8428 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 10196 0 10252 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 12404 0 12460 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 3956 0 4012 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 60000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 1743156
string GDS_START 286082
<< end >>

