MACRO MUX2X1
 CLASS CORE ;
 FOREIGN MUX2X1 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 8.64000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 8.64000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 5.13500000 1.20500000 5.42500000 1.49500000 ;
        RECT 5.21000000 1.49500000 5.35000000 2.15000000 ;
        RECT 5.13500000 2.15000000 5.42500000 2.44000000 ;
    END
  END Y

  PIN S
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 4.25000000 0.47000000 6.31000000 0.61000000 ;
        RECT 4.25000000 0.61000000 4.39000000 0.80000000 ;
        RECT 1.29500000 0.80000000 1.58500000 0.87500000 ;
        RECT 4.17500000 0.80000000 4.46500000 0.87500000 ;
        RECT 1.29500000 0.87500000 4.46500000 1.01500000 ;
        RECT 1.29500000 1.01500000 1.58500000 1.09000000 ;
        RECT 4.17500000 1.01500000 4.46500000 1.09000000 ;
        RECT 5.61500000 1.74500000 5.90500000 1.82000000 ;
        RECT 6.17000000 0.61000000 6.31000000 1.82000000 ;
        RECT 5.61500000 1.82000000 6.31000000 1.96000000 ;
        RECT 5.61500000 1.96000000 5.90500000 2.03500000 ;
    END
  END S

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 7.05500000 0.80000000 7.34500000 1.09000000 ;
        RECT 7.13000000 1.09000000 7.27000000 1.74500000 ;
        RECT 7.05500000 1.74500000 7.34500000 2.03500000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.73500000 1.20500000 3.02500000 1.49500000 ;
    END
  END A


END MUX2X1
