VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.756000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.995 1.585 2.070 ;
        RECT 2.735 1.995 3.025 2.070 ;
        RECT 4.175 1.995 4.465 2.070 ;
        RECT 5.615 1.995 5.905 2.070 ;
        RECT 1.295 1.855 5.905 1.995 ;
        RECT 1.295 1.780 1.585 1.855 ;
        RECT 2.735 1.780 3.025 1.855 ;
        RECT 4.175 1.780 4.465 1.855 ;
        RECT 5.615 1.780 5.905 1.855 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 2.810 1.135 2.950 1.780 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 5.690 1.135 5.830 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
        RECT 2.735 0.845 3.025 1.135 ;
        RECT 4.175 0.845 4.465 1.135 ;
        RECT 5.615 0.845 5.905 1.135 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 1.124200 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 1.850 0.240 1.990 0.440 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 7.200 3.570 ;
        RECT 1.775 2.735 2.065 3.090 ;
        RECT 4.655 2.735 4.945 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.155 3.215 7.045 3.245 ;
        RECT 0.155 3.090 4.465 3.215 ;
        RECT 5.135 3.090 7.045 3.215 ;
        RECT 1.755 2.715 2.085 3.090 ;
      LAYER mcon ;
        RECT 1.835 3.245 2.005 3.415 ;
        RECT 1.835 2.795 2.005 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 3.724950 ;
    PORT
      LAYER met1 ;
        RECT 0.815 2.410 1.105 2.485 ;
        RECT 3.695 2.410 3.985 2.485 ;
        RECT 6.095 2.410 6.385 2.485 ;
        RECT 0.815 2.270 6.385 2.410 ;
        RECT 0.815 2.195 1.105 2.270 ;
        RECT 3.695 2.195 3.985 2.270 ;
        RECT 6.095 2.195 6.385 2.270 ;
        RECT 0.890 0.730 1.030 2.195 ;
        RECT 6.170 0.730 6.310 2.195 ;
        RECT 0.815 0.440 1.105 0.730 ;
        RECT 3.695 0.655 3.985 0.730 ;
        RECT 6.095 0.655 6.385 0.730 ;
        RECT 3.695 0.515 6.385 0.655 ;
        RECT 3.695 0.440 3.985 0.515 ;
        RECT 6.095 0.440 6.385 0.515 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 7.200 3.330 ;
      LAYER li1 ;
        RECT 4.635 2.715 4.965 3.045 ;
        RECT 0.795 2.175 1.125 2.505 ;
        RECT 3.675 2.260 4.005 2.505 ;
        RECT 6.075 2.260 6.405 2.505 ;
        RECT 3.675 2.175 3.985 2.260 ;
        RECT 6.095 2.175 6.405 2.260 ;
        RECT 1.295 2.005 1.605 2.090 ;
        RECT 1.275 1.760 1.605 2.005 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 5.595 0.920 5.925 1.155 ;
        RECT 4.175 0.825 4.465 0.920 ;
        RECT 5.595 0.825 5.905 0.920 ;
        RECT 0.795 0.655 1.105 0.750 ;
        RECT 0.795 0.420 1.125 0.655 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.675 0.420 4.005 0.750 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 6.075 0.420 6.405 0.750 ;
        RECT 4.715 0.240 4.885 0.420 ;
        RECT 0.155 0.085 7.045 0.240 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 4.715 2.795 4.885 2.965 ;
        RECT 0.875 2.255 1.045 2.425 ;
        RECT 3.755 2.255 3.925 2.425 ;
        RECT 6.155 2.255 6.325 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 5.675 1.840 5.845 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 0.875 0.500 1.045 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 3.755 0.500 3.925 0.670 ;
        RECT 6.155 0.500 6.325 0.670 ;
        RECT 4.715 -0.085 4.885 0.085 ;
  END
END INVX8
END LIBRARY

