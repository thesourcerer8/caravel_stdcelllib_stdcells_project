magic
tech sky130A
magscale 1 2
timestamp 1636962376
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 3168 666
<< nmos >>
rect 273 48 303 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1713 48 1743 132
rect 2001 48 2031 132
rect 2289 48 2319 132
rect 2865 48 2895 132
<< pmos >>
rect 273 450 303 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1713 450 1743 618
rect 2001 450 2031 618
rect 2289 450 2319 618
rect 2865 450 2895 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 355 134 413 146
rect 355 132 367 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 691 134 749 146
rect 401 100 461 132
rect 303 48 461 100
rect 691 100 703 134
rect 737 132 749 134
rect 1219 134 1277 146
rect 1219 132 1231 134
rect 737 100 849 132
rect 691 48 849 100
rect 879 48 1137 132
rect 1167 100 1231 132
rect 1265 132 1277 134
rect 1555 134 1613 146
rect 1265 100 1325 132
rect 1167 48 1325 100
rect 1555 100 1567 134
rect 1601 132 1613 134
rect 1891 134 1949 146
rect 1891 132 1903 134
rect 1601 100 1713 132
rect 1555 48 1713 100
rect 1743 100 1903 132
rect 1937 132 1949 134
rect 2083 134 2141 146
rect 2083 132 2095 134
rect 1937 100 2001 132
rect 1743 48 2001 100
rect 2031 100 2095 132
rect 2129 132 2141 134
rect 2371 134 2429 146
rect 2371 132 2383 134
rect 2129 100 2289 132
rect 2031 48 2289 100
rect 2319 100 2383 132
rect 2417 132 2429 134
rect 2707 134 2765 146
rect 2417 100 2477 132
rect 2319 48 2477 100
rect 2707 100 2719 134
rect 2753 132 2765 134
rect 2947 134 3005 146
rect 2947 132 2959 134
rect 2753 100 2865 132
rect 2707 48 2865 100
rect 2895 100 2959 132
rect 2993 132 3005 134
rect 2993 100 3053 132
rect 2895 48 3053 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 593 461 618
rect 303 559 367 593
rect 401 559 461 593
rect 303 450 461 559
rect 691 485 849 618
rect 691 451 703 485
rect 737 451 849 485
rect 691 450 849 451
rect 879 593 1137 618
rect 879 559 943 593
rect 977 559 1137 593
rect 879 450 1137 559
rect 1167 485 1325 618
rect 1167 451 1231 485
rect 1265 451 1325 485
rect 1167 450 1325 451
rect 1555 593 1713 618
rect 1555 559 1567 593
rect 1601 559 1713 593
rect 1555 450 1713 559
rect 1743 485 2001 618
rect 1743 451 1903 485
rect 1937 451 2001 485
rect 1743 450 2001 451
rect 2031 450 2289 618
rect 2319 593 2477 618
rect 2319 559 2383 593
rect 2417 559 2477 593
rect 2319 450 2477 559
rect 2707 593 2865 618
rect 2707 559 2719 593
rect 2753 559 2865 593
rect 2707 450 2865 559
rect 2895 485 3053 618
rect 2895 451 2959 485
rect 2993 451 3053 485
rect 2895 450 3053 451
rect 115 439 173 450
rect 691 439 749 450
rect 1219 439 1277 450
rect 1891 439 1949 450
rect 2947 439 3005 450
<< ndiffc >>
rect 127 100 161 134
rect 367 100 401 134
rect 703 100 737 134
rect 1231 100 1265 134
rect 1567 100 1601 134
rect 1903 100 1937 134
rect 2095 100 2129 134
rect 2383 100 2417 134
rect 2719 100 2753 134
rect 2959 100 2993 134
<< pdiffc >>
rect 127 451 161 485
rect 367 559 401 593
rect 703 451 737 485
rect 943 559 977 593
rect 1231 451 1265 485
rect 1567 559 1601 593
rect 1903 451 1937 485
rect 2383 559 2417 593
rect 2719 559 2753 593
rect 2959 451 2993 485
<< poly >>
rect 273 618 303 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1713 618 1743 644
rect 2001 618 2031 644
rect 2289 618 2319 644
rect 2865 618 2895 644
rect 273 418 303 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1713 418 1743 450
rect 2001 418 2031 450
rect 2289 418 2319 450
rect 2865 418 2895 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 2847 402 2913 418
rect 2847 368 2863 402
rect 2897 368 2913 402
rect 2847 352 2913 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 2271 215 2337 231
rect 2271 181 2287 215
rect 2321 181 2337 215
rect 2271 165 2337 181
rect 2847 215 2913 231
rect 2847 181 2863 215
rect 2897 181 2913 215
rect 2847 165 2913 181
rect 273 132 303 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1713 132 1743 165
rect 2001 132 2031 165
rect 2289 132 2319 165
rect 2865 132 2895 165
rect 273 22 303 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1713 22 1743 48
rect 2001 22 2031 48
rect 2289 22 2319 48
rect 2865 22 2895 48
<< polycont >>
rect 271 368 305 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 2287 368 2321 402
rect 2863 368 2897 402
rect 271 181 305 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 2287 181 2321 215
rect 2863 181 2897 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3168 683
rect 31 643 3137 649
rect 31 618 2333 643
rect 2467 618 3137 643
rect 351 593 417 618
rect 351 559 367 593
rect 401 559 417 593
rect 927 593 993 618
rect 351 543 417 559
rect 927 559 943 593
rect 977 559 993 593
rect 927 543 993 559
rect 1551 593 1617 618
rect 1551 559 1567 593
rect 1601 559 1617 593
rect 1551 543 1617 559
rect 2367 593 2433 609
rect 2367 559 2383 593
rect 2417 559 2433 593
rect 2367 543 2433 559
rect 2703 593 2769 618
rect 2703 559 2719 593
rect 2753 559 2769 593
rect 2703 543 2769 559
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 687 485 753 501
rect 687 451 703 485
rect 737 451 753 485
rect 687 435 753 451
rect 847 418 881 532
rect 1215 485 1281 501
rect 1215 452 1231 485
rect 1219 451 1231 452
rect 1265 451 1281 485
rect 1219 435 1281 451
rect 1887 485 1953 501
rect 1887 451 1903 485
rect 1937 452 1953 485
rect 2943 485 3009 501
rect 2943 452 2959 485
rect 1937 451 1949 452
rect 1887 435 1949 451
rect 2947 451 2959 452
rect 2993 451 3009 485
rect 2947 435 3009 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 2847 402 2913 418
rect 2847 368 2863 402
rect 2897 368 2913 402
rect 2847 352 2913 368
rect 1711 231 1745 352
rect 1999 231 2033 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 184 321 215
rect 831 215 897 231
rect 305 181 317 184
rect 255 165 317 181
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1983 215 2049 231
rect 1983 184 1999 215
rect 1695 165 1761 181
rect 1987 181 1999 184
rect 2033 184 2049 215
rect 2033 181 2045 184
rect 1987 165 2045 181
rect 2095 150 2129 262
rect 2271 215 2337 231
rect 2271 181 2287 215
rect 2321 184 2337 215
rect 2847 215 2913 231
rect 2321 181 2333 184
rect 2271 165 2333 181
rect 2847 181 2863 215
rect 2897 184 2913 215
rect 2897 181 2909 184
rect 2847 165 2909 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 351 134 417 150
rect 351 100 367 134
rect 401 100 417 134
rect 351 84 417 100
rect 687 134 753 150
rect 687 100 703 134
rect 737 100 753 134
rect 1219 134 1281 150
rect 1219 131 1231 134
rect 687 84 753 100
rect 1215 100 1231 131
rect 1265 100 1281 134
rect 1215 84 1281 100
rect 1551 134 1617 150
rect 1551 100 1567 134
rect 1601 100 1617 134
rect 1551 84 1617 100
rect 1887 134 1953 150
rect 1887 100 1903 134
rect 1937 100 1953 134
rect 1887 84 1953 100
rect 2079 134 2145 150
rect 2079 100 2095 134
rect 2129 100 2145 134
rect 2079 84 2145 100
rect 2367 134 2433 150
rect 2367 100 2383 134
rect 2417 100 2433 134
rect 2367 84 2433 100
rect 2703 134 2769 150
rect 2703 100 2719 134
rect 2753 100 2769 134
rect 2703 84 2769 100
rect 2943 134 3009 150
rect 2943 100 2959 134
rect 2993 100 3009 134
rect 2943 84 3009 100
rect 31 17 3137 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3168 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 367 559 401 593
rect 847 532 881 566
rect 2383 559 2417 593
rect 2719 559 2753 593
rect 127 451 161 485
rect 703 451 737 485
rect 1231 451 1265 485
rect 1903 451 1937 485
rect 2959 451 2993 485
rect 271 368 305 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 2287 368 2321 402
rect 2863 368 2897 402
rect 2095 262 2129 296
rect 271 181 305 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 2287 181 2321 215
rect 2863 181 2897 215
rect 127 100 161 134
rect 367 100 401 134
rect 703 100 737 134
rect 1231 100 1265 134
rect 1567 100 1601 134
rect 1903 100 1937 134
rect 2383 100 2417 134
rect 2719 100 2753 134
rect 2959 100 2993 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3168 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3168 683
rect 0 618 3168 649
rect 355 593 413 618
rect 355 559 367 593
rect 401 559 413 593
rect 2371 593 2429 618
rect 355 547 413 559
rect 835 566 893 578
rect 835 532 847 566
rect 881 563 893 566
rect 881 535 2030 563
rect 2371 559 2383 593
rect 2417 559 2429 593
rect 2371 547 2429 559
rect 2707 593 2765 618
rect 2707 559 2719 593
rect 2753 559 2765 593
rect 2707 547 2765 559
rect 881 532 893 535
rect 835 520 893 532
rect 115 485 173 497
rect 115 451 127 485
rect 161 451 173 485
rect 115 439 173 451
rect 691 485 749 497
rect 691 451 703 485
rect 737 482 749 485
rect 1219 485 1277 497
rect 1219 482 1231 485
rect 737 454 1231 482
rect 737 451 749 454
rect 691 439 749 451
rect 1219 451 1231 454
rect 1265 482 1277 485
rect 1891 485 1949 497
rect 1265 454 1742 482
rect 1265 451 1277 454
rect 1219 439 1277 451
rect 130 146 158 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 274 227 302 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 212 317 215
rect 706 212 734 439
rect 1714 414 1742 454
rect 1891 451 1903 485
rect 1937 451 1949 485
rect 1891 439 1949 451
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 1123 402 1181 414
rect 1123 368 1135 402
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 1699 402 1757 414
rect 1699 368 1711 402
rect 1745 368 1757 402
rect 1699 356 1757 368
rect 850 227 878 356
rect 1138 227 1166 356
rect 1906 293 1934 439
rect 2002 414 2030 535
rect 2947 485 3005 497
rect 2098 454 2894 482
rect 1987 402 2045 414
rect 1987 368 1999 402
rect 2033 368 2045 402
rect 1987 356 2045 368
rect 2098 308 2126 454
rect 2866 414 2894 454
rect 2947 451 2959 485
rect 2993 451 3005 485
rect 2947 439 3005 451
rect 2275 402 2333 414
rect 2275 368 2287 402
rect 2321 368 2333 402
rect 2275 356 2333 368
rect 2851 402 2909 414
rect 2851 368 2863 402
rect 2897 368 2909 402
rect 2851 356 2909 368
rect 2083 296 2141 308
rect 2083 293 2095 296
rect 1906 265 2095 293
rect 2083 262 2095 265
rect 2129 262 2141 296
rect 2083 250 2141 262
rect 2290 227 2318 356
rect 2866 227 2894 356
rect 305 184 734 212
rect 305 181 317 184
rect 259 169 317 181
rect 706 146 734 184
rect 835 215 893 227
rect 835 181 847 215
rect 881 181 893 215
rect 835 169 893 181
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 212 1181 215
rect 2275 215 2333 227
rect 2275 212 2287 215
rect 1169 184 2287 212
rect 1169 181 1181 184
rect 1123 169 1181 181
rect 2275 181 2287 184
rect 2321 181 2333 215
rect 2275 169 2333 181
rect 2851 215 2909 227
rect 2851 181 2863 215
rect 2897 181 2909 215
rect 2851 169 2909 181
rect 2962 146 2990 439
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 355 134 413 146
rect 355 100 367 134
rect 401 100 413 134
rect 355 88 413 100
rect 691 134 749 146
rect 691 100 703 134
rect 737 100 749 134
rect 691 88 749 100
rect 1219 134 1277 146
rect 1219 100 1231 134
rect 1265 100 1277 134
rect 1219 88 1277 100
rect 1555 134 1613 146
rect 1555 100 1567 134
rect 1601 100 1613 134
rect 1555 88 1613 100
rect 1891 134 1949 146
rect 1891 100 1903 134
rect 1937 131 1949 134
rect 2371 134 2429 146
rect 2371 131 2383 134
rect 1937 103 2383 131
rect 1937 100 1949 103
rect 1891 88 1949 100
rect 2371 100 2383 103
rect 2417 100 2429 134
rect 2371 88 2429 100
rect 2707 134 2765 146
rect 2707 100 2719 134
rect 2753 100 2765 134
rect 2707 88 2765 100
rect 2947 134 3005 146
rect 2947 100 2959 134
rect 2993 100 3005 134
rect 2947 88 3005 100
rect 370 48 398 88
rect 1234 48 1262 88
rect 1570 48 1598 88
rect 2722 48 2750 88
rect 0 17 3168 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3168 17
rect 0 -48 3168 -17
<< labels >>
rlabel metal1 0 618 3168 714 0 VPWR
port 3 se
rlabel metal1 0 618 3168 714 0 VPWR
port 3 se
rlabel metal1 0 -48 3168 48 0 VGND
port 2 se
rlabel metal1 0 -48 3168 48 0 VGND
port 2 se
rlabel metal1 115 88 173 146 0 YC
port 4 se
rlabel metal1 130 146 158 439 0 YC
port 4 se
rlabel metal1 115 439 173 497 0 YC
port 4 se
rlabel metal1 2947 88 3005 146 0 YS
port 5 se
rlabel metal1 2962 146 2990 439 0 YS
port 5 se
rlabel metal1 2947 439 3005 497 0 YS
port 5 se
rlabel metal1 835 169 893 227 0 B
port 1 se
rlabel metal1 850 227 878 356 0 B
port 1 se
rlabel metal1 835 356 893 414 0 B
port 1 se
rlabel metal1 1123 169 1181 184 0 A
port 0 se
rlabel metal1 2275 169 2333 184 0 A
port 0 se
rlabel metal1 1123 184 2333 212 0 A
port 0 se
rlabel metal1 1123 212 1181 227 0 A
port 0 se
rlabel metal1 2275 212 2333 227 0 A
port 0 se
rlabel metal1 1138 227 1166 356 0 A
port 0 se
rlabel metal1 2290 227 2318 356 0 A
port 0 se
rlabel metal1 1123 356 1181 414 0 A
port 0 se
rlabel metal1 2275 356 2333 414 0 A
port 0 se
rlabel locali 0 -17 3168 17 4 VGND
port 2 se ground default abutment
rlabel locali 31 17 3137 48 4 VGND
port 2 se ground default abutment
rlabel locali 0 649 3168 683 4 VPWR
port 3 se power default abutment
rlabel metal1 31 618 3137 649 4 VGND
port 2 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 3168 666
<< end >>
