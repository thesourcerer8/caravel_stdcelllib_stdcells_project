magic
tech sky130A
timestamp 1623602988
<< nwell >>
rect 0 179 432 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
<< ndiff >>
rect 82 66 111 69
rect 322 66 351 69
rect 58 63 137 66
rect 58 46 88 63
rect 105 46 137 63
rect 58 24 137 46
rect 152 36 281 66
rect 152 24 184 36
rect 178 19 184 24
rect 201 24 281 36
rect 296 63 375 66
rect 296 46 328 63
rect 345 46 375 63
rect 296 24 375 46
rect 201 19 207 24
rect 178 13 207 19
<< pdiff >>
rect 58 309 87 312
rect 58 306 137 309
rect 58 289 64 306
rect 81 289 137 306
rect 58 225 137 289
rect 152 225 281 309
rect 296 238 375 309
rect 296 225 328 238
rect 322 221 328 225
rect 345 225 375 238
rect 345 221 351 225
rect 322 215 351 221
<< ndiffc >>
rect 88 46 105 63
rect 184 19 201 36
rect 328 46 345 63
<< pdiffc >>
rect 64 289 81 306
rect 328 221 345 238
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 137 206 152 225
rect 281 206 296 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 137 66 152 78
rect 281 66 296 78
rect 137 11 152 24
rect 281 11 296 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 136 86 153 103
rect 280 86 297 103
<< locali >>
rect 56 306 89 314
rect 56 289 64 306
rect 81 289 89 306
rect 56 281 89 289
rect 320 238 353 246
rect 320 221 328 238
rect 345 221 353 238
rect 320 213 353 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 303 206
rect 272 181 280 198
rect 297 196 303 198
rect 297 181 305 196
rect 272 173 305 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 88 305 103
rect 297 86 303 88
rect 272 78 303 86
rect 80 63 111 71
rect 80 46 88 63
rect 105 61 111 63
rect 320 63 353 71
rect 105 46 113 61
rect 80 38 113 46
rect 320 46 328 63
rect 345 46 353 63
rect 176 36 209 44
rect 320 38 353 46
rect 176 11 184 36
rect 201 11 209 36
<< viali >>
rect 64 289 81 306
rect 328 221 345 238
rect 136 181 153 198
rect 280 181 297 198
rect 136 86 153 103
rect 280 86 297 103
rect 88 46 105 63
rect 328 46 345 63
rect 184 19 201 22
rect 184 5 201 19
<< metal1 >>
rect 0 309 432 357
rect 58 306 87 309
rect 58 289 64 306
rect 81 289 87 306
rect 58 283 87 289
rect 322 238 351 244
rect 322 221 328 238
rect 345 221 351 238
rect 322 215 351 221
rect 130 198 159 204
rect 130 181 136 198
rect 153 181 159 198
rect 130 175 159 181
rect 274 198 303 204
rect 274 181 280 198
rect 297 181 303 198
rect 274 175 303 181
rect 137 109 151 175
rect 281 109 295 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 86 159 103
rect 130 80 159 86
rect 274 103 303 109
rect 274 86 280 103
rect 297 86 303 103
rect 274 80 303 86
rect 329 69 343 215
rect 82 63 111 69
rect 82 46 88 63
rect 105 61 111 63
rect 322 63 351 69
rect 322 61 328 63
rect 105 47 328 61
rect 105 46 111 47
rect 82 40 111 46
rect 322 46 328 47
rect 345 46 351 63
rect 322 40 351 46
rect 178 24 207 28
rect 0 22 432 24
rect 0 5 184 22
rect 201 5 432 22
rect 0 -24 432 5
<< labels >>
rlabel metal1 0 309 432 357 0 VDD
port 1 se
rlabel metal1 0 -24 432 24 0 GND
port 2 se
rlabel metal1 82 40 111 47 0 Y
port 3 se
rlabel metal1 322 40 351 47 0 Y
port 4 se
rlabel metal1 82 47 351 61 0 Y
port 5 se
rlabel metal1 82 61 111 69 0 Y
port 6 se
rlabel metal1 322 61 351 69 0 Y
port 7 se
rlabel metal1 329 69 343 215 0 Y
port 8 se
rlabel metal1 322 215 351 244 0 Y
port 9 se
rlabel metal1 130 80 159 109 0 A
port 10 se
rlabel metal1 137 109 151 175 0 A
port 11 se
rlabel metal1 130 175 159 204 0 A
port 12 se
rlabel metal1 274 80 303 109 0 B
port 13 se
rlabel metal1 281 109 295 175 0 B
port 14 se
rlabel metal1 274 175 303 204 0 B
port 15 se
<< properties >>
string FIXED_BBOX 0 0 432 333
<< end >>
