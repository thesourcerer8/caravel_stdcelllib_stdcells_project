VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF2
  CLASS CORE ;
  FOREIGN CLKBUF2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.720 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 18.720 3.570 ;
        RECT 0.580 2.970 0.870 3.090 ;
        RECT 0.580 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.870 2.970 ;
        RECT 0.580 2.740 0.870 2.800 ;
        RECT 3.220 2.970 3.510 3.090 ;
        RECT 3.220 2.800 3.280 2.970 ;
        RECT 3.450 2.800 3.510 2.970 ;
        RECT 3.220 2.740 3.510 2.800 ;
        RECT 6.100 2.970 6.390 3.090 ;
        RECT 6.100 2.800 6.160 2.970 ;
        RECT 6.330 2.800 6.390 2.970 ;
        RECT 6.100 2.740 6.390 2.800 ;
        RECT 8.980 2.970 9.270 3.090 ;
        RECT 8.980 2.800 9.040 2.970 ;
        RECT 9.210 2.800 9.270 2.970 ;
        RECT 8.980 2.740 9.270 2.800 ;
        RECT 11.860 2.970 12.150 3.090 ;
        RECT 11.860 2.800 11.920 2.970 ;
        RECT 12.090 2.800 12.150 2.970 ;
        RECT 11.860 2.740 12.150 2.800 ;
        RECT 14.740 2.970 15.030 3.090 ;
        RECT 14.740 2.800 14.800 2.970 ;
        RECT 14.970 2.800 15.030 2.970 ;
        RECT 14.740 2.740 15.030 2.800 ;
        RECT 17.620 2.970 17.910 3.090 ;
        RECT 17.620 2.800 17.680 2.970 ;
        RECT 17.850 2.800 17.910 2.970 ;
        RECT 17.620 2.740 17.910 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 18.720 3.570 ;
        RECT 0.560 2.970 0.890 3.090 ;
        RECT 0.560 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.890 2.970 ;
        RECT 0.560 2.720 0.890 2.800 ;
        RECT 6.080 2.970 6.410 3.090 ;
        RECT 6.080 2.800 6.160 2.970 ;
        RECT 6.330 2.800 6.410 2.970 ;
        RECT 6.080 2.720 6.410 2.800 ;
        RECT 8.960 2.970 9.290 3.090 ;
        RECT 8.960 2.800 9.040 2.970 ;
        RECT 9.210 2.800 9.290 2.970 ;
        RECT 8.960 2.720 9.290 2.800 ;
        RECT 11.840 2.970 12.170 3.090 ;
        RECT 11.840 2.800 11.920 2.970 ;
        RECT 12.090 2.800 12.170 2.970 ;
        RECT 11.840 2.720 12.170 2.800 ;
        RECT 14.720 2.970 15.050 3.090 ;
        RECT 14.720 2.800 14.800 2.970 ;
        RECT 14.970 2.800 15.050 2.970 ;
        RECT 14.720 2.720 15.050 2.800 ;
        RECT 17.600 2.970 17.930 3.090 ;
        RECT 17.600 2.800 17.680 2.970 ;
        RECT 17.850 2.800 17.930 2.970 ;
        RECT 17.600 2.720 17.930 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.870 0.670 ;
        RECT 0.580 0.440 0.870 0.500 ;
        RECT 3.220 0.670 3.510 0.730 ;
        RECT 3.220 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.510 0.670 ;
        RECT 3.220 0.440 3.510 0.500 ;
        RECT 6.100 0.670 6.390 0.730 ;
        RECT 6.100 0.500 6.160 0.670 ;
        RECT 6.330 0.500 6.390 0.670 ;
        RECT 6.100 0.440 6.390 0.500 ;
        RECT 8.980 0.670 9.270 0.730 ;
        RECT 8.980 0.500 9.040 0.670 ;
        RECT 9.210 0.500 9.270 0.670 ;
        RECT 8.980 0.440 9.270 0.500 ;
        RECT 11.860 0.670 12.150 0.730 ;
        RECT 11.860 0.500 11.920 0.670 ;
        RECT 12.090 0.500 12.150 0.670 ;
        RECT 11.860 0.440 12.150 0.500 ;
        RECT 14.740 0.670 15.030 0.730 ;
        RECT 14.740 0.500 14.800 0.670 ;
        RECT 14.970 0.500 15.030 0.670 ;
        RECT 14.740 0.440 15.030 0.500 ;
        RECT 17.620 0.670 17.910 0.730 ;
        RECT 17.620 0.500 17.680 0.670 ;
        RECT 17.850 0.500 17.910 0.670 ;
        RECT 17.620 0.440 17.910 0.500 ;
        RECT 0.650 0.240 0.790 0.440 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 6.170 0.240 6.310 0.440 ;
        RECT 9.050 0.240 9.190 0.440 ;
        RECT 11.930 0.240 12.070 0.440 ;
        RECT 14.810 0.240 14.950 0.440 ;
        RECT 17.690 0.240 17.830 0.440 ;
        RECT 0.000 -0.240 18.720 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.240 18.720 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 16.180 0.440 16.470 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.370 2.680 2.950 2.820 ;
        RECT 1.370 2.070 1.510 2.680 ;
        RECT 2.810 2.070 2.950 2.680 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 3.200 2.970 3.530 3.050 ;
        RECT 3.200 2.800 3.280 2.970 ;
        RECT 3.450 2.800 3.530 2.970 ;
        RECT 3.200 2.720 3.530 2.800 ;
        RECT 1.760 2.430 2.090 2.510 ;
        RECT 1.760 2.260 1.840 2.430 ;
        RECT 2.010 2.260 2.090 2.430 ;
        RECT 1.780 2.180 2.090 2.260 ;
        RECT 4.640 2.430 4.970 2.510 ;
        RECT 4.640 2.260 4.720 2.430 ;
        RECT 4.890 2.260 4.970 2.430 ;
        RECT 4.640 2.180 4.970 2.260 ;
        RECT 5.680 2.090 5.850 2.660 ;
        RECT 7.520 2.430 7.850 2.510 ;
        RECT 7.520 2.260 7.600 2.430 ;
        RECT 7.770 2.260 7.850 2.430 ;
        RECT 7.540 2.180 7.850 2.260 ;
        RECT 8.560 2.090 8.730 2.660 ;
        RECT 10.400 2.430 10.730 2.510 ;
        RECT 10.400 2.260 10.480 2.430 ;
        RECT 10.650 2.260 10.730 2.430 ;
        RECT 10.420 2.180 10.730 2.260 ;
        RECT 11.440 2.090 11.610 2.660 ;
        RECT 13.280 2.430 13.610 2.510 ;
        RECT 13.280 2.260 13.360 2.430 ;
        RECT 13.530 2.260 13.610 2.430 ;
        RECT 13.300 2.180 13.610 2.260 ;
        RECT 14.320 2.090 14.490 2.660 ;
        RECT 16.160 2.430 16.490 2.510 ;
        RECT 16.160 2.260 16.240 2.430 ;
        RECT 16.410 2.260 16.490 2.430 ;
        RECT 16.160 2.180 16.490 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.470 2.090 ;
        RECT 5.600 2.010 5.930 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 7.040 2.010 7.370 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 8.480 2.010 8.810 2.090 ;
        RECT 8.480 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.810 2.010 ;
        RECT 8.480 1.760 8.810 1.840 ;
        RECT 9.920 2.010 10.250 2.090 ;
        RECT 9.920 1.840 10.000 2.010 ;
        RECT 10.170 1.840 10.250 2.010 ;
        RECT 9.920 1.760 10.250 1.840 ;
        RECT 11.360 2.010 11.690 2.090 ;
        RECT 11.360 1.840 11.440 2.010 ;
        RECT 11.610 1.840 11.690 2.010 ;
        RECT 11.360 1.760 11.690 1.840 ;
        RECT 12.800 2.010 13.130 2.090 ;
        RECT 12.800 1.840 12.880 2.010 ;
        RECT 13.050 1.840 13.130 2.010 ;
        RECT 12.800 1.760 13.130 1.840 ;
        RECT 14.240 2.010 14.570 2.090 ;
        RECT 14.240 1.840 14.320 2.010 ;
        RECT 14.490 1.840 14.570 2.010 ;
        RECT 14.240 1.760 14.570 1.840 ;
        RECT 15.680 2.010 15.990 2.090 ;
        RECT 15.680 1.840 15.760 2.010 ;
        RECT 15.930 1.840 16.010 2.010 ;
        RECT 15.680 1.760 16.010 1.840 ;
        RECT 2.800 1.160 2.970 1.760 ;
        RECT 5.680 1.620 5.850 1.760 ;
        RECT 8.560 1.620 8.730 1.760 ;
        RECT 11.440 1.620 11.610 1.760 ;
        RECT 14.320 1.620 14.490 1.760 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.920 1.610 1.080 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 1.530 0.910 1.590 0.920 ;
        RECT 1.280 0.830 1.590 0.910 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.920 4.490 1.080 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 4.410 0.910 4.470 0.920 ;
        RECT 4.160 0.830 4.470 0.910 ;
        RECT 5.600 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.600 0.830 5.930 0.910 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.920 7.370 1.080 ;
        RECT 8.480 1.080 8.810 1.160 ;
        RECT 7.290 0.910 7.350 0.920 ;
        RECT 7.040 0.830 7.350 0.910 ;
        RECT 8.480 0.910 8.560 1.080 ;
        RECT 8.730 0.920 8.810 1.080 ;
        RECT 9.920 1.080 10.250 1.160 ;
        RECT 8.730 0.910 8.790 0.920 ;
        RECT 8.480 0.830 8.790 0.910 ;
        RECT 9.920 0.910 10.000 1.080 ;
        RECT 10.170 0.920 10.250 1.080 ;
        RECT 11.360 1.080 11.690 1.160 ;
        RECT 10.170 0.910 10.230 0.920 ;
        RECT 9.920 0.830 10.230 0.910 ;
        RECT 11.360 0.910 11.440 1.080 ;
        RECT 11.610 0.910 11.690 1.080 ;
        RECT 11.360 0.830 11.690 0.910 ;
        RECT 12.800 1.080 13.130 1.160 ;
        RECT 12.800 0.910 12.880 1.080 ;
        RECT 13.050 0.920 13.130 1.080 ;
        RECT 14.240 1.080 14.570 1.160 ;
        RECT 13.050 0.910 13.110 0.920 ;
        RECT 12.800 0.830 13.110 0.910 ;
        RECT 14.240 0.910 14.320 1.080 ;
        RECT 14.490 0.920 14.570 1.080 ;
        RECT 15.680 1.080 16.010 1.160 ;
        RECT 14.490 0.910 14.550 0.920 ;
        RECT 14.240 0.830 14.550 0.910 ;
        RECT 15.680 0.910 15.760 1.080 ;
        RECT 15.930 0.920 16.010 1.080 ;
        RECT 15.930 0.910 15.990 0.920 ;
        RECT 15.680 0.830 15.990 0.910 ;
        RECT 16.240 0.750 16.410 2.180 ;
        RECT 17.120 2.010 17.450 2.090 ;
        RECT 17.120 1.840 17.200 2.010 ;
        RECT 17.370 1.840 17.450 2.010 ;
        RECT 17.120 1.760 17.450 1.840 ;
        RECT 17.120 1.080 17.450 1.160 ;
        RECT 17.120 0.910 17.200 1.080 ;
        RECT 17.370 0.910 17.450 1.080 ;
        RECT 17.120 0.830 17.450 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 1.760 0.670 2.090 0.750 ;
        RECT 1.760 0.500 1.840 0.670 ;
        RECT 2.010 0.500 2.090 0.670 ;
        RECT 3.220 0.670 3.530 0.750 ;
        RECT 3.220 0.660 3.280 0.670 ;
        RECT 1.760 0.420 2.090 0.500 ;
        RECT 3.200 0.500 3.280 0.660 ;
        RECT 3.450 0.500 3.530 0.670 ;
        RECT 3.200 0.420 3.530 0.500 ;
        RECT 4.640 0.670 4.970 0.750 ;
        RECT 4.640 0.500 4.720 0.670 ;
        RECT 4.890 0.500 4.970 0.670 ;
        RECT 6.100 0.670 6.410 0.750 ;
        RECT 6.100 0.660 6.160 0.670 ;
        RECT 4.640 0.420 4.970 0.500 ;
        RECT 6.080 0.500 6.160 0.660 ;
        RECT 6.330 0.500 6.410 0.670 ;
        RECT 6.080 0.420 6.410 0.500 ;
        RECT 7.520 0.670 7.850 0.750 ;
        RECT 7.520 0.500 7.600 0.670 ;
        RECT 7.770 0.500 7.850 0.670 ;
        RECT 7.520 0.420 7.850 0.500 ;
        RECT 8.960 0.670 9.290 0.750 ;
        RECT 8.960 0.500 9.040 0.670 ;
        RECT 9.210 0.500 9.290 0.670 ;
        RECT 8.960 0.420 9.290 0.500 ;
        RECT 10.400 0.670 10.730 0.750 ;
        RECT 10.400 0.500 10.480 0.670 ;
        RECT 10.650 0.500 10.730 0.670 ;
        RECT 11.860 0.670 12.170 0.750 ;
        RECT 11.860 0.660 11.920 0.670 ;
        RECT 10.400 0.420 10.730 0.500 ;
        RECT 11.840 0.500 11.920 0.660 ;
        RECT 12.090 0.500 12.170 0.670 ;
        RECT 11.840 0.420 12.170 0.500 ;
        RECT 13.280 0.670 13.610 0.750 ;
        RECT 13.280 0.500 13.360 0.670 ;
        RECT 13.530 0.500 13.610 0.670 ;
        RECT 13.280 0.420 13.610 0.500 ;
        RECT 14.720 0.670 15.050 0.750 ;
        RECT 14.720 0.500 14.800 0.670 ;
        RECT 14.970 0.500 15.050 0.670 ;
        RECT 14.720 0.420 15.050 0.500 ;
        RECT 16.160 0.670 16.490 0.750 ;
        RECT 16.160 0.500 16.240 0.670 ;
        RECT 16.410 0.500 16.490 0.670 ;
        RECT 17.620 0.670 17.930 0.750 ;
        RECT 17.620 0.660 17.680 0.670 ;
        RECT 16.160 0.420 16.490 0.500 ;
        RECT 17.600 0.500 17.680 0.660 ;
        RECT 17.850 0.500 17.930 0.670 ;
        RECT 17.600 0.420 17.930 0.500 ;
      LAYER met1 ;
        RECT 5.620 2.830 5.910 2.890 ;
        RECT 5.620 2.820 5.680 2.830 ;
        RECT 4.250 2.680 5.680 2.820 ;
        RECT 1.780 2.430 2.070 2.490 ;
        RECT 1.780 2.260 1.840 2.430 ;
        RECT 2.010 2.260 2.070 2.430 ;
        RECT 1.780 2.200 2.070 2.260 ;
        RECT 1.850 1.060 1.990 2.200 ;
        RECT 4.250 2.070 4.390 2.680 ;
        RECT 5.620 2.660 5.680 2.680 ;
        RECT 5.850 2.660 5.910 2.830 ;
        RECT 8.500 2.830 8.790 2.890 ;
        RECT 8.500 2.820 8.560 2.830 ;
        RECT 5.620 2.600 5.910 2.660 ;
        RECT 7.130 2.680 8.560 2.820 ;
        RECT 4.660 2.430 4.950 2.490 ;
        RECT 4.660 2.260 4.720 2.430 ;
        RECT 4.890 2.260 4.950 2.430 ;
        RECT 4.660 2.200 4.950 2.260 ;
        RECT 4.180 2.010 4.470 2.070 ;
        RECT 4.180 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.470 2.010 ;
        RECT 4.180 1.780 4.470 1.840 ;
        RECT 4.730 2.000 4.870 2.200 ;
        RECT 7.130 2.070 7.270 2.680 ;
        RECT 8.500 2.660 8.560 2.680 ;
        RECT 8.730 2.660 8.790 2.830 ;
        RECT 11.380 2.830 11.670 2.890 ;
        RECT 11.380 2.820 11.440 2.830 ;
        RECT 8.500 2.600 8.790 2.660 ;
        RECT 10.010 2.680 11.440 2.820 ;
        RECT 7.540 2.430 7.830 2.490 ;
        RECT 7.540 2.260 7.600 2.430 ;
        RECT 7.770 2.260 7.830 2.430 ;
        RECT 7.540 2.200 7.830 2.260 ;
        RECT 7.060 2.010 7.350 2.070 ;
        RECT 7.060 2.000 7.120 2.010 ;
        RECT 4.730 1.860 7.120 2.000 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 4.180 1.080 4.470 1.140 ;
        RECT 4.180 1.060 4.240 1.080 ;
        RECT 1.850 0.920 4.240 1.060 ;
        RECT 1.850 0.730 1.990 0.920 ;
        RECT 4.180 0.910 4.240 0.920 ;
        RECT 4.410 0.910 4.470 1.080 ;
        RECT 4.180 0.850 4.470 0.910 ;
        RECT 4.730 0.730 4.870 1.860 ;
        RECT 7.060 1.840 7.120 1.860 ;
        RECT 7.290 1.840 7.350 2.010 ;
        RECT 7.060 1.780 7.350 1.840 ;
        RECT 7.610 2.000 7.750 2.200 ;
        RECT 10.010 2.070 10.150 2.680 ;
        RECT 11.380 2.660 11.440 2.680 ;
        RECT 11.610 2.660 11.670 2.830 ;
        RECT 14.260 2.830 14.550 2.890 ;
        RECT 14.260 2.820 14.320 2.830 ;
        RECT 11.380 2.600 11.670 2.660 ;
        RECT 12.890 2.680 14.320 2.820 ;
        RECT 10.420 2.430 10.710 2.490 ;
        RECT 10.420 2.260 10.480 2.430 ;
        RECT 10.650 2.260 10.710 2.430 ;
        RECT 10.420 2.200 10.710 2.260 ;
        RECT 9.940 2.010 10.230 2.070 ;
        RECT 9.940 2.000 10.000 2.010 ;
        RECT 7.610 1.860 10.000 2.000 ;
        RECT 5.620 1.620 5.910 1.680 ;
        RECT 5.620 1.450 5.680 1.620 ;
        RECT 5.850 1.450 5.910 1.620 ;
        RECT 5.620 1.390 5.910 1.450 ;
        RECT 5.690 1.140 5.830 1.390 ;
        RECT 7.130 1.140 7.270 1.780 ;
        RECT 5.620 1.080 5.910 1.140 ;
        RECT 5.620 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.910 1.080 ;
        RECT 5.620 0.850 5.910 0.910 ;
        RECT 7.060 1.080 7.350 1.140 ;
        RECT 7.060 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.350 1.080 ;
        RECT 7.060 0.850 7.350 0.910 ;
        RECT 7.610 0.730 7.750 1.860 ;
        RECT 9.940 1.840 10.000 1.860 ;
        RECT 10.170 1.840 10.230 2.010 ;
        RECT 9.940 1.780 10.230 1.840 ;
        RECT 10.490 2.000 10.630 2.200 ;
        RECT 12.890 2.070 13.030 2.680 ;
        RECT 14.260 2.660 14.320 2.680 ;
        RECT 14.490 2.660 14.550 2.830 ;
        RECT 14.260 2.600 14.550 2.660 ;
        RECT 13.300 2.430 13.590 2.490 ;
        RECT 13.300 2.260 13.360 2.430 ;
        RECT 13.530 2.260 13.590 2.430 ;
        RECT 13.300 2.200 13.590 2.260 ;
        RECT 12.820 2.010 13.110 2.070 ;
        RECT 12.820 2.000 12.880 2.010 ;
        RECT 10.490 1.860 12.880 2.000 ;
        RECT 8.500 1.620 8.790 1.680 ;
        RECT 8.500 1.450 8.560 1.620 ;
        RECT 8.730 1.450 8.790 1.620 ;
        RECT 8.500 1.390 8.790 1.450 ;
        RECT 8.570 1.140 8.710 1.390 ;
        RECT 10.010 1.140 10.150 1.780 ;
        RECT 8.500 1.080 8.790 1.140 ;
        RECT 8.500 0.910 8.560 1.080 ;
        RECT 8.730 0.910 8.790 1.080 ;
        RECT 8.500 0.850 8.790 0.910 ;
        RECT 9.940 1.080 10.230 1.140 ;
        RECT 9.940 0.910 10.000 1.080 ;
        RECT 10.170 0.910 10.230 1.080 ;
        RECT 9.940 0.850 10.230 0.910 ;
        RECT 10.490 0.730 10.630 1.860 ;
        RECT 12.820 1.840 12.880 1.860 ;
        RECT 13.050 1.840 13.110 2.010 ;
        RECT 12.820 1.780 13.110 1.840 ;
        RECT 13.370 2.000 13.510 2.200 ;
        RECT 15.700 2.010 15.990 2.070 ;
        RECT 15.700 2.000 15.760 2.010 ;
        RECT 13.370 1.860 15.760 2.000 ;
        RECT 11.380 1.620 11.670 1.680 ;
        RECT 11.380 1.450 11.440 1.620 ;
        RECT 11.610 1.450 11.670 1.620 ;
        RECT 11.380 1.390 11.670 1.450 ;
        RECT 11.450 1.140 11.590 1.390 ;
        RECT 12.890 1.140 13.030 1.780 ;
        RECT 11.380 1.080 11.670 1.140 ;
        RECT 11.380 0.910 11.440 1.080 ;
        RECT 11.610 0.910 11.670 1.080 ;
        RECT 11.380 0.850 11.670 0.910 ;
        RECT 12.820 1.080 13.110 1.140 ;
        RECT 12.820 0.910 12.880 1.080 ;
        RECT 13.050 0.910 13.110 1.080 ;
        RECT 12.820 0.850 13.110 0.910 ;
        RECT 13.370 0.730 13.510 1.860 ;
        RECT 15.700 1.840 15.760 1.860 ;
        RECT 15.930 2.000 15.990 2.010 ;
        RECT 17.140 2.010 17.430 2.070 ;
        RECT 17.140 2.000 17.200 2.010 ;
        RECT 15.930 1.860 17.200 2.000 ;
        RECT 15.930 1.840 15.990 1.860 ;
        RECT 15.700 1.780 15.990 1.840 ;
        RECT 17.140 1.840 17.200 1.860 ;
        RECT 17.370 1.840 17.430 2.010 ;
        RECT 17.140 1.780 17.430 1.840 ;
        RECT 14.260 1.620 14.550 1.680 ;
        RECT 14.260 1.450 14.320 1.620 ;
        RECT 14.490 1.450 14.550 1.620 ;
        RECT 14.260 1.390 14.550 1.450 ;
        RECT 14.330 1.140 14.470 1.390 ;
        RECT 15.770 1.140 15.910 1.780 ;
        RECT 17.210 1.140 17.350 1.780 ;
        RECT 14.260 1.080 14.550 1.140 ;
        RECT 14.260 0.910 14.320 1.080 ;
        RECT 14.490 0.910 14.550 1.080 ;
        RECT 14.260 0.850 14.550 0.910 ;
        RECT 15.700 1.080 15.990 1.140 ;
        RECT 15.700 0.910 15.760 1.080 ;
        RECT 15.930 0.910 15.990 1.080 ;
        RECT 15.700 0.850 15.990 0.910 ;
        RECT 17.140 1.080 17.430 1.140 ;
        RECT 17.140 0.910 17.200 1.080 ;
        RECT 17.370 0.910 17.430 1.080 ;
        RECT 17.140 0.850 17.430 0.910 ;
        RECT 1.780 0.670 2.070 0.730 ;
        RECT 1.780 0.500 1.840 0.670 ;
        RECT 2.010 0.500 2.070 0.670 ;
        RECT 1.780 0.440 2.070 0.500 ;
        RECT 4.660 0.670 4.950 0.730 ;
        RECT 4.660 0.500 4.720 0.670 ;
        RECT 4.890 0.500 4.950 0.670 ;
        RECT 4.660 0.440 4.950 0.500 ;
        RECT 7.540 0.670 7.830 0.730 ;
        RECT 7.540 0.500 7.600 0.670 ;
        RECT 7.770 0.500 7.830 0.670 ;
        RECT 7.540 0.440 7.830 0.500 ;
        RECT 10.420 0.670 10.710 0.730 ;
        RECT 10.420 0.500 10.480 0.670 ;
        RECT 10.650 0.500 10.710 0.670 ;
        RECT 10.420 0.440 10.710 0.500 ;
        RECT 13.300 0.670 13.590 0.730 ;
        RECT 13.300 0.500 13.360 0.670 ;
        RECT 13.530 0.500 13.590 0.670 ;
        RECT 13.300 0.440 13.590 0.500 ;
  END
END CLKBUF2
END LIBRARY

