magic
tech sky130A
magscale 1 2
timestamp 1636962382
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1728 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 355 134 413 146
rect 355 132 367 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 931 134 989 146
rect 931 132 943 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 48 849 132
rect 879 100 943 132
rect 977 132 989 134
rect 1507 134 1565 146
rect 1507 132 1519 134
rect 977 100 1137 132
rect 879 48 1137 100
rect 1167 48 1425 132
rect 1455 100 1519 132
rect 1553 132 1565 134
rect 1553 100 1613 132
rect 1455 48 1613 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 593 561 618
rect 303 559 367 593
rect 401 559 561 593
rect 303 450 561 559
rect 591 450 849 618
rect 879 485 1137 618
rect 879 451 943 485
rect 977 451 1137 485
rect 879 450 1137 451
rect 1167 450 1425 618
rect 1455 593 1613 618
rect 1455 559 1519 593
rect 1553 559 1613 593
rect 1455 450 1613 559
rect 115 439 173 450
rect 931 439 989 450
<< ndiffc >>
rect 127 100 161 134
rect 367 100 401 134
rect 943 100 977 134
rect 1519 100 1553 134
<< pdiffc >>
rect 127 451 161 485
rect 367 559 401 593
rect 943 451 977 485
rect 1519 559 1553 593
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1728 683
rect 31 643 1697 649
rect 31 618 1469 643
rect 1603 618 1697 643
rect 351 593 417 618
rect 351 559 367 593
rect 401 559 417 593
rect 351 543 417 559
rect 1503 593 1569 609
rect 1503 559 1519 593
rect 1553 559 1569 593
rect 1503 543 1569 559
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 927 485 993 501
rect 927 451 943 485
rect 977 451 993 485
rect 927 436 993 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 893 418
rect 1119 402 1185 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 271 231 305 352
rect 559 296 593 352
rect 559 231 593 262
rect 255 215 321 231
rect 255 181 271 215
rect 305 184 321 215
rect 543 215 609 231
rect 305 181 317 184
rect 255 165 317 181
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 184 897 215
rect 881 181 893 184
rect 831 165 893 181
rect 943 150 977 368
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 184 1473 215
rect 1457 181 1469 184
rect 1407 165 1469 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 351 134 417 150
rect 351 100 367 134
rect 401 100 417 134
rect 351 84 417 100
rect 927 134 993 150
rect 927 100 943 134
rect 977 100 993 134
rect 927 84 993 100
rect 1503 134 1569 150
rect 1503 100 1519 134
rect 1553 100 1569 134
rect 1503 84 1569 100
rect 31 17 1697 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1728 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 367 559 401 593
rect 1519 559 1553 593
rect 127 451 161 485
rect 943 451 977 485
rect 847 368 881 402
rect 943 368 977 402
rect 559 262 593 296
rect 271 181 305 215
rect 847 181 881 215
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 127 100 161 134
rect 367 100 401 134
rect 1519 100 1553 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1728 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1728 683
rect 0 618 1728 649
rect 355 593 413 618
rect 355 559 367 593
rect 401 559 413 593
rect 355 547 413 559
rect 1507 593 1565 618
rect 1507 559 1519 593
rect 1553 559 1565 593
rect 1507 547 1565 559
rect 115 485 173 497
rect 115 451 127 485
rect 161 451 173 485
rect 115 439 173 451
rect 931 485 989 497
rect 931 451 943 485
rect 977 451 989 485
rect 130 399 158 439
rect 835 402 893 414
rect 835 399 847 402
rect 130 371 847 399
rect 130 146 158 371
rect 835 368 847 371
rect 881 368 893 402
rect 835 356 893 368
rect 931 402 989 451
rect 931 368 943 402
rect 977 368 989 402
rect 931 356 989 368
rect 1123 402 1181 414
rect 1123 368 1135 402
rect 1169 399 1181 402
rect 1411 402 1469 414
rect 1169 371 1262 399
rect 1169 368 1181 371
rect 1123 356 1181 368
rect 850 320 878 356
rect 547 296 605 308
rect 547 262 559 296
rect 593 262 605 296
rect 850 292 1166 320
rect 547 250 605 262
rect 1138 227 1166 292
rect 259 215 317 227
rect 259 181 271 215
rect 305 212 317 215
rect 835 215 893 227
rect 835 212 847 215
rect 305 184 847 212
rect 305 181 317 184
rect 259 169 317 181
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 355 134 413 146
rect 355 100 367 134
rect 401 100 413 134
rect 850 131 878 169
rect 1234 131 1262 371
rect 1411 368 1423 402
rect 1457 368 1469 402
rect 1411 356 1469 368
rect 1426 227 1454 356
rect 1411 215 1469 227
rect 1411 181 1423 215
rect 1457 181 1469 215
rect 1411 169 1469 181
rect 850 103 1262 131
rect 1507 134 1565 146
rect 355 88 413 100
rect 1507 100 1519 134
rect 1553 100 1565 134
rect 1507 88 1565 100
rect 370 48 398 88
rect 1522 48 1550 88
rect 0 17 1728 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1728 17
rect 0 -48 1728 -17
<< labels >>
rlabel metal1 0 618 1728 714 0 VPWR
port 4 se
rlabel metal1 0 618 1728 714 0 VPWR
port 4 se
rlabel metal1 0 -48 1728 48 0 VGND
port 3 se
rlabel metal1 0 -48 1728 48 0 VGND
port 3 se
rlabel metal1 931 356 989 497 0 Y
port 5 se
rlabel metal1 1411 169 1469 227 0 B
port 1 se
rlabel metal1 1426 227 1454 356 0 B
port 1 se
rlabel metal1 1411 356 1469 414 0 B
port 1 se
rlabel metal1 850 103 1262 131 0 S
port 2 se
rlabel metal1 850 131 878 169 0 S
port 2 se
rlabel metal1 259 169 317 184 0 S
port 2 se
rlabel metal1 835 169 893 184 0 S
port 2 se
rlabel metal1 259 184 893 212 0 S
port 2 se
rlabel metal1 259 212 317 227 0 S
port 2 se
rlabel metal1 835 212 893 227 0 S
port 2 se
rlabel metal1 1123 356 1181 371 0 S
port 2 se
rlabel metal1 1234 131 1262 371 0 S
port 2 se
rlabel metal1 1123 371 1262 399 0 S
port 2 se
rlabel metal1 1123 399 1181 414 0 S
port 2 se
rlabel metal1 547 250 605 308 0 A
port 0 se
rlabel locali 0 -17 1728 17 4 VGND
port 3 se ground default abutment
rlabel locali 31 17 1697 48 4 VGND
port 3 se ground default abutment
rlabel locali 0 649 1728 683 4 VPWR
port 4 se power default abutment
rlabel metal1 31 618 1697 649 4 VGND
port 3 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1728 666
<< end >>
