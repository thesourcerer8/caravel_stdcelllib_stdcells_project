VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.370 0.870 2.440 ;
        RECT 3.220 2.370 3.510 2.440 ;
        RECT 0.580 2.230 3.510 2.370 ;
        RECT 0.580 2.150 0.870 2.230 ;
        RECT 3.220 2.150 3.510 2.230 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 3.290 0.690 3.430 2.150 ;
        RECT 0.580 0.400 0.870 0.690 ;
        RECT 3.220 0.400 3.510 0.690 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.960 1.590 2.040 ;
        RECT 2.740 1.960 3.030 2.040 ;
        RECT 1.300 1.820 3.030 1.960 ;
        RECT 1.300 1.750 1.590 1.820 ;
        RECT 2.740 1.750 3.030 1.820 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
        RECT 2.740 0.800 3.030 1.090 ;
    END
  END A
END INVX4
END LIBRARY

