magic
tech sky130A
magscale 1 2
timestamp 1624196784
<< locali >>
rect 34111 38090 34145 38204
rect 32575 32096 32609 32210
rect 8095 22442 8383 22476
rect 8095 22180 8129 22442
rect 27199 22254 27233 22442
rect 34399 20774 34433 20888
rect 8191 19812 8225 19852
rect 8191 19778 8383 19812
rect 8417 18520 8513 18554
rect 8479 18480 8513 18520
rect 8479 18446 8575 18480
rect 7903 17148 7937 17188
rect 8191 17148 8225 17188
rect 7903 17114 8225 17148
rect 56959 10340 56993 10454
rect 7711 9196 7937 9230
rect 7711 9156 7745 9196
rect 7903 9156 7937 9196
rect 8191 9196 8513 9230
rect 8191 9156 8225 9196
rect 7903 9122 8225 9156
rect 8479 9156 8513 9196
rect 42751 8786 42785 8900
rect 14527 8120 14561 8530
rect 8479 7864 8801 7898
rect 8479 7824 8513 7864
rect 8383 7790 8513 7824
rect 8767 7824 8801 7864
rect 8383 7676 8417 7790
rect 39487 6936 39521 7124
rect 7903 6532 8225 6566
rect 7903 6492 7937 6532
rect 7745 6458 7937 6492
rect 8191 6492 8225 6532
rect 8479 6492 8513 6532
rect 8191 6458 8513 6492
rect 11551 5456 11585 5718
rect 21631 5530 21665 5644
rect 26623 5530 26657 5644
rect 7711 5160 7745 5200
rect 7903 5200 8225 5234
rect 7903 5160 7937 5200
rect 7711 5126 7937 5160
rect 8191 5160 8225 5200
rect 8479 5160 8513 5200
rect 8191 5126 8513 5160
rect 53119 2866 53153 3054
<< viali >>
rect 9919 57000 9953 57034
rect 13951 57000 13985 57034
rect 21535 57000 21569 57034
rect 32671 57000 32705 57034
rect 1951 56926 1985 56960
rect 2815 56926 2849 56960
rect 5311 56926 5345 56960
rect 5791 56926 5825 56960
rect 7423 56926 7457 56960
rect 8095 56926 8129 56960
rect 11455 56926 11489 56960
rect 13183 56926 13217 56960
rect 15103 56926 15137 56960
rect 16351 56926 16385 56960
rect 17791 56926 17825 56960
rect 19519 56926 19553 56960
rect 20671 56926 20705 56960
rect 23551 56926 23585 56960
rect 24031 56926 24065 56960
rect 26239 56926 26273 56960
rect 27007 56926 27041 56960
rect 29023 56926 29057 56960
rect 30079 56926 30113 56960
rect 32095 56926 32129 56960
rect 34303 56926 34337 56960
rect 35263 56926 35297 56960
rect 36607 56926 36641 56960
rect 41983 56926 42017 56960
rect 47551 56926 47585 56960
rect 52735 56926 52769 56960
rect 1759 56852 1793 56886
rect 2623 56852 2657 56886
rect 5119 56852 5153 56886
rect 7231 56852 7265 56886
rect 11263 56852 11297 56886
rect 12991 56852 13025 56886
rect 13759 56852 13793 56886
rect 14047 56852 14081 56886
rect 16159 56852 16193 56886
rect 19327 56852 19361 56886
rect 21343 56852 21377 56886
rect 21631 56852 21665 56886
rect 23359 56852 23393 56886
rect 26047 56852 26081 56886
rect 28831 56852 28865 56886
rect 31903 56852 31937 56886
rect 32767 56852 32801 56886
rect 34111 56852 34145 56886
rect 35071 56852 35105 56886
rect 38239 56852 38273 56886
rect 40063 56852 40097 56886
rect 40735 56852 40769 56886
rect 41023 56852 41057 56886
rect 43231 56852 43265 56886
rect 45055 56852 45089 56886
rect 46303 56852 46337 56886
rect 48991 56852 49025 56886
rect 51103 56852 51137 56886
rect 54271 56852 54305 56886
rect 55807 56852 55841 56886
rect 57055 56852 57089 56886
rect 9823 56704 9857 56738
rect 37951 56704 37985 56738
rect 39775 56704 39809 56738
rect 40447 56704 40481 56738
rect 40831 56704 40865 56738
rect 42943 56704 42977 56738
rect 44767 56704 44801 56738
rect 46015 56704 46049 56738
rect 48703 56704 48737 56738
rect 50815 56704 50849 56738
rect 53983 56704 54017 56738
rect 55519 56704 55553 56738
rect 56767 56704 56801 56738
rect 1663 56482 1697 56516
rect 2431 56482 2465 56516
rect 3199 56482 3233 56516
rect 4447 56482 4481 56516
rect 5503 56482 5537 56516
rect 6271 56482 6305 56516
rect 7135 56482 7169 56516
rect 8479 56482 8513 56516
rect 10303 56482 10337 56516
rect 11071 56482 11105 56516
rect 11839 56482 11873 56516
rect 12607 56482 12641 56516
rect 13471 56482 13505 56516
rect 15007 56482 15041 56516
rect 17119 56482 17153 56516
rect 18751 56482 18785 56516
rect 20287 56482 20321 56516
rect 21343 56482 21377 56516
rect 22207 56482 22241 56516
rect 22879 56482 22913 56516
rect 24319 56482 24353 56516
rect 26047 56482 26081 56516
rect 26815 56482 26849 56516
rect 27679 56482 27713 56516
rect 28543 56482 28577 56516
rect 29695 56482 29729 56516
rect 30847 56482 30881 56516
rect 32383 56482 32417 56516
rect 33151 56482 33185 56516
rect 33919 56482 33953 56516
rect 34687 56482 34721 56516
rect 36127 56482 36161 56516
rect 36991 56482 37025 56516
rect 37759 56482 37793 56516
rect 38815 56482 38849 56516
rect 40255 56482 40289 56516
rect 41887 56482 41921 56516
rect 42751 56482 42785 56516
rect 43423 56482 43457 56516
rect 44287 56482 44321 56516
rect 45055 56482 45089 56516
rect 46783 56482 46817 56516
rect 48127 56482 48161 56516
rect 48991 56482 49025 56516
rect 49759 56482 49793 56516
rect 50623 56482 50657 56516
rect 53023 56482 53057 56516
rect 53791 56482 53825 56516
rect 54463 56482 54497 56516
rect 55327 56482 55361 56516
rect 55999 56482 56033 56516
rect 33247 56334 33281 56368
rect 56095 56334 56129 56368
rect 7231 56260 7265 56294
rect 15487 56260 15521 56294
rect 15775 56260 15809 56294
rect 45151 56260 45185 56294
rect 49855 56260 49889 56294
rect 52255 56260 52289 56294
rect 57151 56260 57185 56294
rect 1759 56186 1793 56220
rect 2239 56186 2273 56220
rect 2527 56186 2561 56220
rect 3007 56186 3041 56220
rect 3295 56186 3329 56220
rect 4543 56186 4577 56220
rect 5215 56186 5249 56220
rect 5599 56186 5633 56220
rect 6079 56186 6113 56220
rect 6367 56186 6401 56220
rect 8287 56186 8321 56220
rect 8575 56186 8609 56220
rect 10399 56186 10433 56220
rect 10783 56186 10817 56220
rect 11167 56186 11201 56220
rect 11935 56186 11969 56220
rect 12703 56186 12737 56220
rect 13279 56186 13313 56220
rect 13567 56186 13601 56220
rect 15103 56186 15137 56220
rect 15871 56186 15905 56220
rect 16831 56186 16865 56220
rect 17215 56186 17249 56220
rect 18463 56186 18497 56220
rect 18655 56186 18689 56220
rect 20095 56186 20129 56220
rect 20383 56186 20417 56220
rect 21151 56186 21185 56220
rect 21439 56186 21473 56220
rect 21919 56186 21953 56220
rect 22111 56186 22145 56220
rect 22975 56186 23009 56220
rect 24415 56186 24449 56220
rect 26143 56186 26177 56220
rect 26911 56186 26945 56220
rect 27487 56186 27521 56220
rect 27775 56186 27809 56220
rect 28159 56186 28193 56220
rect 28447 56186 28481 56220
rect 29407 56186 29441 56220
rect 29599 56186 29633 56220
rect 30943 56186 30977 56220
rect 31327 56186 31361 56220
rect 31615 56186 31649 56220
rect 31711 56186 31745 56220
rect 32479 56186 32513 56220
rect 34015 56186 34049 56220
rect 34495 56186 34529 56220
rect 34783 56186 34817 56220
rect 36223 56186 36257 56220
rect 36703 56186 36737 56220
rect 36895 56186 36929 56220
rect 37471 56186 37505 56220
rect 37663 56186 37697 56220
rect 37951 56186 37985 56220
rect 38431 56186 38465 56220
rect 38719 56186 38753 56220
rect 39871 56186 39905 56220
rect 40159 56186 40193 56220
rect 41695 56186 41729 56220
rect 41983 56186 42017 56220
rect 42463 56186 42497 56220
rect 42655 56186 42689 56220
rect 43519 56186 43553 56220
rect 43999 56186 44033 56220
rect 44191 56186 44225 56220
rect 44479 56186 44513 56220
rect 46495 56186 46529 56220
rect 46687 56186 46721 56220
rect 48223 56186 48257 56220
rect 48607 56186 48641 56220
rect 48895 56186 48929 56220
rect 50239 56186 50273 56220
rect 50527 56186 50561 56220
rect 51679 56186 51713 56220
rect 51967 56186 52001 56220
rect 52063 56186 52097 56220
rect 52735 56186 52769 56220
rect 52927 56186 52961 56220
rect 53503 56186 53537 56220
rect 53695 56186 53729 56220
rect 53983 56186 54017 56220
rect 54559 56186 54593 56220
rect 54943 56186 54977 56220
rect 55231 56186 55265 56220
rect 1663 55668 1697 55702
rect 4447 55668 4481 55702
rect 7615 55668 7649 55702
rect 9343 55668 9377 55702
rect 13951 55668 13985 55702
rect 20383 55668 20417 55702
rect 23455 55668 23489 55702
rect 25087 55668 25121 55702
rect 39295 55668 39329 55702
rect 40831 55668 40865 55702
rect 45631 55668 45665 55702
rect 46303 55668 46337 55702
rect 47167 55668 47201 55702
rect 51871 55668 51905 55702
rect 56671 55668 56705 55702
rect 57727 55668 57761 55702
rect 46783 55594 46817 55628
rect 47071 55594 47105 55628
rect 1759 55520 1793 55554
rect 4255 55520 4289 55554
rect 4543 55520 4577 55554
rect 7711 55520 7745 55554
rect 9247 55520 9281 55554
rect 14047 55520 14081 55554
rect 17791 55520 17825 55554
rect 20287 55520 20321 55554
rect 20959 55520 20993 55554
rect 23263 55520 23297 55554
rect 23551 55520 23585 55554
rect 24799 55520 24833 55554
rect 24991 55520 25025 55554
rect 39007 55520 39041 55554
rect 39199 55520 39233 55554
rect 39871 55520 39905 55554
rect 40927 55520 40961 55554
rect 45535 55520 45569 55554
rect 51967 55520 52001 55554
rect 55807 55520 55841 55554
rect 56575 55520 56609 55554
rect 57631 55520 57665 55554
rect 39679 55446 39713 55480
rect 1951 55372 1985 55406
rect 7327 55372 7361 55406
rect 8959 55372 8993 55406
rect 17407 55372 17441 55406
rect 20095 55372 20129 55406
rect 20767 55372 20801 55406
rect 45343 55372 45377 55406
rect 45823 55372 45857 55406
rect 55615 55372 55649 55406
rect 56287 55372 56321 55406
rect 57343 55372 57377 55406
rect 57919 55150 57953 55184
rect 42367 55002 42401 55036
rect 57631 54854 57665 54888
rect 57823 54854 57857 54888
rect 25663 54780 25697 54814
rect 7231 54706 7265 54740
rect 7519 54706 7553 54740
rect 20191 54706 20225 54740
rect 20479 54706 20513 54740
rect 22399 54706 22433 54740
rect 22783 54706 22817 54740
rect 57919 54336 57953 54370
rect 57823 54188 57857 54222
rect 57631 54040 57665 54074
rect 58111 54040 58145 54074
rect 57919 53818 57953 53852
rect 57823 53522 57857 53556
rect 57631 53374 57665 53408
rect 58111 53374 58145 53408
rect 29983 53004 30017 53038
rect 1759 52856 1793 52890
rect 2047 52856 2081 52890
rect 51487 52856 51521 52890
rect 2527 51524 2561 51558
rect 2815 51524 2849 51558
rect 43903 51376 43937 51410
rect 12511 51154 12545 51188
rect 31999 50858 32033 50892
rect 37375 50710 37409 50744
rect 37663 50710 37697 50744
rect 56959 50710 56993 50744
rect 57151 50710 57185 50744
rect 4159 50414 4193 50448
rect 40927 50192 40961 50226
rect 40831 50044 40865 50078
rect 6271 49526 6305 49560
rect 44863 49378 44897 49412
rect 45247 49378 45281 49412
rect 48031 49378 48065 49412
rect 48127 49378 48161 49412
rect 7231 49008 7265 49042
rect 1759 48860 1793 48894
rect 41407 48860 41441 48894
rect 41599 48860 41633 48894
rect 1951 48712 1985 48746
rect 28543 48712 28577 48746
rect 4255 48046 4289 48080
rect 4543 48046 4577 48080
rect 58015 48046 58049 48080
rect 17407 47602 17441 47636
rect 17695 47602 17729 47636
rect 23551 47528 23585 47562
rect 31711 46862 31745 46896
rect 13663 46788 13697 46822
rect 13951 46788 13985 46822
rect 4543 46714 4577 46748
rect 4831 46714 4865 46748
rect 15391 46714 15425 46748
rect 15679 46714 15713 46748
rect 45343 46714 45377 46748
rect 45439 46714 45473 46748
rect 28255 46196 28289 46230
rect 27967 46122 28001 46156
rect 40255 46048 40289 46082
rect 38911 44864 38945 44898
rect 39103 44864 39137 44898
rect 46783 44050 46817 44084
rect 46975 44050 47009 44084
rect 47743 44050 47777 44084
rect 47839 44050 47873 44084
rect 37087 43606 37121 43640
rect 37375 43606 37409 43640
rect 13759 43532 13793 43566
rect 38623 43532 38657 43566
rect 52063 43532 52097 43566
rect 38431 43384 38465 43418
rect 10975 42718 11009 42752
rect 11263 42718 11297 42752
rect 25951 42718 25985 42752
rect 26239 42718 26273 42752
rect 45247 42718 45281 42752
rect 45439 42718 45473 42752
rect 16255 42200 16289 42234
rect 16543 42200 16577 42234
rect 48223 42200 48257 42234
rect 39007 41756 39041 41790
rect 33247 41386 33281 41420
rect 33439 41386 33473 41420
rect 33535 40942 33569 40976
rect 1855 40868 1889 40902
rect 2047 40868 2081 40902
rect 34111 40868 34145 40902
rect 33919 40720 33953 40754
rect 44959 40498 44993 40532
rect 26623 40054 26657 40088
rect 26815 40054 26849 40088
rect 57343 40054 57377 40088
rect 57535 40054 57569 40088
rect 57823 39536 57857 39570
rect 57727 39388 57761 39422
rect 30751 39166 30785 39200
rect 26623 38870 26657 38904
rect 10399 38722 10433 38756
rect 10687 38722 10721 38756
rect 24127 38722 24161 38756
rect 24415 38722 24449 38756
rect 31327 38722 31361 38756
rect 31615 38722 31649 38756
rect 57631 38722 57665 38756
rect 57823 38722 57857 38756
rect 34111 38204 34145 38238
rect 34399 38204 34433 38238
rect 54655 38204 54689 38238
rect 55423 38204 55457 38238
rect 55231 38130 55265 38164
rect 34111 38056 34145 38090
rect 34207 38056 34241 38090
rect 5023 37390 5057 37424
rect 5791 37390 5825 37424
rect 6079 37390 6113 37424
rect 43327 37390 43361 37424
rect 14623 36872 14657 36906
rect 14911 36872 14945 36906
rect 24031 36872 24065 36906
rect 23839 36724 23873 36758
rect 9823 36206 9857 36240
rect 16927 36132 16961 36166
rect 17119 36132 17153 36166
rect 20671 36058 20705 36092
rect 20863 36058 20897 36092
rect 44383 36058 44417 36092
rect 44575 36058 44609 36092
rect 10687 35540 10721 35574
rect 10879 35540 10913 35574
rect 20383 35540 20417 35574
rect 20671 35540 20705 35574
rect 21055 35540 21089 35574
rect 21343 35540 21377 35574
rect 52639 35540 52673 35574
rect 52831 35540 52865 35574
rect 56671 35540 56705 35574
rect 56575 35392 56609 35426
rect 30943 34800 30977 34834
rect 15583 34726 15617 34760
rect 15871 34726 15905 34760
rect 31423 34726 31457 34760
rect 31519 34726 31553 34760
rect 53119 34726 53153 34760
rect 53215 34726 53249 34760
rect 57055 34726 57089 34760
rect 57247 34726 57281 34760
rect 28255 34208 28289 34242
rect 58015 34208 58049 34242
rect 26719 33468 26753 33502
rect 16831 33394 16865 33428
rect 35935 33394 35969 33428
rect 36223 33394 36257 33428
rect 39583 32728 39617 32762
rect 32575 32210 32609 32244
rect 26239 32136 26273 32170
rect 5887 32062 5921 32096
rect 21631 32062 21665 32096
rect 27391 32062 27425 32096
rect 32575 32062 32609 32096
rect 52831 31692 52865 31726
rect 20575 30878 20609 30912
rect 53407 30804 53441 30838
rect 6943 30730 6977 30764
rect 19039 30730 19073 30764
rect 52063 30730 52097 30764
rect 55327 30730 55361 30764
rect 38911 30360 38945 30394
rect 4351 30286 4385 30320
rect 4639 30286 4673 30320
rect 36415 29472 36449 29506
rect 6271 29398 6305 29432
rect 37087 29398 37121 29432
rect 18463 28880 18497 28914
rect 37567 28880 37601 28914
rect 10975 28066 11009 28100
rect 11167 28066 11201 28100
rect 36223 28066 36257 28100
rect 24223 27844 24257 27878
rect 24319 27844 24353 27878
rect 18271 27622 18305 27656
rect 56383 27548 56417 27582
rect 57055 27548 57089 27582
rect 27967 27400 28001 27434
rect 28063 27400 28097 27434
rect 18751 26956 18785 26990
rect 18943 26956 18977 26990
rect 15103 26734 15137 26768
rect 16639 26734 16673 26768
rect 57343 25402 57377 25436
rect 46783 25180 46817 25214
rect 46975 25180 47009 25214
rect 54271 24958 54305 24992
rect 54463 24958 54497 24992
rect 25471 24884 25505 24918
rect 50527 24884 50561 24918
rect 55327 24884 55361 24918
rect 42655 24070 42689 24104
rect 42847 24070 42881 24104
rect 38815 22812 38849 22846
rect 13567 22738 13601 22772
rect 17791 22738 17825 22772
rect 26911 22738 26945 22772
rect 30943 22738 30977 22772
rect 41119 22738 41153 22772
rect 41311 22738 41345 22772
rect 8383 22442 8417 22476
rect 27199 22442 27233 22476
rect 15583 22220 15617 22254
rect 26815 22220 26849 22254
rect 27103 22220 27137 22254
rect 27199 22220 27233 22254
rect 8095 22146 8129 22180
rect 7615 21184 7649 21218
rect 33535 20888 33569 20922
rect 34399 20888 34433 20922
rect 50719 20888 50753 20922
rect 50911 20888 50945 20922
rect 34399 20740 34433 20774
rect 22015 20518 22049 20552
rect 22207 20518 22241 20552
rect 9823 20074 9857 20108
rect 45151 20074 45185 20108
rect 49663 20074 49697 20108
rect 7615 19852 7649 19886
rect 8191 19852 8225 19886
rect 8383 19778 8417 19812
rect 12127 19630 12161 19664
rect 12415 19630 12449 19664
rect 18943 19556 18977 19590
rect 30559 19556 30593 19590
rect 7711 18742 7745 18776
rect 44959 18742 44993 18776
rect 8383 18520 8417 18554
rect 8575 18446 8609 18480
rect 18271 18224 18305 18258
rect 30847 18224 30881 18258
rect 42847 18224 42881 18258
rect 46015 18224 46049 18258
rect 7615 18076 7649 18110
rect 45823 18076 45857 18110
rect 22303 17558 22337 17592
rect 22495 17558 22529 17592
rect 23359 17410 23393 17444
rect 7615 17188 7649 17222
rect 7903 17188 7937 17222
rect 8191 17188 8225 17222
rect 35359 16966 35393 17000
rect 35551 16966 35585 17000
rect 19423 16892 19457 16926
rect 44191 16152 44225 16186
rect 44479 16152 44513 16186
rect 49567 16078 49601 16112
rect 35071 15856 35105 15890
rect 35263 15856 35297 15890
rect 7615 15782 7649 15816
rect 36703 15190 36737 15224
rect 36991 15190 37025 15224
rect 7903 14746 7937 14780
rect 20479 14746 20513 14780
rect 21151 14746 21185 14780
rect 52639 14746 52673 14780
rect 36607 14524 36641 14558
rect 36799 14524 36833 14558
rect 7615 14376 7649 14410
rect 3007 13562 3041 13596
rect 3295 13562 3329 13596
rect 7519 13488 7553 13522
rect 7807 13488 7841 13522
rect 6847 13414 6881 13448
rect 11455 13414 11489 13448
rect 7615 13118 7649 13152
rect 29023 12970 29057 13004
rect 57919 12970 57953 13004
rect 57343 12526 57377 12560
rect 57631 12378 57665 12412
rect 57919 12378 57953 12412
rect 57727 12230 57761 12264
rect 20383 12082 20417 12116
rect 31039 12082 31073 12116
rect 44575 12082 44609 12116
rect 2047 11860 2081 11894
rect 2335 11860 2369 11894
rect 55519 11860 55553 11894
rect 7615 11786 7649 11820
rect 33919 11712 33953 11746
rect 39775 11712 39809 11746
rect 40063 11712 40097 11746
rect 55711 11712 55745 11746
rect 56575 11712 56609 11746
rect 56959 11638 56993 11672
rect 57247 11638 57281 11672
rect 3007 11564 3041 11598
rect 56191 11564 56225 11598
rect 56479 11564 56513 11598
rect 56767 11564 56801 11598
rect 57343 11416 57377 11450
rect 56095 11046 56129 11080
rect 57055 10972 57089 11006
rect 57343 10972 57377 11006
rect 55999 10898 56033 10932
rect 57247 10898 57281 10932
rect 41887 10824 41921 10858
rect 2911 10750 2945 10784
rect 3199 10750 3233 10784
rect 44767 10750 44801 10784
rect 54751 10750 54785 10784
rect 56959 10454 56993 10488
rect 57055 10454 57089 10488
rect 54847 10380 54881 10414
rect 55039 10380 55073 10414
rect 55135 10380 55169 10414
rect 55519 10306 55553 10340
rect 55807 10306 55841 10340
rect 56095 10306 56129 10340
rect 56959 10306 56993 10340
rect 57343 10306 57377 10340
rect 17695 10232 17729 10266
rect 56671 10232 56705 10266
rect 7615 10084 7649 10118
rect 55903 10084 55937 10118
rect 56575 10084 56609 10118
rect 57439 10084 57473 10118
rect 54847 9862 54881 9896
rect 54463 9714 54497 9748
rect 55135 9714 55169 9748
rect 55999 9640 56033 9674
rect 57631 9640 57665 9674
rect 54367 9566 54401 9600
rect 55231 9566 55265 9600
rect 55903 9566 55937 9600
rect 46687 9492 46721 9526
rect 46975 9492 47009 9526
rect 53119 9418 53153 9452
rect 53791 9418 53825 9452
rect 3103 9196 3137 9230
rect 7615 9122 7649 9156
rect 7711 9122 7745 9156
rect 8479 9122 8513 9156
rect 37471 9122 37505 9156
rect 30079 9048 30113 9082
rect 30367 9048 30401 9082
rect 36511 9048 36545 9082
rect 36799 9048 36833 9082
rect 54655 9048 54689 9082
rect 49375 8974 49409 9008
rect 53327 8974 53361 9008
rect 56575 8974 56609 9008
rect 57247 8974 57281 9008
rect 42751 8900 42785 8934
rect 44095 8900 44129 8934
rect 53407 8900 53441 8934
rect 55423 8900 55457 8934
rect 42751 8752 42785 8786
rect 54559 8752 54593 8786
rect 55327 8752 55361 8786
rect 2047 8530 2081 8564
rect 13567 8530 13601 8564
rect 14527 8530 14561 8564
rect 42079 8530 42113 8564
rect 48607 8530 48641 8564
rect 52447 8530 52481 8564
rect 1759 8382 1793 8416
rect 3007 8382 3041 8416
rect 3295 8382 3329 8416
rect 4255 8382 4289 8416
rect 4543 8382 4577 8416
rect 10591 8382 10625 8416
rect 11071 8382 11105 8416
rect 11359 8382 11393 8416
rect 11839 8382 11873 8416
rect 12127 8382 12161 8416
rect 12895 8382 12929 8416
rect 13663 8382 13697 8416
rect 9823 8308 9857 8342
rect 1663 8234 1697 8268
rect 2431 8234 2465 8268
rect 2527 8234 2561 8268
rect 3199 8234 3233 8268
rect 4447 8234 4481 8268
rect 7807 8234 7841 8268
rect 7903 8234 7937 8268
rect 9743 8234 9777 8268
rect 10495 8234 10529 8268
rect 11263 8234 11297 8268
rect 12031 8234 12065 8268
rect 12799 8234 12833 8268
rect 39487 8456 39521 8490
rect 34111 8382 34145 8416
rect 34399 8382 34433 8416
rect 35071 8382 35105 8416
rect 39679 8382 39713 8416
rect 42175 8382 42209 8416
rect 48223 8382 48257 8416
rect 52543 8382 52577 8416
rect 53311 8382 53345 8416
rect 16255 8308 16289 8342
rect 17023 8308 17057 8342
rect 49759 8308 49793 8342
rect 54079 8308 54113 8342
rect 55231 8308 55265 8342
rect 55999 8308 56033 8342
rect 57151 8308 57185 8342
rect 16159 8234 16193 8268
rect 16927 8234 16961 8268
rect 48127 8234 48161 8268
rect 48895 8234 48929 8268
rect 48991 8234 49025 8268
rect 49663 8234 49697 8268
rect 53215 8234 53249 8268
rect 53983 8234 54017 8268
rect 33631 8160 33665 8194
rect 6175 8086 6209 8120
rect 6943 8086 6977 8120
rect 9535 8086 9569 8120
rect 14527 8086 14561 8120
rect 17791 8086 17825 8120
rect 22111 8086 22145 8120
rect 25951 8086 25985 8120
rect 2911 7864 2945 7898
rect 29023 7864 29057 7898
rect 36511 7864 36545 7898
rect 39199 7864 39233 7898
rect 40063 7864 40097 7898
rect 46111 7864 46145 7898
rect 51487 7864 51521 7898
rect 7615 7790 7649 7824
rect 8767 7790 8801 7824
rect 24319 7790 24353 7824
rect 25087 7790 25121 7824
rect 2527 7716 2561 7750
rect 3295 7716 3329 7750
rect 4063 7716 4097 7750
rect 4831 7716 4865 7750
rect 5311 7716 5345 7750
rect 5599 7716 5633 7750
rect 10207 7716 10241 7750
rect 10975 7716 11009 7750
rect 12415 7716 12449 7750
rect 13855 7716 13889 7750
rect 15583 7716 15617 7750
rect 15871 7716 15905 7750
rect 20959 7716 20993 7750
rect 23647 7716 23681 7750
rect 23935 7716 23969 7750
rect 24607 7716 24641 7750
rect 25375 7716 25409 7750
rect 25471 7716 25505 7750
rect 25951 7716 25985 7750
rect 26143 7716 26177 7750
rect 29311 7716 29345 7750
rect 30175 7716 30209 7750
rect 33823 7716 33857 7750
rect 34591 7716 34625 7750
rect 35359 7716 35393 7750
rect 36127 7716 36161 7750
rect 36799 7716 36833 7750
rect 39583 7716 39617 7750
rect 41023 7716 41057 7750
rect 41119 7716 41153 7750
rect 42655 7716 42689 7750
rect 44095 7716 44129 7750
rect 44863 7716 44897 7750
rect 45631 7716 45665 7750
rect 46303 7716 46337 7750
rect 46399 7716 46433 7750
rect 47071 7716 47105 7750
rect 49375 7716 49409 7750
rect 50143 7716 50177 7750
rect 51775 7716 51809 7750
rect 52639 7716 52673 7750
rect 53407 7716 53441 7750
rect 1567 7642 1601 7676
rect 8383 7642 8417 7676
rect 9439 7642 9473 7676
rect 12895 7642 12929 7676
rect 13183 7642 13217 7676
rect 28351 7642 28385 7676
rect 39487 7642 39521 7676
rect 55135 7642 55169 7676
rect 55807 7642 55841 7676
rect 56575 7642 56609 7676
rect 57343 7642 57377 7676
rect 7135 7568 7169 7602
rect 13951 7568 13985 7602
rect 15199 7568 15233 7602
rect 21727 7568 21761 7602
rect 23263 7568 23297 7602
rect 27007 7568 27041 7602
rect 31231 7568 31265 7602
rect 32383 7568 32417 7602
rect 38815 7568 38849 7602
rect 40255 7568 40289 7602
rect 41887 7568 41921 7602
rect 46879 7568 46913 7602
rect 47167 7568 47201 7602
rect 47935 7568 47969 7602
rect 51103 7568 51137 7602
rect 10127 7494 10161 7528
rect 2431 7420 2465 7454
rect 3199 7420 3233 7454
rect 3967 7420 4001 7454
rect 4735 7420 4769 7454
rect 5503 7420 5537 7454
rect 9343 7420 9377 7454
rect 10879 7420 10913 7454
rect 12319 7420 12353 7454
rect 13087 7420 13121 7454
rect 15775 7420 15809 7454
rect 20863 7420 20897 7454
rect 23839 7420 23873 7454
rect 24703 7420 24737 7454
rect 26239 7420 26273 7454
rect 26911 7420 26945 7454
rect 28255 7420 28289 7454
rect 29407 7420 29441 7454
rect 30079 7420 30113 7454
rect 31135 7420 31169 7454
rect 33727 7420 33761 7454
rect 34495 7420 34529 7454
rect 35263 7420 35297 7454
rect 36031 7420 36065 7454
rect 36895 7420 36929 7454
rect 38719 7420 38753 7454
rect 40351 7420 40385 7454
rect 41791 7420 41825 7454
rect 42559 7420 42593 7454
rect 43999 7420 44033 7454
rect 44767 7420 44801 7454
rect 45535 7420 45569 7454
rect 47839 7420 47873 7454
rect 49279 7420 49313 7454
rect 50047 7420 50081 7454
rect 51007 7420 51041 7454
rect 51871 7420 51905 7454
rect 52543 7420 52577 7454
rect 53311 7420 53345 7454
rect 17791 7124 17825 7158
rect 19999 7124 20033 7158
rect 22303 7124 22337 7158
rect 23167 7124 23201 7158
rect 23839 7124 23873 7158
rect 26047 7124 26081 7158
rect 26815 7124 26849 7158
rect 27583 7124 27617 7158
rect 30559 7124 30593 7158
rect 38143 7124 38177 7158
rect 39487 7124 39521 7158
rect 39679 7124 39713 7158
rect 41887 7124 41921 7158
rect 42255 7124 42289 7158
rect 44959 7124 44993 7158
rect 4255 7050 4289 7084
rect 4543 7050 4577 7084
rect 6559 7050 6593 7084
rect 6847 7050 6881 7084
rect 7615 7050 7649 7084
rect 8383 7050 8417 7084
rect 9823 7050 9857 7084
rect 10303 7050 10337 7084
rect 10591 7050 10625 7084
rect 13663 7050 13697 7084
rect 14815 7050 14849 7084
rect 15007 7050 15041 7084
rect 15871 7050 15905 7084
rect 16351 7050 16385 7084
rect 16639 7050 16673 7084
rect 17311 7050 17345 7084
rect 18079 7050 18113 7084
rect 18847 7050 18881 7084
rect 20287 7050 20321 7084
rect 21151 7050 21185 7084
rect 21631 7050 21665 7084
rect 21919 7050 21953 7084
rect 22687 7050 22721 7084
rect 23359 7050 23393 7084
rect 24127 7050 24161 7084
rect 25375 7050 25409 7084
rect 25663 7050 25697 7084
rect 26431 7050 26465 7084
rect 27103 7050 27137 7084
rect 27967 7050 28001 7084
rect 29503 7050 29537 7084
rect 30847 7050 30881 7084
rect 31423 7050 31457 7084
rect 31615 7050 31649 7084
rect 32479 7050 32513 7084
rect 34015 7050 34049 7084
rect 36223 7050 36257 7084
rect 36991 7050 37025 7084
rect 37759 7050 37793 7084
rect 38431 7050 38465 7084
rect 1663 6976 1697 7010
rect 2527 6976 2561 7010
rect 6079 6976 6113 7010
rect 11263 6976 11297 7010
rect 12703 6976 12737 7010
rect 28735 6976 28769 7010
rect 33247 6976 33281 7010
rect 39295 6976 39329 7010
rect 39967 7050 40001 7084
rect 41503 7050 41537 7084
rect 43039 7050 43073 7084
rect 43711 7050 43745 7084
rect 44191 7050 44225 7084
rect 44479 7050 44513 7084
rect 45247 7050 45281 7084
rect 46783 7050 46817 7084
rect 48319 7050 48353 7084
rect 49087 7050 49121 7084
rect 50335 7050 50369 7084
rect 52063 7050 52097 7084
rect 52831 7050 52865 7084
rect 42175 6976 42209 7010
rect 47551 6976 47585 7010
rect 54079 6976 54113 7010
rect 54751 6976 54785 7010
rect 55519 6976 55553 7010
rect 57823 6976 57857 7010
rect 4447 6902 4481 6936
rect 5215 6902 5249 6936
rect 5311 6902 5345 6936
rect 5983 6902 6017 6936
rect 6751 6902 6785 6936
rect 7519 6902 7553 6936
rect 8287 6902 8321 6936
rect 9727 6902 9761 6936
rect 10495 6902 10529 6936
rect 13567 6902 13601 6936
rect 15103 6902 15137 6936
rect 15775 6902 15809 6936
rect 17215 6902 17249 6936
rect 17983 6902 18017 6936
rect 18751 6902 18785 6936
rect 20383 6902 20417 6936
rect 21055 6902 21089 6936
rect 21823 6902 21857 6936
rect 22591 6902 22625 6936
rect 23455 6902 23489 6936
rect 24223 6902 24257 6936
rect 25567 6902 25601 6936
rect 26335 6902 26369 6936
rect 27199 6902 27233 6936
rect 27871 6902 27905 6936
rect 28639 6902 28673 6936
rect 29407 6902 29441 6936
rect 30943 6902 30977 6936
rect 31711 6902 31745 6936
rect 32383 6902 32417 6936
rect 33151 6902 33185 6936
rect 33919 6902 33953 6936
rect 34687 6902 34721 6936
rect 34783 6902 34817 6936
rect 36127 6902 36161 6936
rect 36895 6902 36929 6936
rect 37663 6902 37697 6936
rect 38527 6902 38561 6936
rect 39199 6902 39233 6936
rect 39487 6902 39521 6936
rect 40063 6902 40097 6936
rect 41407 6902 41441 6936
rect 42943 6902 42977 6936
rect 43807 6902 43841 6936
rect 44575 6902 44609 6936
rect 45343 6902 45377 6936
rect 46687 6902 46721 6936
rect 47455 6902 47489 6936
rect 48223 6902 48257 6936
rect 48991 6902 49025 6936
rect 50239 6902 50273 6936
rect 51967 6902 52001 6936
rect 52735 6902 52769 6936
rect 43423 6754 43457 6788
rect 7615 6458 7649 6492
rect 7711 6458 7745 6492
rect 8479 6532 8513 6566
rect 15103 6532 15137 6566
rect 15871 6532 15905 6566
rect 20479 6532 20513 6566
rect 24127 6532 24161 6566
rect 27871 6532 27905 6566
rect 33151 6532 33185 6566
rect 34687 6532 34721 6566
rect 35839 6532 35873 6566
rect 5407 6384 5441 6418
rect 5695 6384 5729 6418
rect 6847 6384 6881 6418
rect 7135 6384 7169 6418
rect 13951 6384 13985 6418
rect 14719 6384 14753 6418
rect 15487 6384 15521 6418
rect 16159 6384 16193 6418
rect 16255 6384 16289 6418
rect 17407 6384 17441 6418
rect 17695 6384 17729 6418
rect 18175 6384 18209 6418
rect 18463 6384 18497 6418
rect 18943 6384 18977 6418
rect 19231 6384 19265 6418
rect 19999 6384 20033 6418
rect 20671 6384 20705 6418
rect 20767 6384 20801 6418
rect 21535 6384 21569 6418
rect 22975 6384 23009 6418
rect 23455 6384 23489 6418
rect 23647 6384 23681 6418
rect 24415 6384 24449 6418
rect 28159 6384 28193 6418
rect 28735 6384 28769 6418
rect 29023 6384 29057 6418
rect 33439 6384 33473 6418
rect 34303 6384 34337 6418
rect 34975 6384 35009 6418
rect 35071 6384 35105 6418
rect 37279 6384 37313 6418
rect 41023 6384 41057 6418
rect 41215 6384 41249 6418
rect 42847 6384 42881 6418
rect 44095 6384 44129 6418
rect 44863 6384 44897 6418
rect 50623 6384 50657 6418
rect 50815 6384 50849 6418
rect 51391 6384 51425 6418
rect 51583 6384 51617 6418
rect 1567 6310 1601 6344
rect 2335 6310 2369 6344
rect 3199 6310 3233 6344
rect 3967 6310 4001 6344
rect 4735 6310 4769 6344
rect 9439 6310 9473 6344
rect 10207 6310 10241 6344
rect 10975 6310 11009 6344
rect 12223 6310 12257 6344
rect 12991 6310 13025 6344
rect 25663 6310 25697 6344
rect 26815 6310 26849 6344
rect 29695 6310 29729 6344
rect 31231 6310 31265 6344
rect 36319 6310 36353 6344
rect 38911 6310 38945 6344
rect 40351 6310 40385 6344
rect 41887 6310 41921 6344
rect 45535 6310 45569 6344
rect 46975 6310 47009 6344
rect 47743 6310 47777 6344
rect 49183 6310 49217 6344
rect 49951 6310 49985 6344
rect 53311 6310 53345 6344
rect 54463 6310 54497 6344
rect 55231 6310 55265 6344
rect 55999 6310 56033 6344
rect 57055 6310 57089 6344
rect 57823 6310 57857 6344
rect 30655 6236 30689 6270
rect 32191 6236 32225 6270
rect 37183 6236 37217 6270
rect 52447 6236 52481 6270
rect 5599 6088 5633 6122
rect 7039 6088 7073 6122
rect 13855 6088 13889 6122
rect 14623 6088 14657 6122
rect 15391 6088 15425 6122
rect 17599 6088 17633 6122
rect 18367 6088 18401 6122
rect 19135 6088 19169 6122
rect 19903 6088 19937 6122
rect 21439 6088 21473 6122
rect 22879 6088 22913 6122
rect 23743 6088 23777 6122
rect 24511 6088 24545 6122
rect 28255 6088 28289 6122
rect 28927 6088 28961 6122
rect 30559 6088 30593 6122
rect 32095 6088 32129 6122
rect 33535 6088 33569 6122
rect 34207 6088 34241 6122
rect 36895 6088 36929 6122
rect 41311 6088 41345 6122
rect 42751 6088 42785 6122
rect 43999 6088 44033 6122
rect 44767 6088 44801 6122
rect 50911 6088 50945 6122
rect 51679 6088 51713 6122
rect 52351 6088 52385 6122
rect 5791 5718 5825 5752
rect 5983 5718 6017 5752
rect 11551 5718 11585 5752
rect 1567 5644 1601 5678
rect 2911 5644 2945 5678
rect 4447 5644 4481 5678
rect 5119 5644 5153 5678
rect 6847 5644 6881 5678
rect 7615 5644 7649 5678
rect 8383 5644 8417 5678
rect 9631 5644 9665 5678
rect 10399 5644 10433 5678
rect 11167 5644 11201 5678
rect 6079 5570 6113 5604
rect 12607 5644 12641 5678
rect 13375 5644 13409 5678
rect 15007 5644 15041 5678
rect 15871 5644 15905 5678
rect 16543 5644 16577 5678
rect 17311 5644 17345 5678
rect 18751 5644 18785 5678
rect 20191 5644 20225 5678
rect 20959 5644 20993 5678
rect 21631 5644 21665 5678
rect 21727 5644 21761 5678
rect 22495 5644 22529 5678
rect 23263 5644 23297 5678
rect 24031 5644 24065 5678
rect 25471 5644 25505 5678
rect 26239 5644 26273 5678
rect 26623 5644 26657 5678
rect 27007 5644 27041 5678
rect 27775 5644 27809 5678
rect 28543 5644 28577 5678
rect 29311 5644 29345 5678
rect 30751 5644 30785 5678
rect 31519 5644 31553 5678
rect 32287 5644 32321 5678
rect 33151 5644 33185 5678
rect 33823 5644 33857 5678
rect 34687 5644 34721 5678
rect 36031 5644 36065 5678
rect 36799 5644 36833 5678
rect 37567 5644 37601 5678
rect 38335 5644 38369 5678
rect 39103 5644 39137 5678
rect 39871 5644 39905 5678
rect 41311 5644 41345 5678
rect 42079 5644 42113 5678
rect 42847 5644 42881 5678
rect 43615 5644 43649 5678
rect 44383 5644 44417 5678
rect 45151 5644 45185 5678
rect 46591 5644 46625 5678
rect 47359 5644 47393 5678
rect 48127 5644 48161 5678
rect 48991 5644 49025 5678
rect 49663 5644 49697 5678
rect 50527 5644 50561 5678
rect 52159 5644 52193 5678
rect 52927 5644 52961 5678
rect 53695 5644 53729 5678
rect 54463 5644 54497 5678
rect 55999 5644 56033 5678
rect 57439 5644 57473 5678
rect 21631 5496 21665 5530
rect 26623 5496 26657 5530
rect 11551 5422 11585 5456
rect 55423 5422 55457 5456
rect 7519 5200 7553 5234
rect 7711 5200 7745 5234
rect 8479 5200 8513 5234
rect 58015 5200 58049 5234
rect 1567 4978 1601 5012
rect 2335 4978 2369 5012
rect 3103 4978 3137 5012
rect 4159 4978 4193 5012
rect 5407 4978 5441 5012
rect 6943 4978 6977 5012
rect 9247 4978 9281 5012
rect 10015 4978 10049 5012
rect 10783 4978 10817 5012
rect 12223 4978 12257 5012
rect 12991 4978 13025 5012
rect 13951 4978 13985 5012
rect 14719 4978 14753 5012
rect 15487 4978 15521 5012
rect 16351 4978 16385 5012
rect 17503 4978 17537 5012
rect 18271 4978 18305 5012
rect 19039 4978 19073 5012
rect 19807 4978 19841 5012
rect 20671 4978 20705 5012
rect 21343 4978 21377 5012
rect 22783 4978 22817 5012
rect 23551 4978 23585 5012
rect 24319 4978 24353 5012
rect 25087 4978 25121 5012
rect 25855 4978 25889 5012
rect 26623 4978 26657 5012
rect 28063 4978 28097 5012
rect 28927 4978 28961 5012
rect 29599 4978 29633 5012
rect 30367 4978 30401 5012
rect 31135 4978 31169 5012
rect 31903 4978 31937 5012
rect 33343 4978 33377 5012
rect 34111 4978 34145 5012
rect 34879 4978 34913 5012
rect 35647 4978 35681 5012
rect 36415 4978 36449 5012
rect 37183 4978 37217 5012
rect 38623 4978 38657 5012
rect 39391 4978 39425 5012
rect 40159 4978 40193 5012
rect 40927 4978 40961 5012
rect 41695 4978 41729 5012
rect 42463 4978 42497 5012
rect 43903 4978 43937 5012
rect 44767 4978 44801 5012
rect 45439 4978 45473 5012
rect 46207 4978 46241 5012
rect 46975 4978 47009 5012
rect 47743 4978 47777 5012
rect 49375 4978 49409 5012
rect 50431 4978 50465 5012
rect 51103 4978 51137 5012
rect 51871 4978 51905 5012
rect 52639 4978 52673 5012
rect 54463 4978 54497 5012
rect 55615 4978 55649 5012
rect 56383 4978 56417 5012
rect 57055 4978 57089 5012
rect 41119 4386 41153 4420
rect 41311 4386 41345 4420
rect 1567 4312 1601 4346
rect 2335 4312 2369 4346
rect 3103 4312 3137 4346
rect 4351 4312 4385 4346
rect 5119 4312 5153 4346
rect 5887 4312 5921 4346
rect 6655 4312 6689 4346
rect 7423 4312 7457 4346
rect 8191 4312 8225 4346
rect 9631 4312 9665 4346
rect 10399 4312 10433 4346
rect 11167 4312 11201 4346
rect 11935 4312 11969 4346
rect 12703 4312 12737 4346
rect 13567 4312 13601 4346
rect 15487 4312 15521 4346
rect 16255 4312 16289 4346
rect 17023 4312 17057 4346
rect 17791 4312 17825 4346
rect 18559 4312 18593 4346
rect 20287 4312 20321 4346
rect 21055 4312 21089 4346
rect 21823 4312 21857 4346
rect 23263 4312 23297 4346
rect 24031 4312 24065 4346
rect 25471 4312 25505 4346
rect 26239 4312 26273 4346
rect 27007 4312 27041 4346
rect 28351 4312 28385 4346
rect 29119 4312 29153 4346
rect 30943 4312 30977 4346
rect 31711 4312 31745 4346
rect 32767 4312 32801 4346
rect 33919 4312 33953 4346
rect 34687 4312 34721 4346
rect 36031 4312 36065 4346
rect 36799 4312 36833 4346
rect 37567 4312 37601 4346
rect 39007 4312 39041 4346
rect 39775 4312 39809 4346
rect 41983 4312 42017 4346
rect 42751 4312 42785 4346
rect 43519 4312 43553 4346
rect 44959 4312 44993 4346
rect 46783 4312 46817 4346
rect 47551 4312 47585 4346
rect 48319 4312 48353 4346
rect 49087 4312 49121 4346
rect 49855 4312 49889 4346
rect 50623 4312 50657 4346
rect 51871 4312 51905 4346
rect 52639 4312 52673 4346
rect 53407 4312 53441 4346
rect 54175 4312 54209 4346
rect 55615 4312 55649 4346
rect 57151 4312 57185 4346
rect 55135 4238 55169 4272
rect 44479 4164 44513 4198
rect 1567 3646 1601 3680
rect 2335 3646 2369 3680
rect 3103 3646 3137 3680
rect 3871 3646 3905 3680
rect 4639 3646 4673 3680
rect 5599 3646 5633 3680
rect 6943 3646 6977 3680
rect 7711 3646 7745 3680
rect 8479 3646 8513 3680
rect 9247 3646 9281 3680
rect 10015 3646 10049 3680
rect 10783 3646 10817 3680
rect 12991 3646 13025 3680
rect 13663 3646 13697 3680
rect 14431 3646 14465 3680
rect 15199 3646 15233 3680
rect 15967 3646 16001 3680
rect 17503 3646 17537 3680
rect 18271 3646 18305 3680
rect 19039 3646 19073 3680
rect 19807 3646 19841 3680
rect 20575 3646 20609 3680
rect 21343 3646 21377 3680
rect 22783 3646 22817 3680
rect 23551 3646 23585 3680
rect 24319 3646 24353 3680
rect 25087 3646 25121 3680
rect 25855 3646 25889 3680
rect 26623 3646 26657 3680
rect 28063 3646 28097 3680
rect 28831 3646 28865 3680
rect 29599 3646 29633 3680
rect 30367 3646 30401 3680
rect 31135 3646 31169 3680
rect 31903 3646 31937 3680
rect 33343 3646 33377 3680
rect 34111 3646 34145 3680
rect 34879 3646 34913 3680
rect 35647 3646 35681 3680
rect 36415 3646 36449 3680
rect 37183 3646 37217 3680
rect 38623 3646 38657 3680
rect 39391 3646 39425 3680
rect 40159 3646 40193 3680
rect 40927 3646 40961 3680
rect 41695 3646 41729 3680
rect 42463 3646 42497 3680
rect 43903 3646 43937 3680
rect 44671 3646 44705 3680
rect 45439 3646 45473 3680
rect 46207 3646 46241 3680
rect 46975 3646 47009 3680
rect 47743 3646 47777 3680
rect 49183 3646 49217 3680
rect 50527 3646 50561 3680
rect 51199 3646 51233 3680
rect 51967 3646 52001 3680
rect 52735 3646 52769 3680
rect 54463 3646 54497 3680
rect 55231 3646 55265 3680
rect 55999 3646 56033 3680
rect 56767 3646 56801 3680
rect 57535 3646 57569 3680
rect 12127 3424 12161 3458
rect 12415 3424 12449 3458
rect 35359 3128 35393 3162
rect 13279 3054 13313 3088
rect 35647 3054 35681 3088
rect 41023 3054 41057 3088
rect 53119 3054 53153 3088
rect 1567 2980 1601 3014
rect 2335 2980 2369 3014
rect 3103 2980 3137 3014
rect 4927 2980 4961 3014
rect 5695 2980 5729 3014
rect 7039 2980 7073 3014
rect 7807 2980 7841 3014
rect 9727 2980 9761 3014
rect 10495 2980 10529 3014
rect 12991 2980 13025 3014
rect 13759 2980 13793 3014
rect 15103 2980 15137 3014
rect 16639 2980 16673 3014
rect 17791 2980 17825 3014
rect 18559 2980 18593 3014
rect 20479 2980 20513 3014
rect 21247 2980 21281 3014
rect 23167 2980 23201 3014
rect 23935 2980 23969 3014
rect 25855 2980 25889 3014
rect 26623 2980 26657 3014
rect 28543 2980 28577 3014
rect 29311 2980 29345 3014
rect 31231 2980 31265 3014
rect 31999 2980 32033 3014
rect 33919 2980 33953 3014
rect 34687 2980 34721 3014
rect 36607 2980 36641 3014
rect 37375 2980 37409 3014
rect 39295 2980 39329 3014
rect 40063 2980 40097 3014
rect 41983 2980 42017 3014
rect 42751 2980 42785 3014
rect 44671 2980 44705 3014
rect 45439 2980 45473 3014
rect 47359 2980 47393 3014
rect 48127 2980 48161 3014
rect 50047 2980 50081 3014
rect 50815 2980 50849 3014
rect 52735 2980 52769 3014
rect 53503 2980 53537 3014
rect 55423 2980 55457 3014
rect 56191 2980 56225 3014
rect 46399 2832 46433 2866
rect 51775 2832 51809 2866
rect 53119 2832 53153 2866
rect 8767 2758 8801 2792
rect 43711 2758 43745 2792
rect 49087 2758 49121 2792
<< metal1 >>
rect 1152 57302 58848 57324
rect 1152 57250 4294 57302
rect 4346 57250 4358 57302
rect 4410 57250 4422 57302
rect 4474 57250 4486 57302
rect 4538 57250 35014 57302
rect 35066 57250 35078 57302
rect 35130 57250 35142 57302
rect 35194 57250 35206 57302
rect 35258 57250 58848 57302
rect 1152 57228 58848 57250
rect 1744 56991 1750 57043
rect 1802 57031 1808 57043
rect 1802 57003 2846 57031
rect 1802 56991 1808 57003
rect 208 56917 214 56969
rect 266 56957 272 56969
rect 2818 56966 2846 57003
rect 3280 56991 3286 57043
rect 3338 57031 3344 57043
rect 3338 57003 5822 57031
rect 3338 56991 3344 57003
rect 1939 56960 1997 56966
rect 1939 56957 1951 56960
rect 266 56929 1951 56957
rect 266 56917 272 56929
rect 1939 56926 1951 56929
rect 1985 56926 1997 56960
rect 1939 56920 1997 56926
rect 2803 56960 2861 56966
rect 2803 56926 2815 56960
rect 2849 56926 2861 56960
rect 2803 56920 2861 56926
rect 4912 56917 4918 56969
rect 4970 56957 4976 56969
rect 5794 56966 5822 57003
rect 9616 56991 9622 57043
rect 9674 57031 9680 57043
rect 9907 57034 9965 57040
rect 9907 57031 9919 57034
rect 9674 57003 9919 57031
rect 9674 56991 9680 57003
rect 9907 57000 9919 57003
rect 9953 57000 9965 57034
rect 9907 56994 9965 57000
rect 11248 56991 11254 57043
rect 11306 57031 11312 57043
rect 13939 57034 13997 57040
rect 11306 57003 11486 57031
rect 11306 56991 11312 57003
rect 5299 56960 5357 56966
rect 5299 56957 5311 56960
rect 4970 56929 5311 56957
rect 4970 56917 4976 56929
rect 5299 56926 5311 56929
rect 5345 56926 5357 56960
rect 5299 56920 5357 56926
rect 5779 56960 5837 56966
rect 5779 56926 5791 56960
rect 5825 56926 5837 56960
rect 5779 56920 5837 56926
rect 6448 56917 6454 56969
rect 6506 56957 6512 56969
rect 7411 56960 7469 56966
rect 7411 56957 7423 56960
rect 6506 56929 7423 56957
rect 6506 56917 6512 56929
rect 7411 56926 7423 56929
rect 7457 56926 7469 56960
rect 8080 56957 8086 56969
rect 8041 56929 8086 56957
rect 7411 56920 7469 56926
rect 8080 56917 8086 56929
rect 8138 56917 8144 56969
rect 11458 56966 11486 57003
rect 13939 57000 13951 57034
rect 13985 57031 13997 57034
rect 16432 57031 16438 57043
rect 13985 57003 16438 57031
rect 13985 57000 13997 57003
rect 13939 56994 13997 57000
rect 16432 56991 16438 57003
rect 16490 56991 16496 57043
rect 18064 56991 18070 57043
rect 18122 57031 18128 57043
rect 21523 57034 21581 57040
rect 21523 57031 21535 57034
rect 18122 57003 21535 57031
rect 18122 56991 18128 57003
rect 21523 57000 21535 57003
rect 21569 57000 21581 57034
rect 21523 56994 21581 57000
rect 29104 56991 29110 57043
rect 29162 57031 29168 57043
rect 32659 57034 32717 57040
rect 32659 57031 32671 57034
rect 29162 57003 32671 57031
rect 29162 56991 29168 57003
rect 32659 57000 32671 57003
rect 32705 57000 32717 57034
rect 32659 56994 32717 57000
rect 11443 56960 11501 56966
rect 11443 56926 11455 56960
rect 11489 56926 11501 56960
rect 11443 56920 11501 56926
rect 12784 56917 12790 56969
rect 12842 56957 12848 56969
rect 13171 56960 13229 56966
rect 13171 56957 13183 56960
rect 12842 56929 13183 56957
rect 12842 56917 12848 56929
rect 13171 56926 13183 56929
rect 13217 56926 13229 56960
rect 13171 56920 13229 56926
rect 14416 56917 14422 56969
rect 14474 56957 14480 56969
rect 15091 56960 15149 56966
rect 15091 56957 15103 56960
rect 14474 56929 15103 56957
rect 14474 56917 14480 56929
rect 15091 56926 15103 56929
rect 15137 56926 15149 56960
rect 15091 56920 15149 56926
rect 15952 56917 15958 56969
rect 16010 56957 16016 56969
rect 16339 56960 16397 56966
rect 16339 56957 16351 56960
rect 16010 56929 16351 56957
rect 16010 56917 16016 56929
rect 16339 56926 16351 56929
rect 16385 56926 16397 56960
rect 16339 56920 16397 56926
rect 17488 56917 17494 56969
rect 17546 56957 17552 56969
rect 17779 56960 17837 56966
rect 17779 56957 17791 56960
rect 17546 56929 17791 56957
rect 17546 56917 17552 56929
rect 17779 56926 17791 56929
rect 17825 56926 17837 56960
rect 17779 56920 17837 56926
rect 19120 56917 19126 56969
rect 19178 56957 19184 56969
rect 19507 56960 19565 56966
rect 19507 56957 19519 56960
rect 19178 56929 19519 56957
rect 19178 56917 19184 56929
rect 19507 56926 19519 56929
rect 19553 56926 19565 56960
rect 20656 56957 20662 56969
rect 20617 56929 20662 56957
rect 19507 56920 19565 56926
rect 20656 56917 20662 56929
rect 20714 56917 20720 56969
rect 22288 56917 22294 56969
rect 22346 56957 22352 56969
rect 23539 56960 23597 56966
rect 23539 56957 23551 56960
rect 22346 56929 23551 56957
rect 22346 56917 22352 56929
rect 23539 56926 23551 56929
rect 23585 56926 23597 56960
rect 23539 56920 23597 56926
rect 23824 56917 23830 56969
rect 23882 56957 23888 56969
rect 24019 56960 24077 56966
rect 24019 56957 24031 56960
rect 23882 56929 24031 56957
rect 23882 56917 23888 56929
rect 24019 56926 24031 56929
rect 24065 56926 24077 56960
rect 24019 56920 24077 56926
rect 25456 56917 25462 56969
rect 25514 56957 25520 56969
rect 26227 56960 26285 56966
rect 26227 56957 26239 56960
rect 25514 56929 26239 56957
rect 25514 56917 25520 56929
rect 26227 56926 26239 56929
rect 26273 56926 26285 56960
rect 26992 56957 26998 56969
rect 26953 56929 26998 56957
rect 26227 56920 26285 56926
rect 26992 56917 26998 56929
rect 27050 56917 27056 56969
rect 28624 56917 28630 56969
rect 28682 56957 28688 56969
rect 29011 56960 29069 56966
rect 29011 56957 29023 56960
rect 28682 56929 29023 56957
rect 28682 56917 28688 56929
rect 29011 56926 29023 56929
rect 29057 56926 29069 56960
rect 29011 56920 29069 56926
rect 30067 56960 30125 56966
rect 30067 56926 30079 56960
rect 30113 56957 30125 56960
rect 30160 56957 30166 56969
rect 30113 56929 30166 56957
rect 30113 56926 30125 56929
rect 30067 56920 30125 56926
rect 30160 56917 30166 56929
rect 30218 56917 30224 56969
rect 31696 56917 31702 56969
rect 31754 56957 31760 56969
rect 32083 56960 32141 56966
rect 32083 56957 32095 56960
rect 31754 56929 32095 56957
rect 31754 56917 31760 56929
rect 32083 56926 32095 56929
rect 32129 56926 32141 56960
rect 32083 56920 32141 56926
rect 33328 56917 33334 56969
rect 33386 56957 33392 56969
rect 34291 56960 34349 56966
rect 34291 56957 34303 56960
rect 33386 56929 34303 56957
rect 33386 56917 33392 56929
rect 34291 56926 34303 56929
rect 34337 56926 34349 56960
rect 34291 56920 34349 56926
rect 34864 56917 34870 56969
rect 34922 56957 34928 56969
rect 35251 56960 35309 56966
rect 35251 56957 35263 56960
rect 34922 56929 35263 56957
rect 34922 56917 34928 56929
rect 35251 56926 35263 56929
rect 35297 56926 35309 56960
rect 35251 56920 35309 56926
rect 36496 56917 36502 56969
rect 36554 56957 36560 56969
rect 36595 56960 36653 56966
rect 36595 56957 36607 56960
rect 36554 56929 36607 56957
rect 36554 56917 36560 56929
rect 36595 56926 36607 56929
rect 36641 56926 36653 56960
rect 36595 56920 36653 56926
rect 41200 56917 41206 56969
rect 41258 56957 41264 56969
rect 41971 56960 42029 56966
rect 41971 56957 41983 56960
rect 41258 56929 41983 56957
rect 41258 56917 41264 56929
rect 41971 56926 41983 56929
rect 42017 56926 42029 56960
rect 41971 56920 42029 56926
rect 47536 56917 47542 56969
rect 47594 56957 47600 56969
rect 47594 56929 47639 56957
rect 47594 56917 47600 56929
rect 52240 56917 52246 56969
rect 52298 56957 52304 56969
rect 52723 56960 52781 56966
rect 52723 56957 52735 56960
rect 52298 56929 52735 56957
rect 52298 56917 52304 56929
rect 52723 56926 52735 56929
rect 52769 56926 52781 56960
rect 52723 56920 52781 56926
rect 1744 56883 1750 56895
rect 1705 56855 1750 56883
rect 1744 56843 1750 56855
rect 1802 56843 1808 56895
rect 2608 56883 2614 56895
rect 2569 56855 2614 56883
rect 2608 56843 2614 56855
rect 2666 56843 2672 56895
rect 5107 56886 5165 56892
rect 5107 56852 5119 56886
rect 5153 56883 5165 56886
rect 7219 56886 7277 56892
rect 5153 56855 6494 56883
rect 5153 56852 5165 56855
rect 5107 56846 5165 56852
rect 6466 56821 6494 56855
rect 7219 56852 7231 56886
rect 7265 56883 7277 56886
rect 8272 56883 8278 56895
rect 7265 56855 8278 56883
rect 7265 56852 7277 56855
rect 7219 56846 7277 56852
rect 8272 56843 8278 56855
rect 8330 56843 8336 56895
rect 11248 56883 11254 56895
rect 11209 56855 11254 56883
rect 11248 56843 11254 56855
rect 11306 56843 11312 56895
rect 12208 56843 12214 56895
rect 12266 56883 12272 56895
rect 12979 56886 13037 56892
rect 12979 56883 12991 56886
rect 12266 56855 12991 56883
rect 12266 56843 12272 56855
rect 12979 56852 12991 56855
rect 13025 56852 13037 56886
rect 12979 56846 13037 56852
rect 13747 56886 13805 56892
rect 13747 56852 13759 56886
rect 13793 56883 13805 56886
rect 14032 56883 14038 56895
rect 13793 56855 14038 56883
rect 13793 56852 13805 56855
rect 13747 56846 13805 56852
rect 14032 56843 14038 56855
rect 14090 56843 14096 56895
rect 16144 56883 16150 56895
rect 16105 56855 16150 56883
rect 16144 56843 16150 56855
rect 16202 56843 16208 56895
rect 19315 56886 19373 56892
rect 19315 56883 19327 56886
rect 17266 56855 19327 56883
rect 6448 56769 6454 56821
rect 6506 56769 6512 56821
rect 12400 56769 12406 56821
rect 12458 56809 12464 56821
rect 17266 56809 17294 56855
rect 19315 56852 19327 56855
rect 19361 56852 19373 56886
rect 19315 56846 19373 56852
rect 21331 56886 21389 56892
rect 21331 56852 21343 56886
rect 21377 56883 21389 56886
rect 21616 56883 21622 56895
rect 21377 56855 21622 56883
rect 21377 56852 21389 56855
rect 21331 56846 21389 56852
rect 21616 56843 21622 56855
rect 21674 56843 21680 56895
rect 23344 56883 23350 56895
rect 23305 56855 23350 56883
rect 23344 56843 23350 56855
rect 23402 56843 23408 56895
rect 26035 56886 26093 56892
rect 26035 56852 26047 56886
rect 26081 56883 26093 56886
rect 26320 56883 26326 56895
rect 26081 56855 26326 56883
rect 26081 56852 26093 56855
rect 26035 56846 26093 56852
rect 26320 56843 26326 56855
rect 26378 56843 26384 56895
rect 28816 56883 28822 56895
rect 28777 56855 28822 56883
rect 28816 56843 28822 56855
rect 28874 56843 28880 56895
rect 31888 56883 31894 56895
rect 31849 56855 31894 56883
rect 31888 56843 31894 56855
rect 31946 56843 31952 56895
rect 32752 56883 32758 56895
rect 32713 56855 32758 56883
rect 32752 56843 32758 56855
rect 32810 56843 32816 56895
rect 34096 56883 34102 56895
rect 34057 56855 34102 56883
rect 34096 56843 34102 56855
rect 34154 56843 34160 56895
rect 35059 56886 35117 56892
rect 35059 56883 35071 56886
rect 34882 56855 35071 56883
rect 34882 56821 34910 56855
rect 35059 56852 35071 56855
rect 35105 56852 35117 56886
rect 35059 56846 35117 56852
rect 38032 56843 38038 56895
rect 38090 56883 38096 56895
rect 38227 56886 38285 56892
rect 38227 56883 38239 56886
rect 38090 56855 38239 56883
rect 38090 56843 38096 56855
rect 38227 56852 38239 56855
rect 38273 56852 38285 56886
rect 38227 56846 38285 56852
rect 39664 56843 39670 56895
rect 39722 56883 39728 56895
rect 40051 56886 40109 56892
rect 40051 56883 40063 56886
rect 39722 56855 40063 56883
rect 39722 56843 39728 56855
rect 40051 56852 40063 56855
rect 40097 56852 40109 56886
rect 40723 56886 40781 56892
rect 40723 56883 40735 56886
rect 40051 56846 40109 56852
rect 40450 56855 40735 56883
rect 12458 56781 17294 56809
rect 12458 56769 12464 56781
rect 34864 56769 34870 56821
rect 34922 56769 34928 56821
rect 40450 56747 40478 56855
rect 40723 56852 40735 56855
rect 40769 56883 40781 56886
rect 41011 56886 41069 56892
rect 41011 56883 41023 56886
rect 40769 56855 41023 56883
rect 40769 56852 40781 56855
rect 40723 56846 40781 56852
rect 41011 56852 41023 56855
rect 41057 56852 41069 56886
rect 41011 56846 41069 56852
rect 42832 56843 42838 56895
rect 42890 56883 42896 56895
rect 43219 56886 43277 56892
rect 43219 56883 43231 56886
rect 42890 56855 43231 56883
rect 42890 56843 42896 56855
rect 43219 56852 43231 56855
rect 43265 56852 43277 56886
rect 43219 56846 43277 56852
rect 44368 56843 44374 56895
rect 44426 56883 44432 56895
rect 45043 56886 45101 56892
rect 45043 56883 45055 56886
rect 44426 56855 45055 56883
rect 44426 56843 44432 56855
rect 45043 56852 45055 56855
rect 45089 56852 45101 56886
rect 45043 56846 45101 56852
rect 45904 56843 45910 56895
rect 45962 56883 45968 56895
rect 46291 56886 46349 56892
rect 46291 56883 46303 56886
rect 45962 56855 46303 56883
rect 45962 56843 45968 56855
rect 46291 56852 46303 56855
rect 46337 56852 46349 56886
rect 46291 56846 46349 56852
rect 48979 56886 49037 56892
rect 48979 56852 48991 56886
rect 49025 56883 49037 56886
rect 49072 56883 49078 56895
rect 49025 56855 49078 56883
rect 49025 56852 49037 56855
rect 48979 56846 49037 56852
rect 49072 56843 49078 56855
rect 49130 56843 49136 56895
rect 50704 56843 50710 56895
rect 50762 56883 50768 56895
rect 51091 56886 51149 56892
rect 51091 56883 51103 56886
rect 50762 56855 51103 56883
rect 50762 56843 50768 56855
rect 51091 56852 51103 56855
rect 51137 56852 51149 56886
rect 51091 56846 51149 56852
rect 53872 56843 53878 56895
rect 53930 56883 53936 56895
rect 54259 56886 54317 56892
rect 54259 56883 54271 56886
rect 53930 56855 54271 56883
rect 53930 56843 53936 56855
rect 54259 56852 54271 56855
rect 54305 56852 54317 56886
rect 54259 56846 54317 56852
rect 55408 56843 55414 56895
rect 55466 56883 55472 56895
rect 55795 56886 55853 56892
rect 55795 56883 55807 56886
rect 55466 56855 55807 56883
rect 55466 56843 55472 56855
rect 55795 56852 55807 56855
rect 55841 56852 55853 56886
rect 55795 56846 55853 56852
rect 57043 56886 57101 56892
rect 57043 56852 57055 56886
rect 57089 56883 57101 56886
rect 58576 56883 58582 56895
rect 57089 56855 58582 56883
rect 57089 56852 57101 56855
rect 57043 56846 57101 56852
rect 58576 56843 58582 56855
rect 58634 56843 58640 56895
rect 9808 56735 9814 56747
rect 9769 56707 9814 56735
rect 9808 56695 9814 56707
rect 9866 56695 9872 56747
rect 37936 56735 37942 56747
rect 37897 56707 37942 56735
rect 37936 56695 37942 56707
rect 37994 56695 38000 56747
rect 39760 56735 39766 56747
rect 39721 56707 39766 56735
rect 39760 56695 39766 56707
rect 39818 56695 39824 56747
rect 40432 56735 40438 56747
rect 40393 56707 40438 56735
rect 40432 56695 40438 56707
rect 40490 56695 40496 56747
rect 40816 56735 40822 56747
rect 40777 56707 40822 56735
rect 40816 56695 40822 56707
rect 40874 56695 40880 56747
rect 42928 56735 42934 56747
rect 42889 56707 42934 56735
rect 42928 56695 42934 56707
rect 42986 56695 42992 56747
rect 44752 56735 44758 56747
rect 44713 56707 44758 56735
rect 44752 56695 44758 56707
rect 44810 56695 44816 56747
rect 46003 56738 46061 56744
rect 46003 56704 46015 56738
rect 46049 56735 46061 56738
rect 46096 56735 46102 56747
rect 46049 56707 46102 56735
rect 46049 56704 46061 56707
rect 46003 56698 46061 56704
rect 46096 56695 46102 56707
rect 46154 56695 46160 56747
rect 48688 56735 48694 56747
rect 48649 56707 48694 56735
rect 48688 56695 48694 56707
rect 48746 56695 48752 56747
rect 50800 56735 50806 56747
rect 50761 56707 50806 56735
rect 50800 56695 50806 56707
rect 50858 56695 50864 56747
rect 53872 56695 53878 56747
rect 53930 56735 53936 56747
rect 53971 56738 54029 56744
rect 53971 56735 53983 56738
rect 53930 56707 53983 56735
rect 53930 56695 53936 56707
rect 53971 56704 53983 56707
rect 54017 56704 54029 56738
rect 55504 56735 55510 56747
rect 55465 56707 55510 56735
rect 53971 56698 54029 56704
rect 55504 56695 55510 56707
rect 55562 56695 55568 56747
rect 56752 56735 56758 56747
rect 56713 56707 56758 56735
rect 56752 56695 56758 56707
rect 56810 56695 56816 56747
rect 1152 56636 58848 56658
rect 1152 56584 19654 56636
rect 19706 56584 19718 56636
rect 19770 56584 19782 56636
rect 19834 56584 19846 56636
rect 19898 56584 50374 56636
rect 50426 56584 50438 56636
rect 50490 56584 50502 56636
rect 50554 56584 50566 56636
rect 50618 56584 58848 56636
rect 1152 56562 58848 56584
rect 688 56473 694 56525
rect 746 56513 752 56525
rect 1651 56516 1709 56522
rect 1651 56513 1663 56516
rect 746 56485 1663 56513
rect 746 56473 752 56485
rect 1651 56482 1663 56485
rect 1697 56482 1709 56516
rect 1651 56476 1709 56482
rect 2224 56473 2230 56525
rect 2282 56513 2288 56525
rect 2419 56516 2477 56522
rect 2419 56513 2431 56516
rect 2282 56485 2431 56513
rect 2282 56473 2288 56485
rect 2419 56482 2431 56485
rect 2465 56482 2477 56516
rect 2419 56476 2477 56482
rect 2800 56473 2806 56525
rect 2858 56513 2864 56525
rect 3187 56516 3245 56522
rect 3187 56513 3199 56516
rect 2858 56485 3199 56513
rect 2858 56473 2864 56485
rect 3187 56482 3199 56485
rect 3233 56482 3245 56516
rect 3187 56476 3245 56482
rect 3856 56473 3862 56525
rect 3914 56513 3920 56525
rect 4435 56516 4493 56522
rect 4435 56513 4447 56516
rect 3914 56485 4447 56513
rect 3914 56473 3920 56485
rect 4435 56482 4447 56485
rect 4481 56482 4493 56516
rect 4435 56476 4493 56482
rect 5392 56473 5398 56525
rect 5450 56513 5456 56525
rect 5491 56516 5549 56522
rect 5491 56513 5503 56516
rect 5450 56485 5503 56513
rect 5450 56473 5456 56485
rect 5491 56482 5503 56485
rect 5537 56482 5549 56516
rect 5491 56476 5549 56482
rect 5968 56473 5974 56525
rect 6026 56513 6032 56525
rect 6259 56516 6317 56522
rect 6259 56513 6271 56516
rect 6026 56485 6271 56513
rect 6026 56473 6032 56485
rect 6259 56482 6271 56485
rect 6305 56482 6317 56516
rect 6259 56476 6317 56482
rect 7024 56473 7030 56525
rect 7082 56513 7088 56525
rect 7123 56516 7181 56522
rect 7123 56513 7135 56516
rect 7082 56485 7135 56513
rect 7082 56473 7088 56485
rect 7123 56482 7135 56485
rect 7169 56482 7181 56516
rect 7123 56476 7181 56482
rect 8467 56516 8525 56522
rect 8467 56482 8479 56516
rect 8513 56513 8525 56516
rect 8560 56513 8566 56525
rect 8513 56485 8566 56513
rect 8513 56482 8525 56485
rect 8467 56476 8525 56482
rect 8560 56473 8566 56485
rect 8618 56473 8624 56525
rect 10192 56473 10198 56525
rect 10250 56513 10256 56525
rect 10291 56516 10349 56522
rect 10291 56513 10303 56516
rect 10250 56485 10303 56513
rect 10250 56473 10256 56485
rect 10291 56482 10303 56485
rect 10337 56482 10349 56516
rect 10291 56476 10349 56482
rect 10672 56473 10678 56525
rect 10730 56513 10736 56525
rect 11059 56516 11117 56522
rect 11059 56513 11071 56516
rect 10730 56485 11071 56513
rect 10730 56473 10736 56485
rect 11059 56482 11071 56485
rect 11105 56482 11117 56516
rect 11059 56476 11117 56482
rect 11728 56473 11734 56525
rect 11786 56513 11792 56525
rect 11827 56516 11885 56522
rect 11827 56513 11839 56516
rect 11786 56485 11839 56513
rect 11786 56473 11792 56485
rect 11827 56482 11839 56485
rect 11873 56482 11885 56516
rect 11827 56476 11885 56482
rect 12304 56473 12310 56525
rect 12362 56513 12368 56525
rect 12595 56516 12653 56522
rect 12595 56513 12607 56516
rect 12362 56485 12607 56513
rect 12362 56473 12368 56485
rect 12595 56482 12607 56485
rect 12641 56482 12653 56516
rect 12595 56476 12653 56482
rect 13360 56473 13366 56525
rect 13418 56513 13424 56525
rect 13459 56516 13517 56522
rect 13459 56513 13471 56516
rect 13418 56485 13471 56513
rect 13418 56473 13424 56485
rect 13459 56482 13471 56485
rect 13505 56482 13517 56516
rect 13459 56476 13517 56482
rect 14896 56473 14902 56525
rect 14954 56513 14960 56525
rect 14995 56516 15053 56522
rect 14995 56513 15007 56516
rect 14954 56485 15007 56513
rect 14954 56473 14960 56485
rect 14995 56482 15007 56485
rect 15041 56482 15053 56516
rect 14995 56476 15053 56482
rect 17008 56473 17014 56525
rect 17066 56513 17072 56525
rect 17107 56516 17165 56522
rect 17107 56513 17119 56516
rect 17066 56485 17119 56513
rect 17066 56473 17072 56485
rect 17107 56482 17119 56485
rect 17153 56482 17165 56516
rect 18736 56513 18742 56525
rect 18697 56485 18742 56513
rect 17107 56476 17165 56482
rect 18736 56473 18742 56485
rect 18794 56473 18800 56525
rect 19984 56473 19990 56525
rect 20042 56513 20048 56525
rect 20275 56516 20333 56522
rect 20275 56513 20287 56516
rect 20042 56485 20287 56513
rect 20042 56473 20048 56485
rect 20275 56482 20287 56485
rect 20321 56482 20333 56516
rect 20275 56476 20333 56482
rect 21232 56473 21238 56525
rect 21290 56513 21296 56525
rect 21331 56516 21389 56522
rect 21331 56513 21343 56516
rect 21290 56485 21343 56513
rect 21290 56473 21296 56485
rect 21331 56482 21343 56485
rect 21377 56482 21389 56516
rect 21331 56476 21389 56482
rect 21712 56473 21718 56525
rect 21770 56513 21776 56525
rect 22195 56516 22253 56522
rect 22195 56513 22207 56516
rect 21770 56485 22207 56513
rect 21770 56473 21776 56485
rect 22195 56482 22207 56485
rect 22241 56482 22253 56516
rect 22195 56476 22253 56482
rect 22768 56473 22774 56525
rect 22826 56513 22832 56525
rect 22867 56516 22925 56522
rect 22867 56513 22879 56516
rect 22826 56485 22879 56513
rect 22826 56473 22832 56485
rect 22867 56482 22879 56485
rect 22913 56482 22925 56516
rect 22867 56476 22925 56482
rect 24307 56516 24365 56522
rect 24307 56482 24319 56516
rect 24353 56513 24365 56516
rect 24400 56513 24406 56525
rect 24353 56485 24406 56513
rect 24353 56482 24365 56485
rect 24307 56476 24365 56482
rect 24400 56473 24406 56485
rect 24458 56473 24464 56525
rect 25936 56473 25942 56525
rect 25994 56513 26000 56525
rect 26035 56516 26093 56522
rect 26035 56513 26047 56516
rect 25994 56485 26047 56513
rect 25994 56473 26000 56485
rect 26035 56482 26047 56485
rect 26081 56482 26093 56516
rect 26035 56476 26093 56482
rect 26512 56473 26518 56525
rect 26570 56513 26576 56525
rect 26803 56516 26861 56522
rect 26803 56513 26815 56516
rect 26570 56485 26815 56513
rect 26570 56473 26576 56485
rect 26803 56482 26815 56485
rect 26849 56482 26861 56516
rect 26803 56476 26861 56482
rect 27568 56473 27574 56525
rect 27626 56513 27632 56525
rect 27667 56516 27725 56522
rect 27667 56513 27679 56516
rect 27626 56485 27679 56513
rect 27626 56473 27632 56485
rect 27667 56482 27679 56485
rect 27713 56482 27725 56516
rect 27667 56476 27725 56482
rect 28048 56473 28054 56525
rect 28106 56513 28112 56525
rect 28531 56516 28589 56522
rect 28531 56513 28543 56516
rect 28106 56485 28543 56513
rect 28106 56473 28112 56485
rect 28531 56482 28543 56485
rect 28577 56482 28589 56516
rect 29680 56513 29686 56525
rect 29641 56485 29686 56513
rect 28531 56476 28589 56482
rect 29680 56473 29686 56485
rect 29738 56473 29744 56525
rect 30640 56473 30646 56525
rect 30698 56513 30704 56525
rect 30835 56516 30893 56522
rect 30835 56513 30847 56516
rect 30698 56485 30847 56513
rect 30698 56473 30704 56485
rect 30835 56482 30847 56485
rect 30881 56482 30893 56516
rect 30835 56476 30893 56482
rect 32272 56473 32278 56525
rect 32330 56513 32336 56525
rect 32371 56516 32429 56522
rect 32371 56513 32383 56516
rect 32330 56485 32383 56513
rect 32330 56473 32336 56485
rect 32371 56482 32383 56485
rect 32417 56482 32429 56516
rect 32371 56476 32429 56482
rect 32848 56473 32854 56525
rect 32906 56513 32912 56525
rect 33139 56516 33197 56522
rect 33139 56513 33151 56516
rect 32906 56485 33151 56513
rect 32906 56473 32912 56485
rect 33139 56482 33151 56485
rect 33185 56482 33197 56516
rect 33139 56476 33197 56482
rect 33808 56473 33814 56525
rect 33866 56513 33872 56525
rect 33907 56516 33965 56522
rect 33907 56513 33919 56516
rect 33866 56485 33919 56513
rect 33866 56473 33872 56485
rect 33907 56482 33919 56485
rect 33953 56482 33965 56516
rect 33907 56476 33965 56482
rect 34384 56473 34390 56525
rect 34442 56513 34448 56525
rect 34675 56516 34733 56522
rect 34675 56513 34687 56516
rect 34442 56485 34687 56513
rect 34442 56473 34448 56485
rect 34675 56482 34687 56485
rect 34721 56482 34733 56516
rect 34675 56476 34733 56482
rect 35440 56473 35446 56525
rect 35498 56513 35504 56525
rect 36115 56516 36173 56522
rect 36115 56513 36127 56516
rect 35498 56485 36127 56513
rect 35498 56473 35504 56485
rect 36115 56482 36127 56485
rect 36161 56482 36173 56516
rect 36115 56476 36173 56482
rect 36979 56516 37037 56522
rect 36979 56482 36991 56516
rect 37025 56482 37037 56516
rect 36979 56476 37037 56482
rect 36016 56399 36022 56451
rect 36074 56439 36080 56451
rect 36994 56439 37022 56476
rect 37552 56473 37558 56525
rect 37610 56513 37616 56525
rect 37747 56516 37805 56522
rect 37747 56513 37759 56516
rect 37610 56485 37759 56513
rect 37610 56473 37616 56485
rect 37747 56482 37759 56485
rect 37793 56482 37805 56516
rect 37747 56476 37805 56482
rect 38608 56473 38614 56525
rect 38666 56513 38672 56525
rect 38803 56516 38861 56522
rect 38803 56513 38815 56516
rect 38666 56485 38815 56513
rect 38666 56473 38672 56485
rect 38803 56482 38815 56485
rect 38849 56482 38861 56516
rect 38803 56476 38861 56482
rect 40144 56473 40150 56525
rect 40202 56513 40208 56525
rect 40243 56516 40301 56522
rect 40243 56513 40255 56516
rect 40202 56485 40255 56513
rect 40202 56473 40208 56485
rect 40243 56482 40255 56485
rect 40289 56482 40301 56516
rect 40243 56476 40301 56482
rect 41776 56473 41782 56525
rect 41834 56513 41840 56525
rect 41875 56516 41933 56522
rect 41875 56513 41887 56516
rect 41834 56485 41887 56513
rect 41834 56473 41840 56485
rect 41875 56482 41887 56485
rect 41921 56482 41933 56516
rect 41875 56476 41933 56482
rect 42256 56473 42262 56525
rect 42314 56513 42320 56525
rect 42739 56516 42797 56522
rect 42739 56513 42751 56516
rect 42314 56485 42751 56513
rect 42314 56473 42320 56485
rect 42739 56482 42751 56485
rect 42785 56482 42797 56516
rect 42739 56476 42797 56482
rect 43312 56473 43318 56525
rect 43370 56513 43376 56525
rect 43411 56516 43469 56522
rect 43411 56513 43423 56516
rect 43370 56485 43423 56513
rect 43370 56473 43376 56485
rect 43411 56482 43423 56485
rect 43457 56482 43469 56516
rect 43411 56476 43469 56482
rect 43888 56473 43894 56525
rect 43946 56513 43952 56525
rect 44275 56516 44333 56522
rect 44275 56513 44287 56516
rect 43946 56485 44287 56513
rect 43946 56473 43952 56485
rect 44275 56482 44287 56485
rect 44321 56482 44333 56516
rect 44275 56476 44333 56482
rect 44944 56473 44950 56525
rect 45002 56513 45008 56525
rect 45043 56516 45101 56522
rect 45043 56513 45055 56516
rect 45002 56485 45055 56513
rect 45002 56473 45008 56485
rect 45043 56482 45055 56485
rect 45089 56482 45101 56516
rect 45043 56476 45101 56482
rect 46480 56473 46486 56525
rect 46538 56513 46544 56525
rect 46771 56516 46829 56522
rect 46771 56513 46783 56516
rect 46538 56485 46783 56513
rect 46538 56473 46544 56485
rect 46771 56482 46783 56485
rect 46817 56482 46829 56516
rect 46771 56476 46829 56482
rect 48016 56473 48022 56525
rect 48074 56513 48080 56525
rect 48115 56516 48173 56522
rect 48115 56513 48127 56516
rect 48074 56485 48127 56513
rect 48074 56473 48080 56485
rect 48115 56482 48127 56485
rect 48161 56482 48173 56516
rect 48115 56476 48173 56482
rect 48592 56473 48598 56525
rect 48650 56513 48656 56525
rect 48979 56516 49037 56522
rect 48979 56513 48991 56516
rect 48650 56485 48991 56513
rect 48650 56473 48656 56485
rect 48979 56482 48991 56485
rect 49025 56482 49037 56516
rect 48979 56476 49037 56482
rect 49648 56473 49654 56525
rect 49706 56513 49712 56525
rect 49747 56516 49805 56522
rect 49747 56513 49759 56516
rect 49706 56485 49759 56513
rect 49706 56473 49712 56485
rect 49747 56482 49759 56485
rect 49793 56482 49805 56516
rect 49747 56476 49805 56482
rect 50128 56473 50134 56525
rect 50186 56513 50192 56525
rect 50611 56516 50669 56522
rect 50611 56513 50623 56516
rect 50186 56485 50623 56513
rect 50186 56473 50192 56485
rect 50611 56482 50623 56485
rect 50657 56482 50669 56516
rect 50611 56476 50669 56482
rect 52816 56473 52822 56525
rect 52874 56513 52880 56525
rect 53011 56516 53069 56522
rect 53011 56513 53023 56516
rect 52874 56485 53023 56513
rect 52874 56473 52880 56485
rect 53011 56482 53023 56485
rect 53057 56482 53069 56516
rect 53011 56476 53069 56482
rect 53296 56473 53302 56525
rect 53354 56513 53360 56525
rect 53779 56516 53837 56522
rect 53779 56513 53791 56516
rect 53354 56485 53791 56513
rect 53354 56473 53360 56485
rect 53779 56482 53791 56485
rect 53825 56482 53837 56516
rect 53779 56476 53837 56482
rect 54352 56473 54358 56525
rect 54410 56513 54416 56525
rect 54451 56516 54509 56522
rect 54451 56513 54463 56516
rect 54410 56485 54463 56513
rect 54410 56473 54416 56485
rect 54451 56482 54463 56485
rect 54497 56482 54509 56516
rect 54451 56476 54509 56482
rect 54928 56473 54934 56525
rect 54986 56513 54992 56525
rect 55315 56516 55373 56522
rect 55315 56513 55327 56516
rect 54986 56485 55327 56513
rect 54986 56473 54992 56485
rect 55315 56482 55327 56485
rect 55361 56482 55373 56516
rect 55984 56513 55990 56525
rect 55945 56485 55990 56513
rect 55315 56476 55373 56482
rect 55984 56473 55990 56485
rect 56042 56473 56048 56525
rect 36074 56411 37022 56439
rect 36074 56399 36080 56411
rect 39568 56399 39574 56451
rect 39626 56439 39632 56451
rect 56752 56439 56758 56451
rect 39626 56411 56758 56439
rect 39626 56399 39632 56411
rect 56752 56399 56758 56411
rect 56810 56399 56816 56451
rect 33235 56368 33293 56374
rect 33235 56334 33247 56368
rect 33281 56365 33293 56368
rect 42352 56365 42358 56377
rect 33281 56337 42358 56365
rect 33281 56334 33293 56337
rect 33235 56328 33293 56334
rect 42352 56325 42358 56337
rect 42410 56325 42416 56377
rect 47056 56325 47062 56377
rect 47114 56365 47120 56377
rect 56083 56368 56141 56374
rect 56083 56365 56095 56368
rect 47114 56337 56095 56365
rect 47114 56325 47120 56337
rect 56083 56334 56095 56337
rect 56129 56334 56141 56368
rect 56083 56328 56141 56334
rect 7219 56294 7277 56300
rect 7219 56260 7231 56294
rect 7265 56291 7277 56294
rect 12496 56291 12502 56303
rect 7265 56263 12502 56291
rect 7265 56260 7277 56263
rect 7219 56254 7277 56260
rect 12496 56251 12502 56263
rect 12554 56251 12560 56303
rect 13744 56251 13750 56303
rect 13802 56291 13808 56303
rect 15475 56294 15533 56300
rect 15475 56291 15487 56294
rect 13802 56263 15487 56291
rect 13802 56251 13808 56263
rect 15475 56260 15487 56263
rect 15521 56291 15533 56294
rect 15763 56294 15821 56300
rect 15763 56291 15775 56294
rect 15521 56263 15775 56291
rect 15521 56260 15533 56263
rect 15475 56254 15533 56260
rect 15763 56260 15775 56263
rect 15809 56260 15821 56294
rect 15763 56254 15821 56260
rect 43888 56251 43894 56303
rect 43946 56291 43952 56303
rect 45139 56294 45197 56300
rect 45139 56291 45151 56294
rect 43946 56263 45151 56291
rect 43946 56251 43952 56263
rect 45139 56260 45151 56263
rect 45185 56260 45197 56294
rect 45139 56254 45197 56260
rect 46864 56251 46870 56303
rect 46922 56291 46928 56303
rect 49843 56294 49901 56300
rect 49843 56291 49855 56294
rect 46922 56263 49855 56291
rect 46922 56251 46928 56263
rect 49843 56260 49855 56263
rect 49889 56260 49901 56294
rect 52243 56294 52301 56300
rect 52243 56291 52255 56294
rect 49843 56254 49901 56260
rect 51970 56263 52255 56291
rect 1747 56220 1805 56226
rect 1747 56186 1759 56220
rect 1793 56217 1805 56220
rect 1840 56217 1846 56229
rect 1793 56189 1846 56217
rect 1793 56186 1805 56189
rect 1747 56180 1805 56186
rect 1840 56177 1846 56189
rect 1898 56177 1904 56229
rect 2227 56220 2285 56226
rect 2227 56186 2239 56220
rect 2273 56217 2285 56220
rect 2515 56220 2573 56226
rect 2515 56217 2527 56220
rect 2273 56189 2527 56217
rect 2273 56186 2285 56189
rect 2227 56180 2285 56186
rect 2515 56186 2527 56189
rect 2561 56217 2573 56220
rect 2704 56217 2710 56229
rect 2561 56189 2710 56217
rect 2561 56186 2573 56189
rect 2515 56180 2573 56186
rect 2704 56177 2710 56189
rect 2762 56177 2768 56229
rect 2992 56217 2998 56229
rect 2953 56189 2998 56217
rect 2992 56177 2998 56189
rect 3050 56217 3056 56229
rect 3283 56220 3341 56226
rect 3283 56217 3295 56220
rect 3050 56189 3295 56217
rect 3050 56177 3056 56189
rect 3283 56186 3295 56189
rect 3329 56186 3341 56220
rect 3283 56180 3341 56186
rect 4531 56220 4589 56226
rect 4531 56186 4543 56220
rect 4577 56217 4589 56220
rect 5008 56217 5014 56229
rect 4577 56189 5014 56217
rect 4577 56186 4589 56189
rect 4531 56180 4589 56186
rect 5008 56177 5014 56189
rect 5066 56177 5072 56229
rect 5200 56217 5206 56229
rect 5161 56189 5206 56217
rect 5200 56177 5206 56189
rect 5258 56217 5264 56229
rect 5587 56220 5645 56226
rect 5587 56217 5599 56220
rect 5258 56189 5599 56217
rect 5258 56177 5264 56189
rect 5587 56186 5599 56189
rect 5633 56186 5645 56220
rect 5587 56180 5645 56186
rect 6067 56220 6125 56226
rect 6067 56186 6079 56220
rect 6113 56217 6125 56220
rect 6352 56217 6358 56229
rect 6113 56189 6358 56217
rect 6113 56186 6125 56189
rect 6067 56180 6125 56186
rect 6352 56177 6358 56189
rect 6410 56177 6416 56229
rect 8275 56220 8333 56226
rect 8275 56186 8287 56220
rect 8321 56217 8333 56220
rect 8560 56217 8566 56229
rect 8321 56189 8566 56217
rect 8321 56186 8333 56189
rect 8275 56180 8333 56186
rect 8560 56177 8566 56189
rect 8618 56177 8624 56229
rect 10384 56217 10390 56229
rect 10345 56189 10390 56217
rect 10384 56177 10390 56189
rect 10442 56177 10448 56229
rect 10768 56217 10774 56229
rect 10729 56189 10774 56217
rect 10768 56177 10774 56189
rect 10826 56217 10832 56229
rect 11155 56220 11213 56226
rect 11155 56217 11167 56220
rect 10826 56189 11167 56217
rect 10826 56177 10832 56189
rect 11155 56186 11167 56189
rect 11201 56186 11213 56220
rect 11920 56217 11926 56229
rect 11881 56189 11926 56217
rect 11155 56180 11213 56186
rect 11920 56177 11926 56189
rect 11978 56177 11984 56229
rect 12688 56217 12694 56229
rect 12649 56189 12694 56217
rect 12688 56177 12694 56189
rect 12746 56177 12752 56229
rect 13267 56220 13325 56226
rect 13267 56186 13279 56220
rect 13313 56217 13325 56220
rect 13552 56217 13558 56229
rect 13313 56189 13558 56217
rect 13313 56186 13325 56189
rect 13267 56180 13325 56186
rect 13552 56177 13558 56189
rect 13610 56177 13616 56229
rect 15091 56220 15149 56226
rect 15091 56186 15103 56220
rect 15137 56217 15149 56220
rect 15184 56217 15190 56229
rect 15137 56189 15190 56217
rect 15137 56186 15149 56189
rect 15091 56180 15149 56186
rect 15184 56177 15190 56189
rect 15242 56177 15248 56229
rect 15859 56220 15917 56226
rect 15859 56186 15871 56220
rect 15905 56186 15917 56220
rect 16816 56217 16822 56229
rect 16777 56189 16822 56217
rect 15859 56180 15917 56186
rect 15376 56103 15382 56155
rect 15434 56143 15440 56155
rect 15874 56143 15902 56180
rect 16816 56177 16822 56189
rect 16874 56217 16880 56229
rect 17203 56220 17261 56226
rect 17203 56217 17215 56220
rect 16874 56189 17215 56217
rect 16874 56177 16880 56189
rect 17203 56186 17215 56189
rect 17249 56186 17261 56220
rect 17203 56180 17261 56186
rect 18451 56220 18509 56226
rect 18451 56186 18463 56220
rect 18497 56217 18509 56220
rect 18640 56217 18646 56229
rect 18497 56189 18646 56217
rect 18497 56186 18509 56189
rect 18451 56180 18509 56186
rect 18640 56177 18646 56189
rect 18698 56177 18704 56229
rect 20083 56220 20141 56226
rect 20083 56186 20095 56220
rect 20129 56217 20141 56220
rect 20371 56220 20429 56226
rect 20371 56217 20383 56220
rect 20129 56189 20383 56217
rect 20129 56186 20141 56189
rect 20083 56180 20141 56186
rect 20371 56186 20383 56189
rect 20417 56217 20429 56220
rect 20848 56217 20854 56229
rect 20417 56189 20854 56217
rect 20417 56186 20429 56189
rect 20371 56180 20429 56186
rect 20848 56177 20854 56189
rect 20906 56177 20912 56229
rect 21139 56220 21197 56226
rect 21139 56186 21151 56220
rect 21185 56217 21197 56220
rect 21424 56217 21430 56229
rect 21185 56189 21430 56217
rect 21185 56186 21197 56189
rect 21139 56180 21197 56186
rect 21424 56177 21430 56189
rect 21482 56177 21488 56229
rect 21907 56220 21965 56226
rect 21907 56186 21919 56220
rect 21953 56217 21965 56220
rect 22096 56217 22102 56229
rect 21953 56189 22102 56217
rect 21953 56186 21965 56189
rect 21907 56180 21965 56186
rect 22096 56177 22102 56189
rect 22154 56177 22160 56229
rect 22960 56177 22966 56229
rect 23018 56217 23024 56229
rect 24400 56217 24406 56229
rect 23018 56189 23063 56217
rect 24361 56189 24406 56217
rect 23018 56177 23024 56189
rect 24400 56177 24406 56189
rect 24458 56177 24464 56229
rect 26128 56217 26134 56229
rect 26089 56189 26134 56217
rect 26128 56177 26134 56189
rect 26186 56177 26192 56229
rect 26896 56217 26902 56229
rect 26857 56189 26902 56217
rect 26896 56177 26902 56189
rect 26954 56177 26960 56229
rect 27475 56220 27533 56226
rect 27475 56186 27487 56220
rect 27521 56217 27533 56220
rect 27760 56217 27766 56229
rect 27521 56189 27766 56217
rect 27521 56186 27533 56189
rect 27475 56180 27533 56186
rect 27760 56177 27766 56189
rect 27818 56177 27824 56229
rect 28144 56217 28150 56229
rect 28105 56189 28150 56217
rect 28144 56177 28150 56189
rect 28202 56217 28208 56229
rect 28435 56220 28493 56226
rect 28435 56217 28447 56220
rect 28202 56189 28447 56217
rect 28202 56177 28208 56189
rect 28435 56186 28447 56189
rect 28481 56186 28493 56220
rect 28435 56180 28493 56186
rect 29395 56220 29453 56226
rect 29395 56186 29407 56220
rect 29441 56217 29453 56220
rect 29584 56217 29590 56229
rect 29441 56189 29590 56217
rect 29441 56186 29453 56189
rect 29395 56180 29453 56186
rect 29584 56177 29590 56189
rect 29642 56177 29648 56229
rect 30928 56217 30934 56229
rect 30889 56189 30934 56217
rect 30928 56177 30934 56189
rect 30986 56177 30992 56229
rect 31312 56217 31318 56229
rect 31273 56189 31318 56217
rect 31312 56177 31318 56189
rect 31370 56217 31376 56229
rect 31603 56220 31661 56226
rect 31603 56217 31615 56220
rect 31370 56189 31615 56217
rect 31370 56177 31376 56189
rect 31603 56186 31615 56189
rect 31649 56186 31661 56220
rect 31603 56180 31661 56186
rect 31699 56220 31757 56226
rect 31699 56186 31711 56220
rect 31745 56186 31757 56220
rect 32464 56217 32470 56229
rect 32425 56189 32470 56217
rect 31699 56180 31757 56186
rect 15434 56115 15902 56143
rect 15434 56103 15440 56115
rect 31216 56103 31222 56155
rect 31274 56143 31280 56155
rect 31714 56143 31742 56180
rect 32464 56177 32470 56189
rect 32522 56177 32528 56229
rect 34000 56217 34006 56229
rect 33961 56189 34006 56217
rect 34000 56177 34006 56189
rect 34058 56177 34064 56229
rect 34483 56220 34541 56226
rect 34483 56186 34495 56220
rect 34529 56217 34541 56220
rect 34768 56217 34774 56229
rect 34529 56189 34774 56217
rect 34529 56186 34541 56189
rect 34483 56180 34541 56186
rect 34768 56177 34774 56189
rect 34826 56177 34832 56229
rect 35344 56177 35350 56229
rect 35402 56217 35408 56229
rect 36211 56220 36269 56226
rect 36211 56217 36223 56220
rect 35402 56189 36223 56217
rect 35402 56177 35408 56189
rect 36211 56186 36223 56189
rect 36257 56186 36269 56220
rect 36211 56180 36269 56186
rect 36691 56220 36749 56226
rect 36691 56186 36703 56220
rect 36737 56217 36749 56220
rect 36880 56217 36886 56229
rect 36737 56189 36886 56217
rect 36737 56186 36749 56189
rect 36691 56180 36749 56186
rect 36880 56177 36886 56189
rect 36938 56177 36944 56229
rect 37456 56177 37462 56229
rect 37514 56217 37520 56229
rect 37651 56220 37709 56226
rect 37651 56217 37663 56220
rect 37514 56189 37663 56217
rect 37514 56177 37520 56189
rect 37651 56186 37663 56189
rect 37697 56217 37709 56220
rect 37939 56220 37997 56226
rect 37939 56217 37951 56220
rect 37697 56189 37951 56217
rect 37697 56186 37709 56189
rect 37651 56180 37709 56186
rect 37939 56186 37951 56189
rect 37985 56186 37997 56220
rect 38416 56217 38422 56229
rect 38377 56189 38422 56217
rect 37939 56180 37997 56186
rect 38416 56177 38422 56189
rect 38474 56217 38480 56229
rect 38707 56220 38765 56226
rect 38707 56217 38719 56220
rect 38474 56189 38719 56217
rect 38474 56177 38480 56189
rect 38707 56186 38719 56189
rect 38753 56186 38765 56220
rect 39856 56217 39862 56229
rect 39817 56189 39862 56217
rect 38707 56180 38765 56186
rect 39856 56177 39862 56189
rect 39914 56217 39920 56229
rect 40147 56220 40205 56226
rect 40147 56217 40159 56220
rect 39914 56189 40159 56217
rect 39914 56177 39920 56189
rect 40147 56186 40159 56189
rect 40193 56186 40205 56220
rect 40147 56180 40205 56186
rect 41683 56220 41741 56226
rect 41683 56186 41695 56220
rect 41729 56217 41741 56220
rect 41971 56220 42029 56226
rect 41971 56217 41983 56220
rect 41729 56189 41983 56217
rect 41729 56186 41741 56189
rect 41683 56180 41741 56186
rect 41971 56186 41983 56189
rect 42017 56217 42029 56220
rect 42064 56217 42070 56229
rect 42017 56189 42070 56217
rect 42017 56186 42029 56189
rect 41971 56180 42029 56186
rect 42064 56177 42070 56189
rect 42122 56177 42128 56229
rect 42451 56220 42509 56226
rect 42451 56186 42463 56220
rect 42497 56217 42509 56220
rect 42640 56217 42646 56229
rect 42497 56189 42646 56217
rect 42497 56186 42509 56189
rect 42451 56180 42509 56186
rect 42640 56177 42646 56189
rect 42698 56177 42704 56229
rect 43504 56217 43510 56229
rect 43465 56189 43510 56217
rect 43504 56177 43510 56189
rect 43562 56177 43568 56229
rect 43987 56220 44045 56226
rect 43987 56186 43999 56220
rect 44033 56217 44045 56220
rect 44176 56217 44182 56229
rect 44033 56189 44182 56217
rect 44033 56186 44045 56189
rect 43987 56180 44045 56186
rect 44176 56177 44182 56189
rect 44234 56217 44240 56229
rect 44467 56220 44525 56226
rect 44467 56217 44479 56220
rect 44234 56189 44479 56217
rect 44234 56177 44240 56189
rect 44467 56186 44479 56189
rect 44513 56186 44525 56220
rect 44467 56180 44525 56186
rect 46483 56220 46541 56226
rect 46483 56186 46495 56220
rect 46529 56217 46541 56220
rect 46672 56217 46678 56229
rect 46529 56189 46678 56217
rect 46529 56186 46541 56189
rect 46483 56180 46541 56186
rect 46672 56177 46678 56189
rect 46730 56177 46736 56229
rect 48208 56217 48214 56229
rect 48169 56189 48214 56217
rect 48208 56177 48214 56189
rect 48266 56177 48272 56229
rect 48592 56217 48598 56229
rect 48553 56189 48598 56217
rect 48592 56177 48598 56189
rect 48650 56217 48656 56229
rect 48883 56220 48941 56226
rect 48883 56217 48895 56220
rect 48650 56189 48895 56217
rect 48650 56177 48656 56189
rect 48883 56186 48895 56189
rect 48929 56186 48941 56220
rect 50224 56217 50230 56229
rect 50185 56189 50230 56217
rect 48883 56180 48941 56186
rect 50224 56177 50230 56189
rect 50282 56217 50288 56229
rect 50515 56220 50573 56226
rect 50515 56217 50527 56220
rect 50282 56189 50527 56217
rect 50282 56177 50288 56189
rect 50515 56186 50527 56189
rect 50561 56186 50573 56220
rect 50515 56180 50573 56186
rect 51280 56177 51286 56229
rect 51338 56217 51344 56229
rect 51970 56226 51998 56263
rect 52243 56260 52255 56263
rect 52289 56260 52301 56294
rect 52243 56254 52301 56260
rect 57040 56251 57046 56303
rect 57098 56291 57104 56303
rect 57139 56294 57197 56300
rect 57139 56291 57151 56294
rect 57098 56263 57151 56291
rect 57098 56251 57104 56263
rect 57139 56260 57151 56263
rect 57185 56260 57197 56294
rect 57139 56254 57197 56260
rect 51667 56220 51725 56226
rect 51667 56217 51679 56220
rect 51338 56189 51679 56217
rect 51338 56177 51344 56189
rect 51667 56186 51679 56189
rect 51713 56217 51725 56220
rect 51955 56220 52013 56226
rect 51955 56217 51967 56220
rect 51713 56189 51967 56217
rect 51713 56186 51725 56189
rect 51667 56180 51725 56186
rect 51955 56186 51967 56189
rect 52001 56186 52013 56220
rect 51955 56180 52013 56186
rect 52051 56220 52109 56226
rect 52051 56186 52063 56220
rect 52097 56186 52109 56220
rect 52051 56180 52109 56186
rect 52723 56220 52781 56226
rect 52723 56186 52735 56220
rect 52769 56217 52781 56220
rect 52912 56217 52918 56229
rect 52769 56189 52918 56217
rect 52769 56186 52781 56189
rect 52723 56180 52781 56186
rect 31274 56115 31742 56143
rect 31274 56103 31280 56115
rect 51184 56103 51190 56155
rect 51242 56143 51248 56155
rect 52066 56143 52094 56180
rect 52912 56177 52918 56189
rect 52970 56177 52976 56229
rect 53491 56220 53549 56226
rect 53491 56186 53503 56220
rect 53537 56217 53549 56220
rect 53683 56220 53741 56226
rect 53683 56217 53695 56220
rect 53537 56189 53695 56217
rect 53537 56186 53549 56189
rect 53491 56180 53549 56186
rect 53683 56186 53695 56189
rect 53729 56217 53741 56220
rect 53968 56217 53974 56229
rect 53729 56189 53974 56217
rect 53729 56186 53741 56189
rect 53683 56180 53741 56186
rect 53968 56177 53974 56189
rect 54026 56177 54032 56229
rect 54544 56217 54550 56229
rect 54505 56189 54550 56217
rect 54544 56177 54550 56189
rect 54602 56177 54608 56229
rect 54928 56217 54934 56229
rect 54889 56189 54934 56217
rect 54928 56177 54934 56189
rect 54986 56217 54992 56229
rect 55219 56220 55277 56226
rect 55219 56217 55231 56220
rect 54986 56189 55231 56217
rect 54986 56177 54992 56189
rect 55219 56186 55231 56189
rect 55265 56186 55277 56220
rect 55219 56180 55277 56186
rect 51242 56115 52094 56143
rect 51242 56103 51248 56115
rect 36976 56029 36982 56081
rect 37034 56069 37040 56081
rect 40816 56069 40822 56081
rect 37034 56041 40822 56069
rect 37034 56029 37040 56041
rect 40816 56029 40822 56041
rect 40874 56029 40880 56081
rect 1152 55970 58848 55992
rect 1152 55918 4294 55970
rect 4346 55918 4358 55970
rect 4410 55918 4422 55970
rect 4474 55918 4486 55970
rect 4538 55918 35014 55970
rect 35066 55918 35078 55970
rect 35130 55918 35142 55970
rect 35194 55918 35206 55970
rect 35258 55918 58848 55970
rect 1152 55896 58848 55918
rect 27346 55745 46334 55773
rect 1168 55659 1174 55711
rect 1226 55699 1232 55711
rect 1651 55702 1709 55708
rect 1651 55699 1663 55702
rect 1226 55671 1663 55699
rect 1226 55659 1232 55671
rect 1651 55668 1663 55671
rect 1697 55668 1709 55702
rect 1651 55662 1709 55668
rect 4435 55702 4493 55708
rect 4435 55668 4447 55702
rect 4481 55699 4493 55702
rect 4624 55699 4630 55711
rect 4481 55671 4630 55699
rect 4481 55668 4493 55671
rect 4435 55662 4493 55668
rect 4624 55659 4630 55671
rect 4682 55659 4688 55711
rect 7504 55659 7510 55711
rect 7562 55699 7568 55711
rect 7603 55702 7661 55708
rect 7603 55699 7615 55702
rect 7562 55671 7615 55699
rect 7562 55659 7568 55671
rect 7603 55668 7615 55671
rect 7649 55668 7661 55702
rect 7603 55662 7661 55668
rect 9136 55659 9142 55711
rect 9194 55699 9200 55711
rect 9331 55702 9389 55708
rect 9331 55699 9343 55702
rect 9194 55671 9343 55699
rect 9194 55659 9200 55671
rect 9331 55668 9343 55671
rect 9377 55668 9389 55702
rect 9331 55662 9389 55668
rect 13840 55659 13846 55711
rect 13898 55699 13904 55711
rect 13939 55702 13997 55708
rect 13939 55699 13951 55702
rect 13898 55671 13951 55699
rect 13898 55659 13904 55671
rect 13939 55668 13951 55671
rect 13985 55668 13997 55702
rect 13939 55662 13997 55668
rect 20176 55659 20182 55711
rect 20234 55699 20240 55711
rect 20371 55702 20429 55708
rect 20371 55699 20383 55702
rect 20234 55671 20383 55699
rect 20234 55659 20240 55671
rect 20371 55668 20383 55671
rect 20417 55668 20429 55702
rect 23440 55699 23446 55711
rect 23401 55671 23446 55699
rect 20371 55662 20429 55668
rect 23440 55659 23446 55671
rect 23498 55659 23504 55711
rect 24880 55659 24886 55711
rect 24938 55699 24944 55711
rect 25075 55702 25133 55708
rect 25075 55699 25087 55702
rect 24938 55671 25087 55699
rect 24938 55659 24944 55671
rect 25075 55668 25087 55671
rect 25121 55668 25133 55702
rect 25075 55662 25133 55668
rect 20560 55585 20566 55637
rect 20618 55625 20624 55637
rect 20618 55597 21086 55625
rect 20618 55585 20624 55597
rect 1747 55554 1805 55560
rect 1747 55520 1759 55554
rect 1793 55520 1805 55554
rect 1747 55514 1805 55520
rect 4243 55554 4301 55560
rect 4243 55520 4255 55554
rect 4289 55551 4301 55554
rect 4531 55554 4589 55560
rect 4531 55551 4543 55554
rect 4289 55523 4543 55551
rect 4289 55520 4301 55523
rect 4243 55514 4301 55520
rect 4531 55520 4543 55523
rect 4577 55551 4589 55554
rect 4624 55551 4630 55563
rect 4577 55523 4630 55551
rect 4577 55520 4589 55523
rect 4531 55514 4589 55520
rect 1762 55403 1790 55514
rect 4624 55511 4630 55523
rect 4682 55511 4688 55563
rect 7699 55554 7757 55560
rect 7699 55551 7711 55554
rect 7330 55523 7711 55551
rect 7330 55415 7358 55523
rect 7699 55520 7711 55523
rect 7745 55520 7757 55554
rect 9235 55554 9293 55560
rect 9235 55551 9247 55554
rect 7699 55514 7757 55520
rect 8962 55523 9247 55551
rect 8962 55415 8990 55523
rect 9235 55520 9247 55523
rect 9281 55520 9293 55554
rect 9235 55514 9293 55520
rect 14035 55554 14093 55560
rect 14035 55520 14047 55554
rect 14081 55551 14093 55554
rect 14128 55551 14134 55563
rect 14081 55523 14134 55551
rect 14081 55520 14093 55523
rect 14035 55514 14093 55520
rect 14128 55511 14134 55523
rect 14186 55511 14192 55563
rect 17779 55554 17837 55560
rect 17779 55551 17791 55554
rect 17410 55523 17791 55551
rect 17410 55415 17438 55523
rect 17779 55520 17791 55523
rect 17825 55520 17837 55554
rect 20275 55554 20333 55560
rect 20275 55551 20287 55554
rect 17779 55514 17837 55520
rect 20098 55523 20287 55551
rect 20098 55415 20126 55523
rect 20275 55520 20287 55523
rect 20321 55520 20333 55554
rect 20947 55554 21005 55560
rect 20947 55551 20959 55554
rect 20275 55514 20333 55520
rect 20770 55523 20959 55551
rect 20770 55415 20798 55523
rect 20947 55520 20959 55523
rect 20993 55520 21005 55554
rect 20947 55514 21005 55520
rect 21058 55477 21086 55597
rect 26128 55585 26134 55637
rect 26186 55625 26192 55637
rect 27346 55625 27374 55745
rect 39088 55659 39094 55711
rect 39146 55699 39152 55711
rect 39283 55702 39341 55708
rect 39283 55699 39295 55702
rect 39146 55671 39295 55699
rect 39146 55659 39152 55671
rect 39283 55668 39295 55671
rect 39329 55668 39341 55702
rect 39283 55662 39341 55668
rect 40720 55659 40726 55711
rect 40778 55699 40784 55711
rect 40819 55702 40877 55708
rect 40819 55699 40831 55702
rect 40778 55671 40831 55699
rect 40778 55659 40784 55671
rect 40819 55668 40831 55671
rect 40865 55668 40877 55702
rect 40819 55662 40877 55668
rect 45424 55659 45430 55711
rect 45482 55699 45488 55711
rect 46306 55708 46334 55745
rect 45619 55702 45677 55708
rect 45619 55699 45631 55702
rect 45482 55671 45631 55699
rect 45482 55659 45488 55671
rect 45619 55668 45631 55671
rect 45665 55668 45677 55702
rect 45619 55662 45677 55668
rect 46291 55702 46349 55708
rect 46291 55668 46303 55702
rect 46337 55668 46349 55702
rect 46291 55662 46349 55668
rect 46960 55659 46966 55711
rect 47018 55699 47024 55711
rect 47155 55702 47213 55708
rect 47155 55699 47167 55702
rect 47018 55671 47167 55699
rect 47018 55659 47024 55671
rect 47155 55668 47167 55671
rect 47201 55668 47213 55702
rect 47155 55662 47213 55668
rect 51760 55659 51766 55711
rect 51818 55699 51824 55711
rect 51859 55702 51917 55708
rect 51859 55699 51871 55702
rect 51818 55671 51871 55699
rect 51818 55659 51824 55671
rect 51859 55668 51871 55671
rect 51905 55668 51917 55702
rect 51859 55662 51917 55668
rect 56464 55659 56470 55711
rect 56522 55699 56528 55711
rect 56659 55702 56717 55708
rect 56659 55699 56671 55702
rect 56522 55671 56671 55699
rect 56522 55659 56528 55671
rect 56659 55668 56671 55671
rect 56705 55668 56717 55702
rect 56659 55662 56717 55668
rect 57520 55659 57526 55711
rect 57578 55699 57584 55711
rect 57715 55702 57773 55708
rect 57715 55699 57727 55702
rect 57578 55671 57727 55699
rect 57578 55659 57584 55671
rect 57715 55668 57727 55671
rect 57761 55668 57773 55702
rect 57715 55662 57773 55668
rect 26186 55597 27374 55625
rect 26186 55585 26192 55597
rect 45328 55585 45334 55637
rect 45386 55625 45392 55637
rect 46771 55628 46829 55634
rect 46771 55625 46783 55628
rect 45386 55597 46783 55625
rect 45386 55585 45392 55597
rect 46771 55594 46783 55597
rect 46817 55625 46829 55628
rect 47059 55628 47117 55634
rect 47059 55625 47071 55628
rect 46817 55597 47071 55625
rect 46817 55594 46829 55597
rect 46771 55588 46829 55594
rect 47059 55594 47071 55597
rect 47105 55594 47117 55628
rect 47059 55588 47117 55594
rect 23251 55554 23309 55560
rect 23251 55520 23263 55554
rect 23297 55551 23309 55554
rect 23539 55554 23597 55560
rect 23539 55551 23551 55554
rect 23297 55523 23551 55551
rect 23297 55520 23309 55523
rect 23251 55514 23309 55520
rect 23539 55520 23551 55523
rect 23585 55551 23597 55554
rect 24304 55551 24310 55563
rect 23585 55523 24310 55551
rect 23585 55520 23597 55523
rect 23539 55514 23597 55520
rect 24304 55511 24310 55523
rect 24362 55511 24368 55563
rect 24787 55554 24845 55560
rect 24787 55520 24799 55554
rect 24833 55551 24845 55554
rect 24976 55551 24982 55563
rect 24833 55523 24982 55551
rect 24833 55520 24845 55523
rect 24787 55514 24845 55520
rect 24976 55511 24982 55523
rect 25034 55511 25040 55563
rect 38995 55554 39053 55560
rect 38995 55520 39007 55554
rect 39041 55551 39053 55554
rect 39184 55551 39190 55563
rect 39041 55523 39190 55551
rect 39041 55520 39053 55523
rect 38995 55514 39053 55520
rect 39184 55511 39190 55523
rect 39242 55511 39248 55563
rect 39859 55554 39917 55560
rect 39859 55520 39871 55554
rect 39905 55520 39917 55554
rect 39859 55514 39917 55520
rect 39667 55480 39725 55486
rect 39667 55477 39679 55480
rect 21058 55449 39679 55477
rect 39667 55446 39679 55449
rect 39713 55477 39725 55480
rect 39874 55477 39902 55514
rect 40816 55511 40822 55563
rect 40874 55551 40880 55563
rect 40915 55554 40973 55560
rect 40915 55551 40927 55554
rect 40874 55523 40927 55551
rect 40874 55511 40880 55523
rect 40915 55520 40927 55523
rect 40961 55520 40973 55554
rect 40915 55514 40973 55520
rect 45523 55554 45581 55560
rect 45523 55520 45535 55554
rect 45569 55520 45581 55554
rect 51952 55551 51958 55563
rect 51913 55523 51958 55551
rect 45523 55514 45581 55520
rect 39713 55449 39902 55477
rect 39713 55446 39725 55449
rect 39667 55440 39725 55446
rect 1936 55403 1942 55415
rect 1762 55375 1942 55403
rect 1936 55363 1942 55375
rect 1994 55363 2000 55415
rect 7312 55403 7318 55415
rect 7273 55375 7318 55403
rect 7312 55363 7318 55375
rect 7370 55363 7376 55415
rect 8944 55403 8950 55415
rect 8905 55375 8950 55403
rect 8944 55363 8950 55375
rect 9002 55363 9008 55415
rect 17392 55403 17398 55415
rect 17353 55375 17398 55403
rect 17392 55363 17398 55375
rect 17450 55363 17456 55415
rect 20080 55403 20086 55415
rect 20041 55375 20086 55403
rect 20080 55363 20086 55375
rect 20138 55363 20144 55415
rect 20752 55403 20758 55415
rect 20713 55375 20758 55403
rect 20752 55363 20758 55375
rect 20810 55363 20816 55415
rect 45331 55406 45389 55412
rect 45331 55372 45343 55406
rect 45377 55403 45389 55406
rect 45538 55403 45566 55514
rect 51952 55511 51958 55523
rect 52010 55511 52016 55563
rect 55795 55554 55853 55560
rect 55795 55551 55807 55554
rect 55618 55523 55807 55551
rect 55618 55415 55646 55523
rect 55795 55520 55807 55523
rect 55841 55520 55853 55554
rect 55795 55514 55853 55520
rect 56563 55554 56621 55560
rect 56563 55520 56575 55554
rect 56609 55520 56621 55554
rect 57619 55554 57677 55560
rect 57619 55551 57631 55554
rect 56563 55514 56621 55520
rect 57346 55523 57631 55551
rect 45808 55403 45814 55415
rect 45377 55375 45814 55403
rect 45377 55372 45389 55375
rect 45331 55366 45389 55372
rect 45808 55363 45814 55375
rect 45866 55363 45872 55415
rect 55600 55403 55606 55415
rect 55561 55375 55606 55403
rect 55600 55363 55606 55375
rect 55658 55363 55664 55415
rect 56272 55403 56278 55415
rect 56233 55375 56278 55403
rect 56272 55363 56278 55375
rect 56330 55403 56336 55415
rect 56578 55403 56606 55514
rect 57346 55415 57374 55523
rect 57619 55520 57631 55523
rect 57665 55520 57677 55554
rect 57619 55514 57677 55520
rect 57328 55403 57334 55415
rect 56330 55375 56606 55403
rect 57289 55375 57334 55403
rect 56330 55363 56336 55375
rect 57328 55363 57334 55375
rect 57386 55363 57392 55415
rect 1152 55304 58848 55326
rect 1152 55252 19654 55304
rect 19706 55252 19718 55304
rect 19770 55252 19782 55304
rect 19834 55252 19846 55304
rect 19898 55252 50374 55304
rect 50426 55252 50438 55304
rect 50490 55252 50502 55304
rect 50554 55252 50566 55304
rect 50618 55252 58848 55304
rect 1152 55230 58848 55252
rect 57907 55184 57965 55190
rect 57907 55150 57919 55184
rect 57953 55181 57965 55184
rect 59152 55181 59158 55193
rect 57953 55153 59158 55181
rect 57953 55150 57965 55153
rect 57907 55144 57965 55150
rect 59152 55141 59158 55153
rect 59210 55141 59216 55193
rect 15088 55067 15094 55119
rect 15146 55107 15152 55119
rect 55600 55107 55606 55119
rect 15146 55079 55606 55107
rect 15146 55067 15152 55079
rect 55600 55067 55606 55079
rect 55658 55067 55664 55119
rect 42352 55033 42358 55045
rect 42313 55005 42358 55033
rect 42352 54993 42358 55005
rect 42410 54993 42416 55045
rect 57619 54888 57677 54894
rect 57619 54854 57631 54888
rect 57665 54885 57677 54888
rect 57808 54885 57814 54897
rect 57665 54857 57814 54885
rect 57665 54854 57677 54857
rect 57619 54848 57677 54854
rect 57808 54845 57814 54857
rect 57866 54845 57872 54897
rect 5008 54771 5014 54823
rect 5066 54811 5072 54823
rect 25651 54814 25709 54820
rect 25651 54811 25663 54814
rect 5066 54783 25663 54811
rect 5066 54771 5072 54783
rect 25651 54780 25663 54783
rect 25697 54780 25709 54814
rect 25651 54774 25709 54780
rect 7219 54740 7277 54746
rect 7219 54706 7231 54740
rect 7265 54737 7277 54740
rect 7507 54740 7565 54746
rect 7507 54737 7519 54740
rect 7265 54709 7519 54737
rect 7265 54706 7277 54709
rect 7219 54700 7277 54706
rect 7507 54706 7519 54709
rect 7553 54737 7565 54740
rect 15280 54737 15286 54749
rect 7553 54709 15286 54737
rect 7553 54706 7565 54709
rect 7507 54700 7565 54706
rect 15280 54697 15286 54709
rect 15338 54697 15344 54749
rect 20179 54740 20237 54746
rect 20179 54706 20191 54740
rect 20225 54737 20237 54740
rect 20464 54737 20470 54749
rect 20225 54709 20470 54737
rect 20225 54706 20237 54709
rect 20179 54700 20237 54706
rect 20464 54697 20470 54709
rect 20522 54697 20528 54749
rect 22384 54737 22390 54749
rect 22345 54709 22390 54737
rect 22384 54697 22390 54709
rect 22442 54737 22448 54749
rect 22771 54740 22829 54746
rect 22771 54737 22783 54740
rect 22442 54709 22783 54737
rect 22442 54697 22448 54709
rect 22771 54706 22783 54709
rect 22817 54706 22829 54740
rect 22771 54700 22829 54706
rect 1152 54638 58848 54660
rect 1152 54586 4294 54638
rect 4346 54586 4358 54638
rect 4410 54586 4422 54638
rect 4474 54586 4486 54638
rect 4538 54586 35014 54638
rect 35066 54586 35078 54638
rect 35130 54586 35142 54638
rect 35194 54586 35206 54638
rect 35258 54586 58848 54638
rect 1152 54564 58848 54586
rect 57907 54370 57965 54376
rect 57907 54336 57919 54370
rect 57953 54367 57965 54370
rect 58096 54367 58102 54379
rect 57953 54339 58102 54367
rect 57953 54336 57965 54339
rect 57907 54330 57965 54336
rect 58096 54327 58102 54339
rect 58154 54327 58160 54379
rect 57811 54222 57869 54228
rect 57811 54188 57823 54222
rect 57857 54188 57869 54222
rect 57811 54182 57869 54188
rect 57619 54074 57677 54080
rect 57619 54040 57631 54074
rect 57665 54071 57677 54074
rect 57826 54071 57854 54182
rect 58096 54071 58102 54083
rect 57665 54043 58102 54071
rect 57665 54040 57677 54043
rect 57619 54034 57677 54040
rect 58096 54031 58102 54043
rect 58154 54031 58160 54083
rect 1152 53972 58848 53994
rect 1152 53920 19654 53972
rect 19706 53920 19718 53972
rect 19770 53920 19782 53972
rect 19834 53920 19846 53972
rect 19898 53920 50374 53972
rect 50426 53920 50438 53972
rect 50490 53920 50502 53972
rect 50554 53920 50566 53972
rect 50618 53920 58848 53972
rect 1152 53898 58848 53920
rect 57907 53852 57965 53858
rect 57907 53818 57919 53852
rect 57953 53849 57965 53852
rect 59632 53849 59638 53861
rect 57953 53821 59638 53849
rect 57953 53818 57965 53821
rect 57907 53812 57965 53818
rect 59632 53809 59638 53821
rect 59690 53809 59696 53861
rect 57811 53556 57869 53562
rect 57811 53522 57823 53556
rect 57857 53522 57869 53556
rect 57811 53516 57869 53522
rect 57619 53408 57677 53414
rect 57619 53374 57631 53408
rect 57665 53405 57677 53408
rect 57712 53405 57718 53417
rect 57665 53377 57718 53405
rect 57665 53374 57677 53377
rect 57619 53368 57677 53374
rect 57712 53365 57718 53377
rect 57770 53405 57776 53417
rect 57826 53405 57854 53516
rect 58099 53408 58157 53414
rect 58099 53405 58111 53408
rect 57770 53377 58111 53405
rect 57770 53365 57776 53377
rect 58099 53374 58111 53377
rect 58145 53374 58157 53408
rect 58099 53368 58157 53374
rect 1152 53306 58848 53328
rect 1152 53254 4294 53306
rect 4346 53254 4358 53306
rect 4410 53254 4422 53306
rect 4474 53254 4486 53306
rect 4538 53254 35014 53306
rect 35066 53254 35078 53306
rect 35130 53254 35142 53306
rect 35194 53254 35206 53306
rect 35258 53254 58848 53306
rect 1152 53232 58848 53254
rect 29971 53038 30029 53044
rect 29971 53004 29983 53038
rect 30017 53035 30029 53038
rect 35344 53035 35350 53047
rect 30017 53007 35350 53035
rect 30017 53004 30029 53007
rect 29971 52998 30029 53004
rect 35344 52995 35350 53007
rect 35402 52995 35408 53047
rect 1747 52890 1805 52896
rect 1747 52856 1759 52890
rect 1793 52887 1805 52890
rect 2035 52890 2093 52896
rect 2035 52887 2047 52890
rect 1793 52859 2047 52887
rect 1793 52856 1805 52859
rect 1747 52850 1805 52856
rect 2035 52856 2047 52859
rect 2081 52887 2093 52890
rect 14992 52887 14998 52899
rect 2081 52859 14998 52887
rect 2081 52856 2093 52859
rect 2035 52850 2093 52856
rect 14992 52847 14998 52859
rect 15050 52847 15056 52899
rect 26896 52847 26902 52899
rect 26954 52887 26960 52899
rect 51475 52890 51533 52896
rect 51475 52887 51487 52890
rect 26954 52859 51487 52887
rect 26954 52847 26960 52859
rect 51475 52856 51487 52859
rect 51521 52856 51533 52890
rect 51475 52850 51533 52856
rect 1152 52640 58848 52662
rect 1152 52588 19654 52640
rect 19706 52588 19718 52640
rect 19770 52588 19782 52640
rect 19834 52588 19846 52640
rect 19898 52588 50374 52640
rect 50426 52588 50438 52640
rect 50490 52588 50502 52640
rect 50554 52588 50566 52640
rect 50618 52588 58848 52640
rect 1152 52566 58848 52588
rect 1152 51974 58848 51996
rect 1152 51922 4294 51974
rect 4346 51922 4358 51974
rect 4410 51922 4422 51974
rect 4474 51922 4486 51974
rect 4538 51922 35014 51974
rect 35066 51922 35078 51974
rect 35130 51922 35142 51974
rect 35194 51922 35206 51974
rect 35258 51922 58848 51974
rect 1152 51900 58848 51922
rect 2515 51558 2573 51564
rect 2515 51524 2527 51558
rect 2561 51555 2573 51558
rect 2803 51558 2861 51564
rect 2803 51555 2815 51558
rect 2561 51527 2815 51555
rect 2561 51524 2573 51527
rect 2515 51518 2573 51524
rect 2803 51524 2815 51527
rect 2849 51555 2861 51558
rect 19408 51555 19414 51567
rect 2849 51527 19414 51555
rect 2849 51524 2861 51527
rect 2803 51518 2861 51524
rect 19408 51515 19414 51527
rect 19466 51515 19472 51567
rect 43891 51410 43949 51416
rect 43891 51376 43903 51410
rect 43937 51407 43949 51410
rect 54544 51407 54550 51419
rect 43937 51379 54550 51407
rect 43937 51376 43949 51379
rect 43891 51370 43949 51376
rect 54544 51367 54550 51379
rect 54602 51367 54608 51419
rect 1152 51308 58848 51330
rect 1152 51256 19654 51308
rect 19706 51256 19718 51308
rect 19770 51256 19782 51308
rect 19834 51256 19846 51308
rect 19898 51256 50374 51308
rect 50426 51256 50438 51308
rect 50490 51256 50502 51308
rect 50554 51256 50566 51308
rect 50618 51256 58848 51308
rect 1152 51234 58848 51256
rect 12496 51185 12502 51197
rect 12457 51157 12502 51185
rect 12496 51145 12502 51157
rect 12554 51145 12560 51197
rect 11920 50849 11926 50901
rect 11978 50889 11984 50901
rect 31987 50892 32045 50898
rect 31987 50889 31999 50892
rect 11978 50861 31999 50889
rect 11978 50849 11984 50861
rect 31987 50858 31999 50861
rect 32033 50858 32045 50892
rect 31987 50852 32045 50858
rect 37363 50744 37421 50750
rect 37363 50710 37375 50744
rect 37409 50741 37421 50744
rect 37651 50744 37709 50750
rect 37651 50741 37663 50744
rect 37409 50713 37663 50741
rect 37409 50710 37421 50713
rect 37363 50704 37421 50710
rect 37651 50710 37663 50713
rect 37697 50741 37709 50744
rect 55024 50741 55030 50753
rect 37697 50713 55030 50741
rect 37697 50710 37709 50713
rect 37651 50704 37709 50710
rect 55024 50701 55030 50713
rect 55082 50701 55088 50753
rect 56848 50701 56854 50753
rect 56906 50741 56912 50753
rect 56947 50744 57005 50750
rect 56947 50741 56959 50744
rect 56906 50713 56959 50741
rect 56906 50701 56912 50713
rect 56947 50710 56959 50713
rect 56993 50741 57005 50744
rect 57139 50744 57197 50750
rect 57139 50741 57151 50744
rect 56993 50713 57151 50741
rect 56993 50710 57005 50713
rect 56947 50704 57005 50710
rect 57139 50710 57151 50713
rect 57185 50710 57197 50744
rect 57139 50704 57197 50710
rect 1152 50642 58848 50664
rect 1152 50590 4294 50642
rect 4346 50590 4358 50642
rect 4410 50590 4422 50642
rect 4474 50590 4486 50642
rect 4538 50590 35014 50642
rect 35066 50590 35078 50642
rect 35130 50590 35142 50642
rect 35194 50590 35206 50642
rect 35258 50590 58848 50642
rect 1152 50568 58848 50590
rect 4147 50448 4205 50454
rect 4147 50414 4159 50448
rect 4193 50445 4205 50448
rect 54928 50445 54934 50457
rect 4193 50417 54934 50445
rect 4193 50414 4205 50417
rect 4147 50408 4205 50414
rect 54928 50405 54934 50417
rect 54986 50405 54992 50457
rect 40915 50226 40973 50232
rect 40915 50192 40927 50226
rect 40961 50192 40973 50226
rect 40915 50186 40973 50192
rect 40930 50087 40958 50186
rect 40819 50078 40877 50084
rect 40819 50044 40831 50078
rect 40865 50075 40877 50078
rect 40912 50075 40918 50087
rect 40865 50047 40918 50075
rect 40865 50044 40877 50047
rect 40819 50038 40877 50044
rect 40912 50035 40918 50047
rect 40970 50035 40976 50087
rect 1152 49976 58848 49998
rect 1152 49924 19654 49976
rect 19706 49924 19718 49976
rect 19770 49924 19782 49976
rect 19834 49924 19846 49976
rect 19898 49924 50374 49976
rect 50426 49924 50438 49976
rect 50490 49924 50502 49976
rect 50554 49924 50566 49976
rect 50618 49924 58848 49976
rect 1152 49902 58848 49924
rect 6259 49560 6317 49566
rect 6259 49526 6271 49560
rect 6305 49557 6317 49560
rect 32464 49557 32470 49569
rect 6305 49529 32470 49557
rect 6305 49526 6317 49529
rect 6259 49520 6317 49526
rect 32464 49517 32470 49529
rect 32522 49517 32528 49569
rect 44848 49409 44854 49421
rect 44809 49381 44854 49409
rect 44848 49369 44854 49381
rect 44906 49409 44912 49421
rect 45235 49412 45293 49418
rect 45235 49409 45247 49412
rect 44906 49381 45247 49409
rect 44906 49369 44912 49381
rect 45235 49378 45247 49381
rect 45281 49378 45293 49412
rect 45235 49372 45293 49378
rect 48019 49412 48077 49418
rect 48019 49378 48031 49412
rect 48065 49409 48077 49412
rect 48112 49409 48118 49421
rect 48065 49381 48118 49409
rect 48065 49378 48077 49381
rect 48019 49372 48077 49378
rect 48112 49369 48118 49381
rect 48170 49369 48176 49421
rect 1152 49310 58848 49332
rect 1152 49258 4294 49310
rect 4346 49258 4358 49310
rect 4410 49258 4422 49310
rect 4474 49258 4486 49310
rect 4538 49258 35014 49310
rect 35066 49258 35078 49310
rect 35130 49258 35142 49310
rect 35194 49258 35206 49310
rect 35258 49258 58848 49310
rect 1152 49236 58848 49258
rect 7216 48999 7222 49051
rect 7274 49039 7280 49051
rect 7274 49011 7319 49039
rect 7274 48999 7280 49011
rect 1747 48894 1805 48900
rect 1747 48860 1759 48894
rect 1793 48860 1805 48894
rect 1747 48854 1805 48860
rect 1762 48743 1790 48854
rect 29680 48851 29686 48903
rect 29738 48891 29744 48903
rect 41395 48894 41453 48900
rect 41395 48891 41407 48894
rect 29738 48863 41407 48891
rect 29738 48851 29744 48863
rect 41395 48860 41407 48863
rect 41441 48891 41453 48894
rect 41587 48894 41645 48900
rect 41587 48891 41599 48894
rect 41441 48863 41599 48891
rect 41441 48860 41453 48863
rect 41395 48854 41453 48860
rect 41587 48860 41599 48863
rect 41633 48860 41645 48894
rect 41587 48854 41645 48860
rect 1939 48746 1997 48752
rect 1939 48743 1951 48746
rect 1762 48715 1951 48743
rect 1939 48712 1951 48715
rect 1985 48743 1997 48746
rect 3568 48743 3574 48755
rect 1985 48715 3574 48743
rect 1985 48712 1997 48715
rect 1939 48706 1997 48712
rect 3568 48703 3574 48715
rect 3626 48703 3632 48755
rect 28531 48746 28589 48752
rect 28531 48712 28543 48746
rect 28577 48743 28589 48746
rect 43504 48743 43510 48755
rect 28577 48715 43510 48743
rect 28577 48712 28589 48715
rect 28531 48706 28589 48712
rect 43504 48703 43510 48715
rect 43562 48703 43568 48755
rect 1152 48644 58848 48666
rect 1152 48592 19654 48644
rect 19706 48592 19718 48644
rect 19770 48592 19782 48644
rect 19834 48592 19846 48644
rect 19898 48592 50374 48644
rect 50426 48592 50438 48644
rect 50490 48592 50502 48644
rect 50554 48592 50566 48644
rect 50618 48592 58848 48644
rect 1152 48570 58848 48592
rect 4243 48080 4301 48086
rect 4243 48046 4255 48080
rect 4289 48077 4301 48080
rect 4531 48080 4589 48086
rect 4531 48077 4543 48080
rect 4289 48049 4543 48077
rect 4289 48046 4301 48049
rect 4243 48040 4301 48046
rect 4531 48046 4543 48049
rect 4577 48077 4589 48080
rect 4720 48077 4726 48089
rect 4577 48049 4726 48077
rect 4577 48046 4589 48049
rect 4531 48040 4589 48046
rect 4720 48037 4726 48049
rect 4778 48037 4784 48089
rect 48880 48037 48886 48089
rect 48938 48077 48944 48089
rect 58003 48080 58061 48086
rect 58003 48077 58015 48080
rect 48938 48049 58015 48077
rect 48938 48037 48944 48049
rect 58003 48046 58015 48049
rect 58049 48046 58061 48080
rect 58003 48040 58061 48046
rect 1152 47978 58848 48000
rect 1152 47926 4294 47978
rect 4346 47926 4358 47978
rect 4410 47926 4422 47978
rect 4474 47926 4486 47978
rect 4538 47926 35014 47978
rect 35066 47926 35078 47978
rect 35130 47926 35142 47978
rect 35194 47926 35206 47978
rect 35258 47926 58848 47978
rect 1152 47904 58848 47926
rect 17395 47636 17453 47642
rect 17395 47602 17407 47636
rect 17441 47633 17453 47636
rect 17683 47636 17741 47642
rect 17683 47633 17695 47636
rect 17441 47605 17695 47633
rect 17441 47602 17453 47605
rect 17395 47596 17453 47602
rect 17683 47602 17695 47605
rect 17729 47633 17741 47636
rect 39664 47633 39670 47645
rect 17729 47605 39670 47633
rect 17729 47602 17741 47605
rect 17683 47596 17741 47602
rect 39664 47593 39670 47605
rect 39722 47593 39728 47645
rect 23539 47562 23597 47568
rect 23539 47528 23551 47562
rect 23585 47559 23597 47562
rect 48208 47559 48214 47571
rect 23585 47531 48214 47559
rect 23585 47528 23597 47531
rect 23539 47522 23597 47528
rect 48208 47519 48214 47531
rect 48266 47519 48272 47571
rect 1152 47312 58848 47334
rect 1152 47260 19654 47312
rect 19706 47260 19718 47312
rect 19770 47260 19782 47312
rect 19834 47260 19846 47312
rect 19898 47260 50374 47312
rect 50426 47260 50438 47312
rect 50490 47260 50502 47312
rect 50554 47260 50566 47312
rect 50618 47260 58848 47312
rect 1152 47238 58848 47260
rect 31699 46896 31757 46902
rect 31699 46862 31711 46896
rect 31745 46893 31757 46896
rect 43888 46893 43894 46905
rect 31745 46865 43894 46893
rect 31745 46862 31757 46865
rect 31699 46856 31757 46862
rect 43888 46853 43894 46865
rect 43946 46853 43952 46905
rect 13651 46822 13709 46828
rect 13651 46788 13663 46822
rect 13697 46819 13709 46822
rect 13939 46822 13997 46828
rect 13939 46819 13951 46822
rect 13697 46791 13951 46819
rect 13697 46788 13709 46791
rect 13651 46782 13709 46788
rect 13939 46788 13951 46791
rect 13985 46819 13997 46822
rect 16624 46819 16630 46831
rect 13985 46791 16630 46819
rect 13985 46788 13997 46791
rect 13939 46782 13997 46788
rect 16624 46779 16630 46791
rect 16682 46779 16688 46831
rect 4531 46748 4589 46754
rect 4531 46714 4543 46748
rect 4577 46745 4589 46748
rect 4816 46745 4822 46757
rect 4577 46717 4822 46745
rect 4577 46714 4589 46717
rect 4531 46708 4589 46714
rect 4816 46705 4822 46717
rect 4874 46705 4880 46757
rect 15379 46748 15437 46754
rect 15379 46714 15391 46748
rect 15425 46745 15437 46748
rect 15667 46748 15725 46754
rect 15667 46745 15679 46748
rect 15425 46717 15679 46745
rect 15425 46714 15437 46717
rect 15379 46708 15437 46714
rect 15667 46714 15679 46717
rect 15713 46745 15725 46748
rect 19984 46745 19990 46757
rect 15713 46717 19990 46745
rect 15713 46714 15725 46717
rect 15667 46708 15725 46714
rect 19984 46705 19990 46717
rect 20042 46705 20048 46757
rect 45331 46748 45389 46754
rect 45331 46714 45343 46748
rect 45377 46745 45389 46748
rect 45424 46745 45430 46757
rect 45377 46717 45430 46745
rect 45377 46714 45389 46717
rect 45331 46708 45389 46714
rect 45424 46705 45430 46717
rect 45482 46705 45488 46757
rect 1152 46646 58848 46668
rect 1152 46594 4294 46646
rect 4346 46594 4358 46646
rect 4410 46594 4422 46646
rect 4474 46594 4486 46646
rect 4538 46594 35014 46646
rect 35066 46594 35078 46646
rect 35130 46594 35142 46646
rect 35194 46594 35206 46646
rect 35258 46594 58848 46646
rect 1152 46572 58848 46594
rect 4816 46483 4822 46535
rect 4874 46523 4880 46535
rect 57136 46523 57142 46535
rect 4874 46495 57142 46523
rect 4874 46483 4880 46495
rect 57136 46483 57142 46495
rect 57194 46483 57200 46535
rect 28243 46230 28301 46236
rect 28243 46196 28255 46230
rect 28289 46196 28301 46230
rect 28243 46190 28301 46196
rect 27952 46153 27958 46165
rect 27913 46125 27958 46153
rect 27952 46113 27958 46125
rect 28010 46153 28016 46165
rect 28258 46153 28286 46190
rect 28010 46125 28286 46153
rect 28010 46113 28016 46125
rect 40243 46082 40301 46088
rect 40243 46048 40255 46082
rect 40289 46079 40301 46082
rect 46960 46079 46966 46091
rect 40289 46051 46966 46079
rect 40289 46048 40301 46051
rect 40243 46042 40301 46048
rect 46960 46039 46966 46051
rect 47018 46039 47024 46091
rect 1152 45980 58848 46002
rect 1152 45928 19654 45980
rect 19706 45928 19718 45980
rect 19770 45928 19782 45980
rect 19834 45928 19846 45980
rect 19898 45928 50374 45980
rect 50426 45928 50438 45980
rect 50490 45928 50502 45980
rect 50554 45928 50566 45980
rect 50618 45928 58848 45980
rect 1152 45906 58848 45928
rect 20464 45373 20470 45425
rect 20522 45413 20528 45425
rect 31600 45413 31606 45425
rect 20522 45385 31606 45413
rect 20522 45373 20528 45385
rect 31600 45373 31606 45385
rect 31658 45373 31664 45425
rect 1152 45314 58848 45336
rect 1152 45262 4294 45314
rect 4346 45262 4358 45314
rect 4410 45262 4422 45314
rect 4474 45262 4486 45314
rect 4538 45262 35014 45314
rect 35066 45262 35078 45314
rect 35130 45262 35142 45314
rect 35194 45262 35206 45314
rect 35258 45262 58848 45314
rect 1152 45240 58848 45262
rect 12112 44855 12118 44907
rect 12170 44895 12176 44907
rect 38899 44898 38957 44904
rect 38899 44895 38911 44898
rect 12170 44867 38911 44895
rect 12170 44855 12176 44867
rect 38899 44864 38911 44867
rect 38945 44895 38957 44898
rect 39091 44898 39149 44904
rect 39091 44895 39103 44898
rect 38945 44867 39103 44895
rect 38945 44864 38957 44867
rect 38899 44858 38957 44864
rect 39091 44864 39103 44867
rect 39137 44864 39149 44898
rect 39091 44858 39149 44864
rect 1152 44648 58848 44670
rect 1152 44596 19654 44648
rect 19706 44596 19718 44648
rect 19770 44596 19782 44648
rect 19834 44596 19846 44648
rect 19898 44596 50374 44648
rect 50426 44596 50438 44648
rect 50490 44596 50502 44648
rect 50554 44596 50566 44648
rect 50618 44596 58848 44648
rect 1152 44574 58848 44596
rect 17968 44041 17974 44093
rect 18026 44081 18032 44093
rect 46771 44084 46829 44090
rect 46771 44081 46783 44084
rect 18026 44053 46783 44081
rect 18026 44041 18032 44053
rect 46771 44050 46783 44053
rect 46817 44081 46829 44084
rect 46963 44084 47021 44090
rect 46963 44081 46975 44084
rect 46817 44053 46975 44081
rect 46817 44050 46829 44053
rect 46771 44044 46829 44050
rect 46963 44050 46975 44053
rect 47009 44050 47021 44084
rect 47728 44081 47734 44093
rect 47641 44053 47734 44081
rect 46963 44044 47021 44050
rect 47728 44041 47734 44053
rect 47786 44081 47792 44093
rect 47827 44084 47885 44090
rect 47827 44081 47839 44084
rect 47786 44053 47839 44081
rect 47786 44041 47792 44053
rect 47827 44050 47839 44053
rect 47873 44050 47885 44084
rect 47827 44044 47885 44050
rect 1152 43982 58848 44004
rect 1152 43930 4294 43982
rect 4346 43930 4358 43982
rect 4410 43930 4422 43982
rect 4474 43930 4486 43982
rect 4538 43930 35014 43982
rect 35066 43930 35078 43982
rect 35130 43930 35142 43982
rect 35194 43930 35206 43982
rect 35258 43930 58848 43982
rect 1152 43908 58848 43930
rect 25648 43819 25654 43871
rect 25706 43859 25712 43871
rect 47728 43859 47734 43871
rect 25706 43831 47734 43859
rect 25706 43819 25712 43831
rect 47728 43819 47734 43831
rect 47786 43819 47792 43871
rect 37075 43640 37133 43646
rect 37075 43606 37087 43640
rect 37121 43637 37133 43640
rect 37363 43640 37421 43646
rect 37363 43637 37375 43640
rect 37121 43609 37375 43637
rect 37121 43606 37133 43609
rect 37075 43600 37133 43606
rect 37363 43606 37375 43609
rect 37409 43637 37421 43640
rect 54064 43637 54070 43649
rect 37409 43609 54070 43637
rect 37409 43606 37421 43609
rect 37363 43600 37421 43606
rect 54064 43597 54070 43609
rect 54122 43597 54128 43649
rect 13648 43523 13654 43575
rect 13706 43563 13712 43575
rect 13747 43566 13805 43572
rect 13747 43563 13759 43566
rect 13706 43535 13759 43563
rect 13706 43523 13712 43535
rect 13747 43532 13759 43535
rect 13793 43532 13805 43566
rect 38611 43566 38669 43572
rect 38611 43563 38623 43566
rect 13747 43526 13805 43532
rect 38434 43535 38623 43563
rect 27346 43461 37454 43489
rect 22288 43375 22294 43427
rect 22346 43415 22352 43427
rect 27346 43415 27374 43461
rect 22346 43387 27374 43415
rect 37426 43415 37454 43461
rect 38434 43424 38462 43535
rect 38611 43532 38623 43535
rect 38657 43532 38669 43566
rect 38611 43526 38669 43532
rect 52051 43566 52109 43572
rect 52051 43532 52063 43566
rect 52097 43563 52109 43566
rect 52240 43563 52246 43575
rect 52097 43535 52246 43563
rect 52097 43532 52109 43535
rect 52051 43526 52109 43532
rect 52240 43523 52246 43535
rect 52298 43523 52304 43575
rect 38419 43418 38477 43424
rect 38419 43415 38431 43418
rect 37426 43387 38431 43415
rect 22346 43375 22352 43387
rect 38419 43384 38431 43387
rect 38465 43384 38477 43418
rect 38419 43378 38477 43384
rect 1152 43316 58848 43338
rect 1152 43264 19654 43316
rect 19706 43264 19718 43316
rect 19770 43264 19782 43316
rect 19834 43264 19846 43316
rect 19898 43264 50374 43316
rect 50426 43264 50438 43316
rect 50490 43264 50502 43316
rect 50554 43264 50566 43316
rect 50618 43264 58848 43316
rect 1152 43242 58848 43264
rect 11440 42783 11446 42835
rect 11498 42823 11504 42835
rect 11498 42795 27374 42823
rect 11498 42783 11504 42795
rect 10963 42752 11021 42758
rect 10963 42718 10975 42752
rect 11009 42749 11021 42752
rect 11251 42752 11309 42758
rect 11251 42749 11263 42752
rect 11009 42721 11263 42749
rect 11009 42718 11021 42721
rect 10963 42712 11021 42718
rect 11251 42718 11263 42721
rect 11297 42749 11309 42752
rect 11344 42749 11350 42761
rect 11297 42721 11350 42749
rect 11297 42718 11309 42721
rect 11251 42712 11309 42718
rect 11344 42709 11350 42721
rect 11402 42709 11408 42761
rect 25936 42749 25942 42761
rect 25897 42721 25942 42749
rect 25936 42709 25942 42721
rect 25994 42749 26000 42761
rect 26227 42752 26285 42758
rect 26227 42749 26239 42752
rect 25994 42721 26239 42749
rect 25994 42709 26000 42721
rect 26227 42718 26239 42721
rect 26273 42718 26285 42752
rect 27346 42749 27374 42795
rect 45235 42752 45293 42758
rect 45235 42749 45247 42752
rect 27346 42721 45247 42749
rect 26227 42712 26285 42718
rect 45235 42718 45247 42721
rect 45281 42749 45293 42752
rect 45427 42752 45485 42758
rect 45427 42749 45439 42752
rect 45281 42721 45439 42749
rect 45281 42718 45293 42721
rect 45235 42712 45293 42718
rect 45427 42718 45439 42721
rect 45473 42718 45485 42752
rect 45427 42712 45485 42718
rect 1152 42650 58848 42672
rect 1152 42598 4294 42650
rect 4346 42598 4358 42650
rect 4410 42598 4422 42650
rect 4474 42598 4486 42650
rect 4538 42598 35014 42650
rect 35066 42598 35078 42650
rect 35130 42598 35142 42650
rect 35194 42598 35206 42650
rect 35258 42598 58848 42650
rect 1152 42576 58848 42598
rect 11344 42487 11350 42539
rect 11402 42527 11408 42539
rect 26128 42527 26134 42539
rect 11402 42499 26134 42527
rect 11402 42487 11408 42499
rect 26128 42487 26134 42499
rect 26186 42487 26192 42539
rect 14128 42265 14134 42317
rect 14186 42305 14192 42317
rect 14186 42277 17294 42305
rect 14186 42265 14192 42277
rect 16243 42234 16301 42240
rect 16243 42200 16255 42234
rect 16289 42231 16301 42234
rect 16528 42231 16534 42243
rect 16289 42203 16534 42231
rect 16289 42200 16301 42203
rect 16243 42194 16301 42200
rect 16528 42191 16534 42203
rect 16586 42191 16592 42243
rect 17266 42231 17294 42277
rect 48211 42234 48269 42240
rect 48211 42231 48223 42234
rect 17266 42203 48223 42231
rect 48211 42200 48223 42203
rect 48257 42200 48269 42234
rect 48211 42194 48269 42200
rect 1152 41984 58848 42006
rect 1152 41932 19654 41984
rect 19706 41932 19718 41984
rect 19770 41932 19782 41984
rect 19834 41932 19846 41984
rect 19898 41932 50374 41984
rect 50426 41932 50438 41984
rect 50490 41932 50502 41984
rect 50554 41932 50566 41984
rect 50618 41932 58848 41984
rect 1152 41910 58848 41932
rect 22960 41747 22966 41799
rect 23018 41787 23024 41799
rect 38995 41790 39053 41796
rect 38995 41787 39007 41790
rect 23018 41759 39007 41787
rect 23018 41747 23024 41759
rect 38995 41756 39007 41759
rect 39041 41756 39053 41790
rect 38995 41750 39053 41756
rect 25168 41377 25174 41429
rect 25226 41417 25232 41429
rect 33235 41420 33293 41426
rect 33235 41417 33247 41420
rect 25226 41389 33247 41417
rect 25226 41377 25232 41389
rect 33235 41386 33247 41389
rect 33281 41417 33293 41420
rect 33427 41420 33485 41426
rect 33427 41417 33439 41420
rect 33281 41389 33439 41417
rect 33281 41386 33293 41389
rect 33235 41380 33293 41386
rect 33427 41386 33439 41389
rect 33473 41386 33485 41420
rect 33427 41380 33485 41386
rect 1152 41318 58848 41340
rect 1152 41266 4294 41318
rect 4346 41266 4358 41318
rect 4410 41266 4422 41318
rect 4474 41266 4486 41318
rect 4538 41266 35014 41318
rect 35066 41266 35078 41318
rect 35130 41266 35142 41318
rect 35194 41266 35206 41318
rect 35258 41266 58848 41318
rect 1152 41244 58848 41266
rect 33523 40976 33581 40982
rect 33523 40942 33535 40976
rect 33569 40973 33581 40976
rect 33569 40945 37454 40973
rect 33569 40942 33581 40945
rect 33523 40936 33581 40942
rect 1843 40902 1901 40908
rect 1843 40868 1855 40902
rect 1889 40899 1901 40902
rect 2035 40902 2093 40908
rect 2035 40899 2047 40902
rect 1889 40871 2047 40899
rect 1889 40868 1901 40871
rect 1843 40862 1901 40868
rect 2035 40868 2047 40871
rect 2081 40899 2093 40902
rect 28912 40899 28918 40911
rect 2081 40871 28918 40899
rect 2081 40868 2093 40871
rect 2035 40862 2093 40868
rect 28912 40859 28918 40871
rect 28970 40859 28976 40911
rect 34099 40902 34157 40908
rect 34099 40868 34111 40902
rect 34145 40868 34157 40902
rect 37426 40899 37454 40945
rect 48304 40899 48310 40911
rect 37426 40871 48310 40899
rect 34099 40862 34157 40868
rect 33904 40751 33910 40763
rect 33865 40723 33910 40751
rect 33904 40711 33910 40723
rect 33962 40751 33968 40763
rect 34114 40751 34142 40862
rect 48304 40859 48310 40871
rect 48362 40859 48368 40911
rect 33962 40723 34142 40751
rect 33962 40711 33968 40723
rect 1152 40652 58848 40674
rect 1152 40600 19654 40652
rect 19706 40600 19718 40652
rect 19770 40600 19782 40652
rect 19834 40600 19846 40652
rect 19898 40600 50374 40652
rect 50426 40600 50438 40652
rect 50490 40600 50502 40652
rect 50554 40600 50566 40652
rect 50618 40600 58848 40652
rect 1152 40578 58848 40600
rect 44947 40532 45005 40538
rect 44947 40498 44959 40532
rect 44993 40529 45005 40532
rect 46864 40529 46870 40541
rect 44993 40501 46870 40529
rect 44993 40498 45005 40501
rect 44947 40492 45005 40498
rect 46864 40489 46870 40501
rect 46922 40489 46928 40541
rect 25072 40045 25078 40097
rect 25130 40085 25136 40097
rect 26611 40088 26669 40094
rect 26611 40085 26623 40088
rect 25130 40057 26623 40085
rect 25130 40045 25136 40057
rect 26611 40054 26623 40057
rect 26657 40085 26669 40088
rect 26803 40088 26861 40094
rect 26803 40085 26815 40088
rect 26657 40057 26815 40085
rect 26657 40054 26669 40057
rect 26611 40048 26669 40054
rect 26803 40054 26815 40057
rect 26849 40054 26861 40088
rect 26803 40048 26861 40054
rect 57232 40045 57238 40097
rect 57290 40085 57296 40097
rect 57331 40088 57389 40094
rect 57331 40085 57343 40088
rect 57290 40057 57343 40085
rect 57290 40045 57296 40057
rect 57331 40054 57343 40057
rect 57377 40085 57389 40088
rect 57523 40088 57581 40094
rect 57523 40085 57535 40088
rect 57377 40057 57535 40085
rect 57377 40054 57389 40057
rect 57331 40048 57389 40054
rect 57523 40054 57535 40057
rect 57569 40054 57581 40088
rect 57523 40048 57581 40054
rect 1152 39986 58848 40008
rect 1152 39934 4294 39986
rect 4346 39934 4358 39986
rect 4410 39934 4422 39986
rect 4474 39934 4486 39986
rect 4538 39934 35014 39986
rect 35066 39934 35078 39986
rect 35130 39934 35142 39986
rect 35194 39934 35206 39986
rect 35258 39934 58848 39986
rect 1152 39912 58848 39934
rect 23728 39823 23734 39875
rect 23786 39863 23792 39875
rect 57232 39863 57238 39875
rect 23786 39835 57238 39863
rect 23786 39823 23792 39835
rect 57232 39823 57238 39835
rect 57290 39823 57296 39875
rect 57811 39570 57869 39576
rect 57811 39536 57823 39570
rect 57857 39536 57869 39570
rect 57811 39530 57869 39536
rect 57715 39422 57773 39428
rect 57715 39388 57727 39422
rect 57761 39419 57773 39422
rect 57826 39419 57854 39530
rect 57904 39419 57910 39431
rect 57761 39391 57910 39419
rect 57761 39388 57773 39391
rect 57715 39382 57773 39388
rect 57904 39379 57910 39391
rect 57962 39379 57968 39431
rect 1152 39320 58848 39342
rect 1152 39268 19654 39320
rect 19706 39268 19718 39320
rect 19770 39268 19782 39320
rect 19834 39268 19846 39320
rect 19898 39268 50374 39320
rect 50426 39268 50438 39320
rect 50490 39268 50502 39320
rect 50554 39268 50566 39320
rect 50618 39268 58848 39320
rect 1152 39246 58848 39268
rect 30739 39200 30797 39206
rect 30739 39166 30751 39200
rect 30785 39197 30797 39200
rect 32752 39197 32758 39209
rect 30785 39169 32758 39197
rect 30785 39166 30797 39169
rect 30739 39160 30797 39166
rect 32752 39157 32758 39169
rect 32810 39157 32816 39209
rect 1840 38861 1846 38913
rect 1898 38901 1904 38913
rect 26611 38904 26669 38910
rect 26611 38901 26623 38904
rect 1898 38873 26623 38901
rect 1898 38861 1904 38873
rect 26611 38870 26623 38873
rect 26657 38870 26669 38904
rect 26611 38864 26669 38870
rect 10387 38756 10445 38762
rect 10387 38722 10399 38756
rect 10433 38753 10445 38756
rect 10672 38753 10678 38765
rect 10433 38725 10678 38753
rect 10433 38722 10445 38725
rect 10387 38716 10445 38722
rect 10672 38713 10678 38725
rect 10730 38713 10736 38765
rect 24115 38756 24173 38762
rect 24115 38722 24127 38756
rect 24161 38753 24173 38756
rect 24403 38756 24461 38762
rect 24403 38753 24415 38756
rect 24161 38725 24415 38753
rect 24161 38722 24173 38725
rect 24115 38716 24173 38722
rect 24403 38722 24415 38725
rect 24449 38753 24461 38756
rect 30544 38753 30550 38765
rect 24449 38725 30550 38753
rect 24449 38722 24461 38725
rect 24403 38716 24461 38722
rect 30544 38713 30550 38725
rect 30602 38713 30608 38765
rect 31315 38756 31373 38762
rect 31315 38722 31327 38756
rect 31361 38753 31373 38756
rect 31504 38753 31510 38765
rect 31361 38725 31510 38753
rect 31361 38722 31373 38725
rect 31315 38716 31373 38722
rect 31504 38713 31510 38725
rect 31562 38753 31568 38765
rect 31603 38756 31661 38762
rect 31603 38753 31615 38756
rect 31562 38725 31615 38753
rect 31562 38713 31568 38725
rect 31603 38722 31615 38725
rect 31649 38722 31661 38756
rect 31603 38716 31661 38722
rect 57616 38713 57622 38765
rect 57674 38753 57680 38765
rect 57811 38756 57869 38762
rect 57811 38753 57823 38756
rect 57674 38725 57823 38753
rect 57674 38713 57680 38725
rect 57811 38722 57823 38725
rect 57857 38722 57869 38756
rect 57811 38716 57869 38722
rect 1152 38654 58848 38676
rect 1152 38602 4294 38654
rect 4346 38602 4358 38654
rect 4410 38602 4422 38654
rect 4474 38602 4486 38654
rect 4538 38602 35014 38654
rect 35066 38602 35078 38654
rect 35130 38602 35142 38654
rect 35194 38602 35206 38654
rect 35258 38602 58848 38654
rect 1152 38580 58848 38602
rect 27346 38281 37454 38309
rect 12688 38195 12694 38247
rect 12746 38235 12752 38247
rect 27346 38235 27374 38281
rect 12746 38207 27374 38235
rect 34099 38238 34157 38244
rect 12746 38195 12752 38207
rect 34099 38204 34111 38238
rect 34145 38235 34157 38238
rect 34387 38238 34445 38244
rect 34387 38235 34399 38238
rect 34145 38207 34399 38235
rect 34145 38204 34157 38207
rect 34099 38198 34157 38204
rect 34387 38204 34399 38207
rect 34433 38204 34445 38238
rect 37426 38235 37454 38281
rect 54643 38238 54701 38244
rect 54643 38235 54655 38238
rect 37426 38207 54655 38235
rect 34387 38198 34445 38204
rect 54643 38204 54655 38207
rect 54689 38204 54701 38238
rect 54643 38198 54701 38204
rect 55411 38238 55469 38244
rect 55411 38204 55423 38238
rect 55457 38204 55469 38238
rect 55411 38198 55469 38204
rect 13840 38121 13846 38173
rect 13898 38161 13904 38173
rect 55219 38164 55277 38170
rect 55219 38161 55231 38164
rect 13898 38133 55231 38161
rect 13898 38121 13904 38133
rect 55219 38130 55231 38133
rect 55265 38161 55277 38164
rect 55426 38161 55454 38198
rect 55265 38133 55454 38161
rect 55265 38130 55277 38133
rect 55219 38124 55277 38130
rect 32656 38047 32662 38099
rect 32714 38087 32720 38099
rect 34099 38090 34157 38096
rect 34099 38087 34111 38090
rect 32714 38059 34111 38087
rect 32714 38047 32720 38059
rect 34099 38056 34111 38059
rect 34145 38087 34157 38090
rect 34195 38090 34253 38096
rect 34195 38087 34207 38090
rect 34145 38059 34207 38087
rect 34145 38056 34157 38059
rect 34099 38050 34157 38056
rect 34195 38056 34207 38059
rect 34241 38056 34253 38090
rect 34195 38050 34253 38056
rect 1152 37988 58848 38010
rect 1152 37936 19654 37988
rect 19706 37936 19718 37988
rect 19770 37936 19782 37988
rect 19834 37936 19846 37988
rect 19898 37936 50374 37988
rect 50426 37936 50438 37988
rect 50490 37936 50502 37988
rect 50554 37936 50566 37988
rect 50618 37936 58848 37988
rect 1152 37914 58848 37936
rect 5008 37421 5014 37433
rect 4969 37393 5014 37421
rect 5008 37381 5014 37393
rect 5066 37381 5072 37433
rect 5779 37424 5837 37430
rect 5779 37390 5791 37424
rect 5825 37421 5837 37424
rect 6064 37421 6070 37433
rect 5825 37393 6070 37421
rect 5825 37390 5837 37393
rect 5779 37384 5837 37390
rect 6064 37381 6070 37393
rect 6122 37381 6128 37433
rect 30928 37381 30934 37433
rect 30986 37421 30992 37433
rect 43315 37424 43373 37430
rect 43315 37421 43327 37424
rect 30986 37393 43327 37421
rect 30986 37381 30992 37393
rect 43315 37390 43327 37393
rect 43361 37390 43373 37424
rect 43315 37384 43373 37390
rect 1152 37322 58848 37344
rect 1152 37270 4294 37322
rect 4346 37270 4358 37322
rect 4410 37270 4422 37322
rect 4474 37270 4486 37322
rect 4538 37270 35014 37322
rect 35066 37270 35078 37322
rect 35130 37270 35142 37322
rect 35194 37270 35206 37322
rect 35258 37270 58848 37322
rect 1152 37248 58848 37270
rect 5008 37159 5014 37211
rect 5066 37199 5072 37211
rect 52912 37199 52918 37211
rect 5066 37171 52918 37199
rect 5066 37159 5072 37171
rect 52912 37159 52918 37171
rect 52970 37159 52976 37211
rect 14611 36906 14669 36912
rect 14611 36872 14623 36906
rect 14657 36903 14669 36906
rect 14896 36903 14902 36915
rect 14657 36875 14902 36903
rect 14657 36872 14669 36875
rect 14611 36866 14669 36872
rect 14896 36863 14902 36875
rect 14954 36863 14960 36915
rect 24019 36906 24077 36912
rect 24019 36903 24031 36906
rect 23842 36875 24031 36903
rect 18448 36715 18454 36767
rect 18506 36755 18512 36767
rect 23842 36764 23870 36875
rect 24019 36872 24031 36875
rect 24065 36872 24077 36906
rect 24019 36866 24077 36872
rect 23827 36758 23885 36764
rect 23827 36755 23839 36758
rect 18506 36727 23839 36755
rect 18506 36715 18512 36727
rect 23827 36724 23839 36727
rect 23873 36724 23885 36758
rect 23827 36718 23885 36724
rect 1152 36656 58848 36678
rect 1152 36604 19654 36656
rect 19706 36604 19718 36656
rect 19770 36604 19782 36656
rect 19834 36604 19846 36656
rect 19898 36604 50374 36656
rect 50426 36604 50438 36656
rect 50490 36604 50502 36656
rect 50554 36604 50566 36656
rect 50618 36604 58848 36656
rect 1152 36582 58848 36604
rect 14896 36493 14902 36545
rect 14954 36533 14960 36545
rect 32368 36533 32374 36545
rect 14954 36505 32374 36533
rect 14954 36493 14960 36505
rect 32368 36493 32374 36505
rect 32426 36493 32432 36545
rect 9811 36240 9869 36246
rect 9811 36206 9823 36240
rect 9857 36237 9869 36240
rect 19504 36237 19510 36249
rect 9857 36209 19510 36237
rect 9857 36206 9869 36209
rect 9811 36200 9869 36206
rect 19504 36197 19510 36209
rect 19562 36197 19568 36249
rect 16915 36166 16973 36172
rect 16915 36163 16927 36166
rect 7186 36135 16927 36163
rect 2896 36049 2902 36101
rect 2954 36089 2960 36101
rect 7186 36089 7214 36135
rect 16915 36132 16927 36135
rect 16961 36163 16973 36166
rect 17107 36166 17165 36172
rect 17107 36163 17119 36166
rect 16961 36135 17119 36163
rect 16961 36132 16973 36135
rect 16915 36126 16973 36132
rect 17107 36132 17119 36135
rect 17153 36132 17165 36166
rect 18640 36163 18646 36175
rect 17107 36126 17165 36132
rect 17266 36135 18646 36163
rect 2954 36061 7214 36089
rect 2954 36049 2960 36061
rect 12496 36049 12502 36101
rect 12554 36089 12560 36101
rect 17266 36089 17294 36135
rect 18640 36123 18646 36135
rect 18698 36123 18704 36175
rect 12554 36061 17294 36089
rect 12554 36049 12560 36061
rect 17872 36049 17878 36101
rect 17930 36089 17936 36101
rect 20659 36092 20717 36098
rect 20659 36089 20671 36092
rect 17930 36061 20671 36089
rect 17930 36049 17936 36061
rect 20659 36058 20671 36061
rect 20705 36089 20717 36092
rect 20851 36092 20909 36098
rect 20851 36089 20863 36092
rect 20705 36061 20863 36089
rect 20705 36058 20717 36061
rect 20659 36052 20717 36058
rect 20851 36058 20863 36061
rect 20897 36058 20909 36092
rect 44368 36089 44374 36101
rect 44329 36061 44374 36089
rect 20851 36052 20909 36058
rect 44368 36049 44374 36061
rect 44426 36089 44432 36101
rect 44563 36092 44621 36098
rect 44563 36089 44575 36092
rect 44426 36061 44575 36089
rect 44426 36049 44432 36061
rect 44563 36058 44575 36061
rect 44609 36058 44621 36092
rect 44563 36052 44621 36058
rect 1152 35990 58848 36012
rect 1152 35938 4294 35990
rect 4346 35938 4358 35990
rect 4410 35938 4422 35990
rect 4474 35938 4486 35990
rect 4538 35938 35014 35990
rect 35066 35938 35078 35990
rect 35130 35938 35142 35990
rect 35194 35938 35206 35990
rect 35258 35938 58848 35990
rect 1152 35916 58848 35938
rect 3280 35531 3286 35583
rect 3338 35571 3344 35583
rect 10675 35574 10733 35580
rect 10675 35571 10687 35574
rect 3338 35543 10687 35571
rect 3338 35531 3344 35543
rect 10675 35540 10687 35543
rect 10721 35571 10733 35574
rect 10867 35574 10925 35580
rect 10867 35571 10879 35574
rect 10721 35543 10879 35571
rect 10721 35540 10733 35543
rect 10675 35534 10733 35540
rect 10867 35540 10879 35543
rect 10913 35540 10925 35574
rect 10867 35534 10925 35540
rect 20371 35574 20429 35580
rect 20371 35540 20383 35574
rect 20417 35571 20429 35574
rect 20656 35571 20662 35583
rect 20417 35543 20662 35571
rect 20417 35540 20429 35543
rect 20371 35534 20429 35540
rect 20656 35531 20662 35543
rect 20714 35531 20720 35583
rect 21043 35574 21101 35580
rect 21043 35540 21055 35574
rect 21089 35571 21101 35574
rect 21331 35574 21389 35580
rect 21331 35571 21343 35574
rect 21089 35543 21343 35571
rect 21089 35540 21101 35543
rect 21043 35534 21101 35540
rect 21331 35540 21343 35543
rect 21377 35571 21389 35574
rect 21712 35571 21718 35583
rect 21377 35543 21718 35571
rect 21377 35540 21389 35543
rect 21331 35534 21389 35540
rect 21712 35531 21718 35543
rect 21770 35531 21776 35583
rect 32560 35531 32566 35583
rect 32618 35571 32624 35583
rect 52627 35574 52685 35580
rect 52627 35571 52639 35574
rect 32618 35543 52639 35571
rect 32618 35531 32624 35543
rect 52627 35540 52639 35543
rect 52673 35571 52685 35574
rect 52819 35574 52877 35580
rect 52819 35571 52831 35574
rect 52673 35543 52831 35571
rect 52673 35540 52685 35543
rect 52627 35534 52685 35540
rect 52819 35540 52831 35543
rect 52865 35540 52877 35574
rect 52819 35534 52877 35540
rect 56659 35574 56717 35580
rect 56659 35540 56671 35574
rect 56705 35540 56717 35574
rect 56659 35534 56717 35540
rect 56674 35435 56702 35534
rect 56563 35426 56621 35432
rect 56563 35392 56575 35426
rect 56609 35423 56621 35426
rect 56656 35423 56662 35435
rect 56609 35395 56662 35423
rect 56609 35392 56621 35395
rect 56563 35386 56621 35392
rect 56656 35383 56662 35395
rect 56714 35383 56720 35435
rect 1152 35324 58848 35346
rect 1152 35272 19654 35324
rect 19706 35272 19718 35324
rect 19770 35272 19782 35324
rect 19834 35272 19846 35324
rect 19898 35272 50374 35324
rect 50426 35272 50438 35324
rect 50490 35272 50502 35324
rect 50554 35272 50566 35324
rect 50618 35272 58848 35324
rect 1152 35250 58848 35272
rect 30931 34834 30989 34840
rect 30931 34800 30943 34834
rect 30977 34831 30989 34834
rect 40816 34831 40822 34843
rect 30977 34803 40822 34831
rect 30977 34800 30989 34803
rect 30931 34794 30989 34800
rect 40816 34791 40822 34803
rect 40874 34791 40880 34843
rect 15571 34760 15629 34766
rect 15571 34726 15583 34760
rect 15617 34757 15629 34760
rect 15859 34760 15917 34766
rect 15859 34757 15871 34760
rect 15617 34729 15871 34757
rect 15617 34726 15629 34729
rect 15571 34720 15629 34726
rect 15859 34726 15871 34729
rect 15905 34757 15917 34760
rect 26800 34757 26806 34769
rect 15905 34729 26806 34757
rect 15905 34726 15917 34729
rect 15859 34720 15917 34726
rect 26800 34717 26806 34729
rect 26858 34717 26864 34769
rect 31408 34757 31414 34769
rect 31369 34729 31414 34757
rect 31408 34717 31414 34729
rect 31466 34757 31472 34769
rect 31507 34760 31565 34766
rect 31507 34757 31519 34760
rect 31466 34729 31519 34757
rect 31466 34717 31472 34729
rect 31507 34726 31519 34729
rect 31553 34726 31565 34760
rect 31507 34720 31565 34726
rect 53107 34760 53165 34766
rect 53107 34726 53119 34760
rect 53153 34757 53165 34760
rect 53200 34757 53206 34769
rect 53153 34729 53206 34757
rect 53153 34726 53165 34729
rect 53107 34720 53165 34726
rect 53200 34717 53206 34729
rect 53258 34717 53264 34769
rect 57040 34757 57046 34769
rect 57001 34729 57046 34757
rect 57040 34717 57046 34729
rect 57098 34757 57104 34769
rect 57235 34760 57293 34766
rect 57235 34757 57247 34760
rect 57098 34729 57247 34757
rect 57098 34717 57104 34729
rect 57235 34726 57247 34729
rect 57281 34726 57293 34760
rect 57235 34720 57293 34726
rect 1152 34658 58848 34680
rect 1152 34606 4294 34658
rect 4346 34606 4358 34658
rect 4410 34606 4422 34658
rect 4474 34606 4486 34658
rect 4538 34606 35014 34658
rect 35066 34606 35078 34658
rect 35130 34606 35142 34658
rect 35194 34606 35206 34658
rect 35258 34606 58848 34658
rect 1152 34584 58848 34606
rect 24400 34273 24406 34325
rect 24458 34313 24464 34325
rect 24458 34285 37454 34313
rect 24458 34273 24464 34285
rect 28243 34242 28301 34248
rect 28243 34208 28255 34242
rect 28289 34208 28301 34242
rect 37426 34239 37454 34285
rect 58003 34242 58061 34248
rect 58003 34239 58015 34242
rect 37426 34211 58015 34239
rect 28243 34202 28301 34208
rect 58003 34208 58015 34211
rect 58049 34208 58061 34242
rect 58003 34202 58061 34208
rect 28258 34165 28286 34202
rect 53392 34165 53398 34177
rect 28258 34137 53398 34165
rect 53392 34125 53398 34137
rect 53450 34125 53456 34177
rect 1152 33992 58848 34014
rect 1152 33940 19654 33992
rect 19706 33940 19718 33992
rect 19770 33940 19782 33992
rect 19834 33940 19846 33992
rect 19898 33940 50374 33992
rect 50426 33940 50438 33992
rect 50490 33940 50502 33992
rect 50554 33940 50566 33992
rect 50618 33940 58848 33992
rect 1152 33918 58848 33940
rect 21712 33829 21718 33881
rect 21770 33869 21776 33881
rect 51472 33869 51478 33881
rect 21770 33841 51478 33869
rect 21770 33829 21776 33841
rect 51472 33829 51478 33841
rect 51530 33829 51536 33881
rect 26707 33502 26765 33508
rect 26707 33468 26719 33502
rect 26753 33499 26765 33502
rect 56272 33499 56278 33511
rect 26753 33471 56278 33499
rect 26753 33468 26765 33471
rect 26707 33462 26765 33468
rect 56272 33459 56278 33471
rect 56330 33459 56336 33511
rect 10576 33385 10582 33437
rect 10634 33425 10640 33437
rect 16819 33428 16877 33434
rect 16819 33425 16831 33428
rect 10634 33397 16831 33425
rect 10634 33385 10640 33397
rect 16819 33394 16831 33397
rect 16865 33394 16877 33428
rect 16819 33388 16877 33394
rect 35923 33428 35981 33434
rect 35923 33394 35935 33428
rect 35969 33425 35981 33428
rect 36211 33428 36269 33434
rect 36211 33425 36223 33428
rect 35969 33397 36223 33425
rect 35969 33394 35981 33397
rect 35923 33388 35981 33394
rect 36211 33394 36223 33397
rect 36257 33425 36269 33428
rect 38128 33425 38134 33437
rect 36257 33397 38134 33425
rect 36257 33394 36269 33397
rect 36211 33388 36269 33394
rect 38128 33385 38134 33397
rect 38186 33385 38192 33437
rect 1152 33326 58848 33348
rect 1152 33274 4294 33326
rect 4346 33274 4358 33326
rect 4410 33274 4422 33326
rect 4474 33274 4486 33326
rect 4538 33274 35014 33326
rect 35066 33274 35078 33326
rect 35130 33274 35142 33326
rect 35194 33274 35206 33326
rect 35258 33274 58848 33326
rect 1152 33252 58848 33274
rect 10384 32719 10390 32771
rect 10442 32759 10448 32771
rect 39571 32762 39629 32768
rect 39571 32759 39583 32762
rect 10442 32731 39583 32759
rect 10442 32719 10448 32731
rect 39571 32728 39583 32731
rect 39617 32728 39629 32762
rect 39571 32722 39629 32728
rect 1152 32660 58848 32682
rect 1152 32608 19654 32660
rect 19706 32608 19718 32660
rect 19770 32608 19782 32660
rect 19834 32608 19846 32660
rect 19898 32608 50374 32660
rect 50426 32608 50438 32660
rect 50490 32608 50502 32660
rect 50554 32608 50566 32660
rect 50618 32608 58848 32660
rect 1152 32586 58848 32608
rect 32563 32244 32621 32250
rect 32563 32241 32575 32244
rect 7186 32213 32575 32241
rect 5875 32096 5933 32102
rect 5875 32062 5887 32096
rect 5921 32093 5933 32096
rect 7186 32093 7214 32213
rect 32563 32210 32575 32213
rect 32609 32210 32621 32244
rect 32563 32204 32621 32210
rect 26227 32170 26285 32176
rect 26227 32136 26239 32170
rect 26273 32167 26285 32170
rect 51952 32167 51958 32179
rect 26273 32139 51958 32167
rect 26273 32136 26285 32139
rect 26227 32130 26285 32136
rect 51952 32127 51958 32139
rect 52010 32127 52016 32179
rect 5921 32065 7214 32093
rect 21619 32096 21677 32102
rect 5921 32062 5933 32065
rect 5875 32056 5933 32062
rect 21619 32062 21631 32096
rect 21665 32093 21677 32096
rect 24496 32093 24502 32105
rect 21665 32065 24502 32093
rect 21665 32062 21677 32065
rect 21619 32056 21677 32062
rect 24496 32053 24502 32065
rect 24554 32053 24560 32105
rect 27376 32053 27382 32105
rect 27434 32093 27440 32105
rect 32563 32096 32621 32102
rect 27434 32065 27479 32093
rect 27434 32053 27440 32065
rect 32563 32062 32575 32096
rect 32609 32093 32621 32096
rect 53296 32093 53302 32105
rect 32609 32065 53302 32093
rect 32609 32062 32621 32065
rect 32563 32056 32621 32062
rect 53296 32053 53302 32065
rect 53354 32053 53360 32105
rect 1152 31994 58848 32016
rect 1152 31942 4294 31994
rect 4346 31942 4358 31994
rect 4410 31942 4422 31994
rect 4474 31942 4486 31994
rect 4538 31942 35014 31994
rect 35066 31942 35078 31994
rect 35130 31942 35142 31994
rect 35194 31942 35206 31994
rect 35258 31942 58848 31994
rect 1152 31920 58848 31942
rect 27376 31831 27382 31883
rect 27434 31871 27440 31883
rect 50128 31871 50134 31883
rect 27434 31843 50134 31871
rect 27434 31831 27440 31843
rect 50128 31831 50134 31843
rect 50186 31831 50192 31883
rect 24496 31757 24502 31809
rect 24554 31797 24560 31809
rect 35440 31797 35446 31809
rect 24554 31769 35446 31797
rect 24554 31757 24560 31769
rect 35440 31757 35446 31769
rect 35498 31757 35504 31809
rect 35344 31683 35350 31735
rect 35402 31723 35408 31735
rect 52819 31726 52877 31732
rect 52819 31723 52831 31726
rect 35402 31695 52831 31723
rect 35402 31683 35408 31695
rect 52819 31692 52831 31695
rect 52865 31692 52877 31726
rect 52819 31686 52877 31692
rect 6448 31609 6454 31661
rect 6506 31649 6512 31661
rect 8080 31649 8086 31661
rect 6506 31621 8086 31649
rect 6506 31609 6512 31621
rect 8080 31609 8086 31621
rect 8138 31609 8144 31661
rect 1152 31328 58848 31350
rect 1152 31276 19654 31328
rect 19706 31276 19718 31328
rect 19770 31276 19782 31328
rect 19834 31276 19846 31328
rect 19898 31276 50374 31328
rect 50426 31276 50438 31328
rect 50490 31276 50502 31328
rect 50554 31276 50566 31328
rect 50618 31276 58848 31328
rect 1152 31254 58848 31276
rect 20563 30912 20621 30918
rect 20563 30878 20575 30912
rect 20609 30909 20621 30912
rect 34000 30909 34006 30921
rect 20609 30881 34006 30909
rect 20609 30878 20621 30881
rect 20563 30872 20621 30878
rect 34000 30869 34006 30881
rect 34058 30869 34064 30921
rect 53395 30838 53453 30844
rect 53395 30835 53407 30838
rect 47506 30807 53407 30835
rect 6931 30764 6989 30770
rect 6931 30730 6943 30764
rect 6977 30761 6989 30764
rect 12592 30761 12598 30773
rect 6977 30733 12598 30761
rect 6977 30730 6989 30733
rect 6931 30724 6989 30730
rect 12592 30721 12598 30733
rect 12650 30721 12656 30773
rect 19024 30761 19030 30773
rect 18985 30733 19030 30761
rect 19024 30721 19030 30733
rect 19082 30721 19088 30773
rect 24016 30721 24022 30773
rect 24074 30761 24080 30773
rect 47506 30761 47534 30807
rect 53395 30804 53407 30807
rect 53441 30804 53453 30838
rect 53395 30798 53453 30804
rect 24074 30733 47534 30761
rect 24074 30721 24080 30733
rect 51856 30721 51862 30773
rect 51914 30761 51920 30773
rect 52051 30764 52109 30770
rect 52051 30761 52063 30764
rect 51914 30733 52063 30761
rect 51914 30721 51920 30733
rect 52051 30730 52063 30733
rect 52097 30730 52109 30764
rect 55312 30761 55318 30773
rect 55273 30733 55318 30761
rect 52051 30724 52109 30730
rect 55312 30721 55318 30733
rect 55370 30721 55376 30773
rect 1152 30662 58848 30684
rect 1152 30610 4294 30662
rect 4346 30610 4358 30662
rect 4410 30610 4422 30662
rect 4474 30610 4486 30662
rect 4538 30610 35014 30662
rect 35066 30610 35078 30662
rect 35130 30610 35142 30662
rect 35194 30610 35206 30662
rect 35258 30610 58848 30662
rect 1152 30588 58848 30610
rect 29488 30499 29494 30551
rect 29546 30539 29552 30551
rect 55312 30539 55318 30551
rect 29546 30511 55318 30539
rect 29546 30499 29552 30511
rect 55312 30499 55318 30511
rect 55370 30499 55376 30551
rect 19024 30425 19030 30477
rect 19082 30465 19088 30477
rect 38224 30465 38230 30477
rect 19082 30437 38230 30465
rect 19082 30425 19088 30437
rect 38224 30425 38230 30437
rect 38282 30425 38288 30477
rect 38899 30394 38957 30400
rect 38899 30360 38911 30394
rect 38945 30391 38957 30394
rect 52144 30391 52150 30403
rect 38945 30363 52150 30391
rect 38945 30360 38957 30363
rect 38899 30354 38957 30360
rect 52144 30351 52150 30363
rect 52202 30351 52208 30403
rect 4339 30320 4397 30326
rect 4339 30286 4351 30320
rect 4385 30317 4397 30320
rect 4627 30320 4685 30326
rect 4627 30317 4639 30320
rect 4385 30289 4639 30317
rect 4385 30286 4397 30289
rect 4339 30280 4397 30286
rect 4627 30286 4639 30289
rect 4673 30317 4685 30320
rect 51568 30317 51574 30329
rect 4673 30289 51574 30317
rect 4673 30286 4685 30289
rect 4627 30280 4685 30286
rect 51568 30277 51574 30289
rect 51626 30277 51632 30329
rect 1152 29996 58848 30018
rect 1152 29944 19654 29996
rect 19706 29944 19718 29996
rect 19770 29944 19782 29996
rect 19834 29944 19846 29996
rect 19898 29944 50374 29996
rect 50426 29944 50438 29996
rect 50490 29944 50502 29996
rect 50554 29944 50566 29996
rect 50618 29944 58848 29996
rect 1152 29922 58848 29944
rect 36403 29506 36461 29512
rect 36403 29472 36415 29506
rect 36449 29503 36461 29506
rect 36449 29475 37454 29503
rect 36449 29472 36461 29475
rect 36403 29466 36461 29472
rect 6256 29429 6262 29441
rect 6217 29401 6262 29429
rect 6256 29389 6262 29401
rect 6314 29389 6320 29441
rect 37072 29429 37078 29441
rect 37033 29401 37078 29429
rect 37072 29389 37078 29401
rect 37130 29389 37136 29441
rect 37426 29429 37454 29475
rect 49072 29429 49078 29441
rect 37426 29401 49078 29429
rect 49072 29389 49078 29401
rect 49130 29389 49136 29441
rect 1152 29330 58848 29352
rect 1152 29278 4294 29330
rect 4346 29278 4358 29330
rect 4410 29278 4422 29330
rect 4474 29278 4486 29330
rect 4538 29278 35014 29330
rect 35066 29278 35078 29330
rect 35130 29278 35142 29330
rect 35194 29278 35206 29330
rect 35258 29278 58848 29330
rect 1152 29256 58848 29278
rect 37072 29167 37078 29219
rect 37130 29207 37136 29219
rect 49360 29207 49366 29219
rect 37130 29179 49366 29207
rect 37130 29167 37136 29179
rect 49360 29167 49366 29179
rect 49418 29167 49424 29219
rect 13936 28871 13942 28923
rect 13994 28911 14000 28923
rect 18451 28914 18509 28920
rect 18451 28911 18463 28914
rect 13994 28883 18463 28911
rect 13994 28871 14000 28883
rect 18451 28880 18463 28883
rect 18497 28880 18509 28914
rect 18451 28874 18509 28880
rect 37555 28914 37613 28920
rect 37555 28880 37567 28914
rect 37601 28911 37613 28914
rect 44080 28911 44086 28923
rect 37601 28883 44086 28911
rect 37601 28880 37613 28883
rect 37555 28874 37613 28880
rect 44080 28871 44086 28883
rect 44138 28871 44144 28923
rect 1152 28664 58848 28686
rect 1152 28612 19654 28664
rect 19706 28612 19718 28664
rect 19770 28612 19782 28664
rect 19834 28612 19846 28664
rect 19898 28612 50374 28664
rect 50426 28612 50438 28664
rect 50490 28612 50502 28664
rect 50554 28612 50566 28664
rect 50618 28612 58848 28664
rect 1152 28590 58848 28612
rect 2992 28057 2998 28109
rect 3050 28097 3056 28109
rect 10963 28100 11021 28106
rect 10963 28097 10975 28100
rect 3050 28069 10975 28097
rect 3050 28057 3056 28069
rect 10963 28066 10975 28069
rect 11009 28097 11021 28100
rect 11155 28100 11213 28106
rect 11155 28097 11167 28100
rect 11009 28069 11167 28097
rect 11009 28066 11021 28069
rect 10963 28060 11021 28066
rect 11155 28066 11167 28069
rect 11201 28066 11213 28100
rect 11155 28060 11213 28066
rect 36211 28100 36269 28106
rect 36211 28066 36223 28100
rect 36257 28097 36269 28100
rect 45616 28097 45622 28109
rect 36257 28069 45622 28097
rect 36257 28066 36269 28069
rect 36211 28060 36269 28066
rect 45616 28057 45622 28069
rect 45674 28057 45680 28109
rect 1152 27998 58848 28020
rect 1152 27946 4294 27998
rect 4346 27946 4358 27998
rect 4410 27946 4422 27998
rect 4474 27946 4486 27998
rect 4538 27946 35014 27998
rect 35066 27946 35078 27998
rect 35130 27946 35142 27998
rect 35194 27946 35206 27998
rect 35258 27946 58848 27998
rect 1152 27924 58848 27946
rect 24211 27878 24269 27884
rect 24211 27844 24223 27878
rect 24257 27875 24269 27878
rect 24304 27875 24310 27887
rect 24257 27847 24310 27875
rect 24257 27844 24269 27847
rect 24211 27838 24269 27844
rect 24304 27835 24310 27847
rect 24362 27835 24368 27887
rect 18259 27656 18317 27662
rect 18259 27622 18271 27656
rect 18305 27653 18317 27656
rect 35536 27653 35542 27665
rect 18305 27625 35542 27653
rect 18305 27622 18317 27625
rect 18259 27616 18317 27622
rect 35536 27613 35542 27625
rect 35594 27613 35600 27665
rect 52528 27539 52534 27591
rect 52586 27579 52592 27591
rect 56371 27582 56429 27588
rect 56371 27579 56383 27582
rect 52586 27551 56383 27579
rect 52586 27539 52592 27551
rect 56371 27548 56383 27551
rect 56417 27548 56429 27582
rect 56371 27542 56429 27548
rect 57043 27582 57101 27588
rect 57043 27548 57055 27582
rect 57089 27548 57101 27582
rect 57043 27542 57101 27548
rect 13552 27465 13558 27517
rect 13610 27505 13616 27517
rect 13610 27477 27374 27505
rect 13610 27465 13616 27477
rect 27346 27431 27374 27477
rect 42736 27465 42742 27517
rect 42794 27505 42800 27517
rect 57058 27505 57086 27542
rect 42794 27477 57086 27505
rect 42794 27465 42800 27477
rect 27955 27434 28013 27440
rect 27955 27431 27967 27434
rect 27346 27403 27967 27431
rect 27955 27400 27967 27403
rect 28001 27431 28013 27434
rect 28051 27434 28109 27440
rect 28051 27431 28063 27434
rect 28001 27403 28063 27431
rect 28001 27400 28013 27403
rect 27955 27394 28013 27400
rect 28051 27400 28063 27403
rect 28097 27400 28109 27434
rect 28051 27394 28109 27400
rect 1152 27332 58848 27354
rect 1152 27280 19654 27332
rect 19706 27280 19718 27332
rect 19770 27280 19782 27332
rect 19834 27280 19846 27332
rect 19898 27280 50374 27332
rect 50426 27280 50438 27332
rect 50490 27280 50502 27332
rect 50554 27280 50566 27332
rect 50618 27280 58848 27332
rect 1152 27258 58848 27280
rect 6352 26947 6358 26999
rect 6410 26987 6416 26999
rect 18739 26990 18797 26996
rect 18739 26987 18751 26990
rect 6410 26959 18751 26987
rect 6410 26947 6416 26959
rect 18739 26956 18751 26959
rect 18785 26987 18797 26990
rect 18931 26990 18989 26996
rect 18931 26987 18943 26990
rect 18785 26959 18943 26987
rect 18785 26956 18797 26959
rect 18739 26950 18797 26956
rect 18931 26956 18943 26959
rect 18977 26956 18989 26990
rect 18931 26950 18989 26956
rect 16816 26873 16822 26925
rect 16874 26913 16880 26925
rect 42160 26913 42166 26925
rect 16874 26885 42166 26913
rect 16874 26873 16880 26885
rect 42160 26873 42166 26885
rect 42218 26873 42224 26925
rect 6832 26799 6838 26851
rect 6890 26839 6896 26851
rect 56656 26839 56662 26851
rect 6890 26811 56662 26839
rect 6890 26799 6896 26811
rect 56656 26799 56662 26811
rect 56714 26799 56720 26851
rect 14896 26725 14902 26777
rect 14954 26765 14960 26777
rect 15091 26768 15149 26774
rect 15091 26765 15103 26768
rect 14954 26737 15103 26765
rect 14954 26725 14960 26737
rect 15091 26734 15103 26737
rect 15137 26734 15149 26768
rect 15091 26728 15149 26734
rect 16048 26725 16054 26777
rect 16106 26765 16112 26777
rect 16627 26768 16685 26774
rect 16627 26765 16639 26768
rect 16106 26737 16639 26765
rect 16106 26725 16112 26737
rect 16627 26734 16639 26737
rect 16673 26734 16685 26768
rect 16627 26728 16685 26734
rect 1152 26666 58848 26688
rect 1152 26614 4294 26666
rect 4346 26614 4358 26666
rect 4410 26614 4422 26666
rect 4474 26614 4486 26666
rect 4538 26614 35014 26666
rect 35066 26614 35078 26666
rect 35130 26614 35142 26666
rect 35194 26614 35206 26666
rect 35258 26614 58848 26666
rect 1152 26592 58848 26614
rect 19408 26059 19414 26111
rect 19466 26099 19472 26111
rect 23824 26099 23830 26111
rect 19466 26071 23830 26099
rect 19466 26059 19472 26071
rect 23824 26059 23830 26071
rect 23882 26059 23888 26111
rect 1152 26000 58848 26022
rect 1152 25948 19654 26000
rect 19706 25948 19718 26000
rect 19770 25948 19782 26000
rect 19834 25948 19846 26000
rect 19898 25948 50374 26000
rect 50426 25948 50438 26000
rect 50490 25948 50502 26000
rect 50554 25948 50566 26000
rect 50618 25948 58848 26000
rect 1152 25926 58848 25948
rect 56944 25393 56950 25445
rect 57002 25433 57008 25445
rect 57331 25436 57389 25442
rect 57331 25433 57343 25436
rect 57002 25405 57343 25433
rect 57002 25393 57008 25405
rect 57331 25402 57343 25405
rect 57377 25402 57389 25436
rect 57331 25396 57389 25402
rect 1152 25334 58848 25356
rect 1152 25282 4294 25334
rect 4346 25282 4358 25334
rect 4410 25282 4422 25334
rect 4474 25282 4486 25334
rect 4538 25282 35014 25334
rect 35066 25282 35078 25334
rect 35130 25282 35142 25334
rect 35194 25282 35206 25334
rect 35258 25282 58848 25334
rect 1152 25260 58848 25282
rect 16624 25171 16630 25223
rect 16682 25211 16688 25223
rect 23632 25211 23638 25223
rect 16682 25183 23638 25211
rect 16682 25171 16688 25183
rect 23632 25171 23638 25183
rect 23690 25171 23696 25223
rect 42064 25171 42070 25223
rect 42122 25211 42128 25223
rect 46771 25214 46829 25220
rect 46771 25211 46783 25214
rect 42122 25183 46783 25211
rect 42122 25171 42128 25183
rect 46771 25180 46783 25183
rect 46817 25211 46829 25214
rect 46963 25214 47021 25220
rect 46963 25211 46975 25214
rect 46817 25183 46975 25211
rect 46817 25180 46829 25183
rect 46771 25174 46829 25180
rect 46963 25180 46975 25183
rect 47009 25180 47021 25214
rect 46963 25174 47021 25180
rect 34768 24949 34774 25001
rect 34826 24989 34832 25001
rect 54259 24992 54317 24998
rect 54259 24989 54271 24992
rect 34826 24961 54271 24989
rect 34826 24949 34832 24961
rect 54259 24958 54271 24961
rect 54305 24989 54317 24992
rect 54451 24992 54509 24998
rect 54451 24989 54463 24992
rect 54305 24961 54463 24989
rect 54305 24958 54317 24961
rect 54259 24952 54317 24958
rect 54451 24958 54463 24961
rect 54497 24958 54509 24992
rect 54451 24952 54509 24958
rect 25456 24915 25462 24927
rect 25417 24887 25462 24915
rect 25456 24875 25462 24887
rect 25514 24875 25520 24927
rect 50515 24918 50573 24924
rect 50515 24884 50527 24918
rect 50561 24915 50573 24918
rect 50704 24915 50710 24927
rect 50561 24887 50710 24915
rect 50561 24884 50573 24887
rect 50515 24878 50573 24884
rect 50704 24875 50710 24887
rect 50762 24875 50768 24927
rect 55315 24918 55373 24924
rect 55315 24884 55327 24918
rect 55361 24884 55373 24918
rect 55315 24878 55373 24884
rect 32464 24801 32470 24853
rect 32522 24841 32528 24853
rect 55330 24841 55358 24878
rect 32522 24813 55358 24841
rect 32522 24801 32528 24813
rect 1152 24668 58848 24690
rect 1152 24616 19654 24668
rect 19706 24616 19718 24668
rect 19770 24616 19782 24668
rect 19834 24616 19846 24668
rect 19898 24616 50374 24668
rect 50426 24616 50438 24668
rect 50490 24616 50502 24668
rect 50554 24616 50566 24668
rect 50618 24616 58848 24668
rect 1152 24594 58848 24616
rect 3568 24283 3574 24335
rect 3626 24323 3632 24335
rect 23248 24323 23254 24335
rect 3626 24295 23254 24323
rect 3626 24283 3632 24295
rect 23248 24283 23254 24295
rect 23306 24283 23312 24335
rect 15280 24209 15286 24261
rect 15338 24249 15344 24261
rect 39088 24249 39094 24261
rect 15338 24221 39094 24249
rect 15338 24209 15344 24221
rect 39088 24209 39094 24221
rect 39146 24209 39152 24261
rect 7120 24135 7126 24187
rect 7178 24175 7184 24187
rect 31408 24175 31414 24187
rect 7178 24147 31414 24175
rect 7178 24135 7184 24147
rect 31408 24135 31414 24147
rect 31466 24135 31472 24187
rect 21424 24061 21430 24113
rect 21482 24101 21488 24113
rect 42643 24104 42701 24110
rect 42643 24101 42655 24104
rect 21482 24073 42655 24101
rect 21482 24061 21488 24073
rect 42643 24070 42655 24073
rect 42689 24101 42701 24104
rect 42835 24104 42893 24110
rect 42835 24101 42847 24104
rect 42689 24073 42847 24101
rect 42689 24070 42701 24073
rect 42643 24064 42701 24070
rect 42835 24070 42847 24073
rect 42881 24070 42893 24104
rect 42835 24064 42893 24070
rect 1152 24002 58848 24024
rect 1152 23950 4294 24002
rect 4346 23950 4358 24002
rect 4410 23950 4422 24002
rect 4474 23950 4486 24002
rect 4538 23950 35014 24002
rect 35066 23950 35078 24002
rect 35130 23950 35142 24002
rect 35194 23950 35206 24002
rect 35258 23950 58848 24002
rect 1152 23928 58848 23950
rect 17392 23839 17398 23891
rect 17450 23879 17456 23891
rect 41872 23879 41878 23891
rect 17450 23851 41878 23879
rect 17450 23839 17456 23851
rect 41872 23839 41878 23851
rect 41930 23839 41936 23891
rect 15952 23765 15958 23817
rect 16010 23805 16016 23817
rect 45424 23805 45430 23817
rect 16010 23777 45430 23805
rect 16010 23765 16016 23777
rect 45424 23765 45430 23777
rect 45482 23765 45488 23817
rect 3664 23691 3670 23743
rect 3722 23731 3728 23743
rect 53200 23731 53206 23743
rect 3722 23703 53206 23731
rect 3722 23691 3728 23703
rect 53200 23691 53206 23703
rect 53258 23691 53264 23743
rect 1152 23336 58848 23358
rect 1152 23284 19654 23336
rect 19706 23284 19718 23336
rect 19770 23284 19782 23336
rect 19834 23284 19846 23336
rect 19898 23284 50374 23336
rect 50426 23284 50438 23336
rect 50490 23284 50502 23336
rect 50554 23284 50566 23336
rect 50618 23284 58848 23336
rect 1152 23262 58848 23284
rect 8560 22877 8566 22929
rect 8618 22917 8624 22929
rect 39568 22917 39574 22929
rect 8618 22889 39574 22917
rect 8618 22877 8624 22889
rect 39568 22877 39574 22889
rect 39626 22877 39632 22929
rect 1936 22803 1942 22855
rect 1994 22843 2000 22855
rect 38803 22846 38861 22852
rect 1994 22815 37454 22843
rect 1994 22803 2000 22815
rect 13552 22769 13558 22781
rect 13513 22741 13558 22769
rect 13552 22729 13558 22741
rect 13610 22729 13616 22781
rect 17776 22769 17782 22781
rect 17737 22741 17782 22769
rect 17776 22729 17782 22741
rect 17834 22729 17840 22781
rect 26896 22769 26902 22781
rect 26857 22741 26902 22769
rect 26896 22729 26902 22741
rect 26954 22729 26960 22781
rect 30928 22769 30934 22781
rect 30889 22741 30934 22769
rect 30928 22729 30934 22741
rect 30986 22729 30992 22781
rect 37426 22769 37454 22815
rect 38803 22812 38815 22846
rect 38849 22843 38861 22846
rect 51088 22843 51094 22855
rect 38849 22815 51094 22843
rect 38849 22812 38861 22815
rect 38803 22806 38861 22812
rect 51088 22803 51094 22815
rect 51146 22803 51152 22855
rect 41107 22772 41165 22778
rect 41107 22769 41119 22772
rect 37426 22741 41119 22769
rect 41107 22738 41119 22741
rect 41153 22769 41165 22772
rect 41299 22772 41357 22778
rect 41299 22769 41311 22772
rect 41153 22741 41311 22769
rect 41153 22738 41165 22741
rect 41107 22732 41165 22738
rect 41299 22738 41311 22741
rect 41345 22738 41357 22772
rect 41299 22732 41357 22738
rect 1152 22670 58848 22692
rect 1152 22618 4294 22670
rect 4346 22618 4358 22670
rect 4410 22618 4422 22670
rect 4474 22618 4486 22670
rect 4538 22618 35014 22670
rect 35066 22618 35078 22670
rect 35130 22618 35142 22670
rect 35194 22618 35206 22670
rect 35258 22618 58848 22670
rect 1152 22596 58848 22618
rect 8848 22507 8854 22559
rect 8906 22507 8912 22559
rect 13552 22507 13558 22559
rect 13610 22547 13616 22559
rect 32752 22547 32758 22559
rect 13610 22519 32758 22547
rect 13610 22507 13616 22519
rect 32752 22507 32758 22519
rect 32810 22507 32816 22559
rect 8371 22476 8429 22482
rect 8371 22442 8383 22476
rect 8417 22473 8429 22476
rect 8560 22473 8566 22485
rect 8417 22445 8566 22473
rect 8417 22442 8429 22445
rect 8371 22436 8429 22442
rect 8560 22433 8566 22445
rect 8618 22433 8624 22485
rect 27187 22476 27245 22482
rect 27187 22442 27199 22476
rect 27233 22473 27245 22476
rect 36880 22473 36886 22485
rect 27233 22445 36886 22473
rect 27233 22442 27245 22445
rect 27187 22436 27245 22442
rect 36880 22433 36886 22445
rect 36938 22433 36944 22485
rect 16528 22359 16534 22411
rect 16586 22399 16592 22411
rect 40240 22399 40246 22411
rect 16586 22371 40246 22399
rect 16586 22359 16592 22371
rect 40240 22359 40246 22371
rect 40298 22359 40304 22411
rect 19504 22285 19510 22337
rect 19562 22325 19568 22337
rect 20944 22325 20950 22337
rect 19562 22297 20950 22325
rect 19562 22285 19568 22297
rect 20944 22285 20950 22297
rect 21002 22285 21008 22337
rect 15571 22254 15629 22260
rect 15571 22220 15583 22254
rect 15617 22251 15629 22254
rect 26803 22254 26861 22260
rect 15617 22223 17294 22251
rect 15617 22220 15629 22223
rect 15571 22214 15629 22220
rect 8083 22180 8141 22186
rect 8083 22146 8095 22180
rect 8129 22146 8141 22180
rect 17266 22177 17294 22223
rect 26803 22220 26815 22254
rect 26849 22251 26861 22254
rect 27091 22254 27149 22260
rect 27091 22251 27103 22254
rect 26849 22223 27103 22251
rect 26849 22220 26861 22223
rect 26803 22214 26861 22220
rect 27091 22220 27103 22223
rect 27137 22251 27149 22254
rect 27187 22254 27245 22260
rect 27187 22251 27199 22254
rect 27137 22223 27199 22251
rect 27137 22220 27149 22223
rect 27091 22214 27149 22220
rect 27187 22220 27199 22223
rect 27233 22220 27245 22254
rect 27187 22214 27245 22220
rect 35632 22177 35638 22189
rect 17266 22149 35638 22177
rect 8083 22140 8141 22146
rect 35632 22137 35638 22149
rect 35690 22137 35696 22189
rect 8752 22063 8758 22115
rect 8810 22063 8816 22115
rect 1152 22004 58848 22026
rect 1152 21952 19654 22004
rect 19706 21952 19718 22004
rect 19770 21952 19782 22004
rect 19834 21952 19846 22004
rect 19898 21952 50374 22004
rect 50426 21952 50438 22004
rect 50490 21952 50502 22004
rect 50554 21952 50566 22004
rect 50618 21952 58848 22004
rect 1152 21930 58848 21952
rect 3568 21841 3574 21893
rect 3626 21881 3632 21893
rect 26896 21881 26902 21893
rect 3626 21853 26902 21881
rect 3626 21841 3632 21853
rect 26896 21841 26902 21853
rect 26954 21841 26960 21893
rect 8752 21545 8758 21597
rect 8810 21585 8816 21597
rect 58096 21585 58102 21597
rect 8810 21557 58102 21585
rect 8810 21545 8816 21557
rect 58096 21545 58102 21557
rect 58154 21545 58160 21597
rect 8368 21471 8374 21523
rect 8426 21511 8432 21523
rect 55504 21511 55510 21523
rect 8426 21483 55510 21511
rect 8426 21471 8432 21483
rect 55504 21471 55510 21483
rect 55562 21471 55568 21523
rect 7984 21397 7990 21449
rect 8042 21437 8048 21449
rect 53872 21437 53878 21449
rect 8042 21409 53878 21437
rect 8042 21397 8048 21409
rect 53872 21397 53878 21409
rect 53930 21397 53936 21449
rect 1152 21338 58848 21360
rect 1152 21286 4294 21338
rect 4346 21286 4358 21338
rect 4410 21286 4422 21338
rect 4474 21286 4486 21338
rect 4538 21286 35014 21338
rect 35066 21286 35078 21338
rect 35130 21286 35142 21338
rect 35194 21286 35206 21338
rect 35258 21286 58848 21338
rect 1152 21264 58848 21286
rect 7603 21218 7661 21224
rect 7603 21184 7615 21218
rect 7649 21215 7661 21218
rect 7649 21187 8270 21215
rect 7649 21184 7661 21187
rect 7603 21178 7661 21184
rect 8242 21141 8270 21187
rect 8752 21141 8758 21153
rect 8242 21113 8758 21141
rect 8752 21101 8758 21113
rect 8810 21101 8816 21153
rect 8368 21067 8374 21079
rect 8256 21039 8374 21067
rect 8368 21027 8374 21039
rect 8426 21027 8432 21079
rect 7942 21005 7994 21011
rect 7942 20947 7994 20953
rect 21616 20879 21622 20931
rect 21674 20919 21680 20931
rect 33523 20922 33581 20928
rect 21674 20891 27374 20919
rect 21674 20879 21680 20891
rect 27346 20845 27374 20891
rect 33523 20888 33535 20922
rect 33569 20919 33581 20922
rect 34387 20922 34445 20928
rect 34387 20919 34399 20922
rect 33569 20891 34399 20919
rect 33569 20888 33581 20891
rect 33523 20882 33581 20888
rect 34387 20888 34399 20891
rect 34433 20888 34445 20922
rect 50707 20922 50765 20928
rect 50707 20919 50719 20922
rect 34387 20882 34445 20888
rect 37426 20891 50719 20919
rect 37426 20845 37454 20891
rect 50707 20888 50719 20891
rect 50753 20919 50765 20922
rect 50899 20922 50957 20928
rect 50899 20919 50911 20922
rect 50753 20891 50911 20919
rect 50753 20888 50765 20891
rect 50707 20882 50765 20888
rect 50899 20888 50911 20891
rect 50945 20888 50957 20922
rect 50899 20882 50957 20888
rect 27346 20817 37454 20845
rect 34387 20774 34445 20780
rect 34387 20740 34399 20774
rect 34433 20771 34445 20774
rect 44656 20771 44662 20783
rect 34433 20743 44662 20771
rect 34433 20740 34445 20743
rect 34387 20734 34445 20740
rect 44656 20731 44662 20743
rect 44714 20731 44720 20783
rect 1152 20672 58848 20694
rect 1152 20620 19654 20672
rect 19706 20620 19718 20672
rect 19770 20620 19782 20672
rect 19834 20620 19846 20672
rect 19898 20620 50374 20672
rect 50426 20620 50438 20672
rect 50490 20620 50502 20672
rect 50554 20620 50566 20672
rect 50618 20620 58848 20672
rect 1152 20598 58848 20620
rect 20848 20509 20854 20561
rect 20906 20549 20912 20561
rect 22003 20552 22061 20558
rect 22003 20549 22015 20552
rect 20906 20521 22015 20549
rect 20906 20509 20912 20521
rect 22003 20518 22015 20521
rect 22049 20549 22061 20552
rect 22195 20552 22253 20558
rect 22195 20549 22207 20552
rect 22049 20521 22207 20549
rect 22049 20518 22061 20521
rect 22003 20512 22061 20518
rect 22195 20518 22207 20521
rect 22241 20518 22253 20552
rect 22195 20512 22253 20518
rect 10864 20287 10870 20339
rect 10922 20327 10928 20339
rect 17968 20327 17974 20339
rect 10922 20299 17974 20327
rect 10922 20287 10928 20299
rect 17968 20287 17974 20299
rect 18026 20287 18032 20339
rect 9811 20108 9869 20114
rect 9811 20074 9823 20108
rect 9857 20105 9869 20108
rect 21520 20105 21526 20117
rect 9857 20077 21526 20105
rect 9857 20074 9869 20077
rect 9811 20068 9869 20074
rect 21520 20065 21526 20077
rect 21578 20065 21584 20117
rect 43888 20065 43894 20117
rect 43946 20105 43952 20117
rect 45139 20108 45197 20114
rect 45139 20105 45151 20108
rect 43946 20077 45151 20105
rect 43946 20065 43952 20077
rect 45139 20074 45151 20077
rect 45185 20074 45197 20108
rect 49648 20105 49654 20117
rect 49609 20077 49654 20105
rect 45139 20068 45197 20074
rect 49648 20065 49654 20077
rect 49706 20065 49712 20117
rect 1152 20006 58848 20028
rect 1152 19954 4294 20006
rect 4346 19954 4358 20006
rect 4410 19954 4422 20006
rect 4474 19954 4486 20006
rect 4538 19954 35014 20006
rect 35066 19954 35078 20006
rect 35130 19954 35142 20006
rect 35194 19954 35206 20006
rect 35258 19954 58848 20006
rect 1152 19932 58848 19954
rect 7603 19886 7661 19892
rect 7603 19852 7615 19886
rect 7649 19883 7661 19886
rect 8179 19886 8237 19892
rect 8179 19883 8191 19886
rect 7649 19855 8191 19883
rect 7649 19852 7661 19855
rect 7603 19846 7661 19852
rect 8179 19852 8191 19855
rect 8225 19852 8237 19886
rect 53968 19883 53974 19895
rect 8179 19846 8237 19852
rect 8626 19855 53974 19883
rect 8272 19769 8278 19821
rect 8330 19769 8336 19821
rect 8371 19812 8429 19818
rect 8371 19778 8383 19812
rect 8417 19809 8429 19812
rect 8626 19809 8654 19855
rect 53968 19843 53974 19855
rect 54026 19843 54032 19895
rect 8417 19795 8654 19809
rect 8417 19781 8640 19795
rect 8417 19778 8429 19781
rect 8371 19772 8429 19778
rect 38224 19769 38230 19821
rect 38282 19809 38288 19821
rect 45040 19809 45046 19821
rect 38282 19781 45046 19809
rect 38282 19769 38288 19781
rect 45040 19769 45046 19781
rect 45098 19769 45104 19821
rect 8290 19735 8318 19769
rect 8256 19707 8318 19735
rect 17776 19695 17782 19747
rect 17834 19735 17840 19747
rect 43984 19735 43990 19747
rect 17834 19707 43990 19735
rect 17834 19695 17840 19707
rect 43984 19695 43990 19707
rect 44042 19695 44048 19747
rect 12115 19664 12173 19670
rect 12115 19630 12127 19664
rect 12161 19661 12173 19664
rect 12403 19664 12461 19670
rect 12403 19661 12415 19664
rect 12161 19633 12415 19661
rect 12161 19630 12173 19633
rect 12115 19624 12173 19630
rect 12403 19630 12415 19633
rect 12449 19661 12461 19664
rect 45808 19661 45814 19673
rect 12449 19633 45814 19661
rect 12449 19630 12461 19633
rect 12403 19624 12461 19630
rect 45808 19621 45814 19633
rect 45866 19621 45872 19673
rect 10960 19547 10966 19599
rect 11018 19587 11024 19599
rect 18931 19590 18989 19596
rect 18931 19587 18943 19590
rect 11018 19559 18943 19587
rect 11018 19547 11024 19559
rect 18931 19556 18943 19559
rect 18977 19556 18989 19590
rect 30547 19590 30605 19596
rect 30547 19587 30559 19590
rect 18931 19550 18989 19556
rect 27346 19559 30559 19587
rect 7936 19473 7942 19525
rect 7994 19473 8000 19525
rect 20848 19399 20854 19451
rect 20906 19439 20912 19451
rect 27346 19439 27374 19559
rect 30547 19556 30559 19559
rect 30593 19556 30605 19590
rect 30547 19550 30605 19556
rect 20906 19411 27374 19439
rect 20906 19399 20912 19411
rect 1152 19340 58848 19362
rect 1152 19288 19654 19340
rect 19706 19288 19718 19340
rect 19770 19288 19782 19340
rect 19834 19288 19846 19340
rect 19898 19288 50374 19340
rect 50426 19288 50438 19340
rect 50490 19288 50502 19340
rect 50554 19288 50566 19340
rect 50618 19288 58848 19340
rect 1152 19266 58848 19288
rect 7984 19177 7990 19229
rect 8042 19217 8048 19229
rect 48688 19217 48694 19229
rect 8042 19189 48694 19217
rect 8042 19177 8048 19189
rect 48688 19177 48694 19189
rect 48746 19177 48752 19229
rect 8272 19029 8278 19081
rect 8330 19069 8336 19081
rect 50800 19069 50806 19081
rect 8330 19041 50806 19069
rect 8330 19029 8336 19041
rect 50800 19029 50806 19041
rect 50858 19029 50864 19081
rect 8656 18955 8662 19007
rect 8714 18995 8720 19007
rect 13456 18995 13462 19007
rect 8714 18967 13462 18995
rect 8714 18955 8720 18967
rect 13456 18955 13462 18967
rect 13514 18955 13520 19007
rect 25936 18807 25942 18859
rect 25994 18847 26000 18859
rect 27856 18847 27862 18859
rect 25994 18819 27862 18847
rect 25994 18807 26000 18819
rect 27856 18807 27862 18819
rect 27914 18807 27920 18859
rect 7699 18776 7757 18782
rect 7699 18742 7711 18776
rect 7745 18773 7757 18776
rect 34672 18773 34678 18785
rect 7745 18745 34678 18773
rect 7745 18742 7757 18745
rect 7699 18736 7757 18742
rect 34672 18733 34678 18745
rect 34730 18733 34736 18785
rect 44947 18776 45005 18782
rect 44947 18742 44959 18776
rect 44993 18773 45005 18776
rect 54640 18773 54646 18785
rect 44993 18745 54646 18773
rect 44993 18742 45005 18745
rect 44947 18736 45005 18742
rect 54640 18733 54646 18745
rect 54698 18733 54704 18785
rect 1152 18674 58848 18696
rect 1152 18622 4294 18674
rect 4346 18622 4358 18674
rect 4410 18622 4422 18674
rect 4474 18622 4486 18674
rect 4538 18622 35014 18674
rect 35066 18622 35078 18674
rect 35130 18622 35142 18674
rect 35194 18622 35206 18674
rect 35258 18622 58848 18674
rect 1152 18600 58848 18622
rect 8371 18554 8429 18560
rect 8371 18551 8383 18554
rect 8194 18523 8383 18551
rect 8194 18489 8222 18523
rect 8371 18520 8383 18523
rect 8417 18520 8429 18554
rect 8371 18514 8429 18520
rect 8176 18437 8182 18489
rect 8234 18437 8240 18489
rect 8563 18480 8621 18486
rect 8563 18446 8575 18480
rect 8609 18477 8621 18480
rect 48592 18477 48598 18489
rect 8609 18449 48598 18477
rect 8609 18446 8621 18449
rect 8563 18440 8621 18446
rect 48592 18437 48598 18449
rect 48650 18437 48656 18489
rect 17296 18215 17302 18267
rect 17354 18255 17360 18267
rect 18259 18258 18317 18264
rect 18259 18255 18271 18258
rect 17354 18227 18271 18255
rect 17354 18215 17360 18227
rect 18259 18224 18271 18227
rect 18305 18224 18317 18258
rect 30832 18255 30838 18267
rect 30793 18227 30838 18255
rect 18259 18218 18317 18224
rect 30832 18215 30838 18227
rect 30890 18215 30896 18267
rect 42832 18255 42838 18267
rect 42793 18227 42838 18255
rect 42832 18215 42838 18227
rect 42890 18215 42896 18267
rect 46003 18258 46061 18264
rect 46003 18224 46015 18258
rect 46049 18224 46061 18258
rect 46003 18218 46061 18224
rect 7936 18141 7942 18193
rect 7994 18141 8000 18193
rect 8368 18181 8374 18193
rect 8256 18153 8374 18181
rect 8368 18141 8374 18153
rect 8426 18141 8432 18193
rect 12016 18181 12022 18193
rect 8544 18153 12022 18181
rect 12016 18141 12022 18153
rect 12074 18141 12080 18193
rect 7603 18110 7661 18116
rect 7603 18076 7615 18110
rect 7649 18107 7661 18110
rect 8176 18107 8182 18119
rect 7649 18079 8182 18107
rect 7649 18076 7661 18079
rect 7603 18070 7661 18076
rect 8176 18067 8182 18079
rect 8234 18067 8240 18119
rect 45808 18107 45814 18119
rect 45769 18079 45814 18107
rect 45808 18067 45814 18079
rect 45866 18107 45872 18119
rect 46018 18107 46046 18218
rect 45866 18079 46046 18107
rect 45866 18067 45872 18079
rect 1152 18008 58848 18030
rect 1152 17956 19654 18008
rect 19706 17956 19718 18008
rect 19770 17956 19782 18008
rect 19834 17956 19846 18008
rect 19898 17956 50374 18008
rect 50426 17956 50438 18008
rect 50490 17956 50502 18008
rect 50554 17956 50566 18008
rect 50618 17956 58848 18008
rect 1152 17934 58848 17956
rect 12016 17771 12022 17823
rect 12074 17811 12080 17823
rect 42928 17811 42934 17823
rect 12074 17783 42934 17811
rect 12074 17771 12080 17783
rect 42928 17771 42934 17783
rect 42986 17771 42992 17823
rect 8368 17697 8374 17749
rect 8426 17737 8432 17749
rect 44752 17737 44758 17749
rect 8426 17709 44758 17737
rect 8426 17697 8432 17709
rect 44752 17697 44758 17709
rect 44810 17697 44816 17749
rect 7984 17623 7990 17675
rect 8042 17663 8048 17675
rect 46096 17663 46102 17675
rect 8042 17635 46102 17663
rect 8042 17623 8048 17635
rect 46096 17623 46102 17635
rect 46154 17623 46160 17675
rect 5200 17549 5206 17601
rect 5258 17589 5264 17601
rect 22291 17592 22349 17598
rect 22291 17589 22303 17592
rect 5258 17561 22303 17589
rect 5258 17549 5264 17561
rect 22291 17558 22303 17561
rect 22337 17589 22349 17592
rect 22483 17592 22541 17598
rect 22483 17589 22495 17592
rect 22337 17561 22495 17589
rect 22337 17558 22349 17561
rect 22291 17552 22349 17558
rect 22483 17558 22495 17561
rect 22529 17558 22541 17592
rect 22483 17552 22541 17558
rect 8560 17475 8566 17527
rect 8618 17515 8624 17527
rect 45808 17515 45814 17527
rect 8618 17487 45814 17515
rect 8618 17475 8624 17487
rect 45808 17475 45814 17487
rect 45866 17475 45872 17527
rect 12400 17401 12406 17453
rect 12458 17441 12464 17453
rect 23347 17444 23405 17450
rect 23347 17441 23359 17444
rect 12458 17413 23359 17441
rect 12458 17401 12464 17413
rect 23347 17410 23359 17413
rect 23393 17410 23405 17444
rect 23347 17404 23405 17410
rect 1152 17342 58848 17364
rect 1152 17290 4294 17342
rect 4346 17290 4358 17342
rect 4410 17290 4422 17342
rect 4474 17290 4486 17342
rect 4538 17290 35014 17342
rect 35066 17290 35078 17342
rect 35130 17290 35142 17342
rect 35194 17290 35206 17342
rect 35258 17290 58848 17342
rect 1152 17268 58848 17290
rect 7603 17222 7661 17228
rect 7603 17188 7615 17222
rect 7649 17219 7661 17222
rect 7891 17222 7949 17228
rect 7891 17219 7903 17222
rect 7649 17191 7903 17219
rect 7649 17188 7661 17191
rect 7603 17182 7661 17188
rect 7891 17188 7903 17191
rect 7937 17188 7949 17222
rect 7891 17182 7949 17188
rect 8179 17222 8237 17228
rect 8179 17188 8191 17222
rect 8225 17219 8237 17222
rect 8225 17191 17294 17219
rect 8225 17188 8237 17191
rect 8179 17182 8237 17188
rect 8194 17131 8222 17182
rect 17266 17145 17294 17191
rect 42640 17145 42646 17157
rect 17266 17117 42646 17145
rect 42640 17105 42646 17117
rect 42698 17105 42704 17157
rect 21520 17031 21526 17083
rect 21578 17071 21584 17083
rect 48592 17071 48598 17083
rect 21578 17043 48598 17071
rect 21578 17031 21584 17043
rect 48592 17031 48598 17043
rect 48650 17031 48656 17083
rect 11056 16957 11062 17009
rect 11114 16997 11120 17009
rect 35347 17000 35405 17006
rect 35347 16997 35359 17000
rect 11114 16969 35359 16997
rect 11114 16957 11120 16969
rect 35347 16966 35359 16969
rect 35393 16997 35405 17000
rect 35539 17000 35597 17006
rect 35539 16997 35551 17000
rect 35393 16969 35551 16997
rect 35393 16966 35405 16969
rect 35347 16960 35405 16966
rect 35539 16966 35551 16969
rect 35585 16966 35597 17000
rect 35539 16960 35597 16966
rect 19411 16926 19469 16932
rect 19411 16892 19423 16926
rect 19457 16923 19469 16926
rect 21520 16923 21526 16935
rect 19457 16895 21526 16923
rect 19457 16892 19469 16895
rect 19411 16886 19469 16892
rect 21520 16883 21526 16895
rect 21578 16883 21584 16935
rect 12016 16849 12022 16861
rect 7954 16775 7982 16835
rect 8256 16821 12022 16849
rect 12016 16809 12022 16821
rect 12074 16809 12080 16861
rect 8176 16775 8182 16787
rect 7954 16747 8182 16775
rect 8176 16735 8182 16747
rect 8234 16735 8240 16787
rect 1152 16676 58848 16698
rect 1152 16624 19654 16676
rect 19706 16624 19718 16676
rect 19770 16624 19782 16676
rect 19834 16624 19846 16676
rect 19898 16624 50374 16676
rect 50426 16624 50438 16676
rect 50490 16624 50502 16676
rect 50554 16624 50566 16676
rect 50618 16624 58848 16676
rect 1152 16602 58848 16624
rect 10000 16513 10006 16565
rect 10058 16553 10064 16565
rect 42832 16553 42838 16565
rect 10058 16525 42838 16553
rect 10058 16513 10064 16525
rect 42832 16513 42838 16525
rect 42890 16513 42896 16565
rect 12016 16439 12022 16491
rect 12074 16479 12080 16491
rect 37936 16479 37942 16491
rect 12074 16451 37942 16479
rect 12074 16439 12080 16451
rect 37936 16439 37942 16451
rect 37994 16439 38000 16491
rect 8176 16365 8182 16417
rect 8234 16405 8240 16417
rect 39760 16405 39766 16417
rect 8234 16377 39766 16405
rect 8234 16365 8240 16377
rect 39760 16365 39766 16377
rect 39818 16365 39824 16417
rect 44179 16186 44237 16192
rect 44179 16152 44191 16186
rect 44225 16183 44237 16186
rect 44467 16186 44525 16192
rect 44467 16183 44479 16186
rect 44225 16155 44479 16183
rect 44225 16152 44237 16155
rect 44179 16146 44237 16152
rect 44467 16152 44479 16155
rect 44513 16183 44525 16186
rect 57328 16183 57334 16195
rect 44513 16155 57334 16183
rect 44513 16152 44525 16155
rect 44467 16146 44525 16152
rect 57328 16143 57334 16155
rect 57386 16143 57392 16195
rect 8272 16069 8278 16121
rect 8330 16109 8336 16121
rect 13936 16109 13942 16121
rect 8330 16081 13942 16109
rect 8330 16069 8336 16081
rect 13936 16069 13942 16081
rect 13994 16069 14000 16121
rect 49552 16109 49558 16121
rect 49513 16081 49558 16109
rect 49552 16069 49558 16081
rect 49610 16069 49616 16121
rect 1152 16010 58848 16032
rect 1152 15958 4294 16010
rect 4346 15958 4358 16010
rect 4410 15958 4422 16010
rect 4474 15958 4486 16010
rect 4538 15958 35014 16010
rect 35066 15958 35078 16010
rect 35130 15958 35142 16010
rect 35194 15958 35206 16010
rect 35258 15958 58848 16010
rect 1152 15936 58848 15958
rect 7714 15859 7934 15887
rect 7603 15816 7661 15822
rect 7603 15782 7615 15816
rect 7649 15813 7661 15816
rect 7714 15813 7742 15859
rect 7649 15785 7742 15813
rect 7906 15813 7934 15859
rect 16624 15847 16630 15899
rect 16682 15887 16688 15899
rect 20080 15887 20086 15899
rect 16682 15859 20086 15887
rect 16682 15847 16688 15859
rect 20080 15847 20086 15859
rect 20138 15847 20144 15899
rect 27760 15847 27766 15899
rect 27818 15887 27824 15899
rect 35059 15890 35117 15896
rect 35059 15887 35071 15890
rect 27818 15859 35071 15887
rect 27818 15847 27824 15859
rect 35059 15856 35071 15859
rect 35105 15887 35117 15890
rect 35251 15890 35309 15896
rect 35251 15887 35263 15890
rect 35105 15859 35263 15887
rect 35105 15856 35117 15859
rect 35059 15850 35117 15856
rect 35251 15856 35263 15859
rect 35297 15856 35309 15890
rect 35251 15850 35309 15856
rect 35728 15847 35734 15899
rect 35786 15887 35792 15899
rect 49552 15887 49558 15899
rect 35786 15859 49558 15887
rect 35786 15847 35792 15859
rect 49552 15847 49558 15859
rect 49610 15847 49616 15899
rect 37456 15813 37462 15825
rect 7906 15785 37462 15813
rect 7649 15782 7661 15785
rect 7603 15776 7661 15782
rect 37456 15773 37462 15785
rect 37514 15773 37520 15825
rect 8368 15591 8374 15603
rect 8257 15563 8374 15591
rect 8368 15551 8374 15563
rect 8426 15551 8432 15603
rect 34096 15517 34102 15529
rect 9120 15489 34102 15517
rect 34096 15477 34102 15489
rect 34154 15477 34160 15529
rect 8752 15403 8758 15455
rect 8810 15403 8816 15455
rect 12976 15403 12982 15455
rect 13034 15443 13040 15455
rect 34864 15443 34870 15455
rect 13034 15415 34870 15443
rect 13034 15403 13040 15415
rect 34864 15403 34870 15415
rect 34922 15403 34928 15455
rect 1152 15344 58848 15366
rect 1152 15292 19654 15344
rect 19706 15292 19718 15344
rect 19770 15292 19782 15344
rect 19834 15292 19846 15344
rect 19898 15292 50374 15344
rect 50426 15292 50438 15344
rect 50490 15292 50502 15344
rect 50554 15292 50566 15344
rect 50618 15292 58848 15344
rect 1152 15270 58848 15292
rect 8752 15181 8758 15233
rect 8810 15221 8816 15233
rect 12976 15221 12982 15233
rect 8810 15193 12982 15221
rect 8810 15181 8816 15193
rect 12976 15181 12982 15193
rect 13034 15181 13040 15233
rect 36691 15224 36749 15230
rect 36691 15190 36703 15224
rect 36737 15221 36749 15224
rect 36979 15224 37037 15230
rect 36979 15221 36991 15224
rect 36737 15193 36991 15221
rect 36737 15190 36749 15193
rect 36691 15184 36749 15190
rect 36979 15190 36991 15193
rect 37025 15221 37037 15224
rect 39856 15221 39862 15233
rect 37025 15193 39862 15221
rect 37025 15190 37037 15193
rect 36979 15184 37037 15190
rect 39856 15181 39862 15193
rect 39914 15181 39920 15233
rect 8368 15107 8374 15159
rect 8426 15147 8432 15159
rect 31888 15147 31894 15159
rect 8426 15119 31894 15147
rect 8426 15107 8432 15119
rect 31888 15107 31894 15119
rect 31946 15107 31952 15159
rect 7312 14811 7318 14863
rect 7370 14851 7376 14863
rect 36592 14851 36598 14863
rect 7370 14823 36598 14851
rect 7370 14811 7376 14823
rect 36592 14811 36598 14823
rect 36650 14811 36656 14863
rect 4048 14737 4054 14789
rect 4106 14777 4112 14789
rect 7891 14780 7949 14786
rect 7891 14777 7903 14780
rect 4106 14749 7903 14777
rect 4106 14737 4112 14749
rect 7891 14746 7903 14749
rect 7937 14746 7949 14780
rect 20464 14777 20470 14789
rect 20425 14749 20470 14777
rect 7891 14740 7949 14746
rect 20464 14737 20470 14749
rect 20522 14737 20528 14789
rect 21139 14780 21197 14786
rect 21139 14746 21151 14780
rect 21185 14777 21197 14780
rect 21232 14777 21238 14789
rect 21185 14749 21238 14777
rect 21185 14746 21197 14749
rect 21139 14740 21197 14746
rect 21232 14737 21238 14749
rect 21290 14737 21296 14789
rect 52627 14780 52685 14786
rect 52627 14746 52639 14780
rect 52673 14777 52685 14780
rect 54448 14777 54454 14789
rect 52673 14749 54454 14777
rect 52673 14746 52685 14749
rect 52627 14740 52685 14746
rect 54448 14737 54454 14749
rect 54506 14737 54512 14789
rect 1152 14678 58848 14700
rect 1152 14626 4294 14678
rect 4346 14626 4358 14678
rect 4410 14626 4422 14678
rect 4474 14626 4486 14678
rect 4538 14626 35014 14678
rect 35066 14626 35078 14678
rect 35130 14626 35142 14678
rect 35194 14626 35206 14678
rect 35258 14626 58848 14678
rect 1152 14604 58848 14626
rect 36592 14555 36598 14567
rect 8194 14527 17294 14555
rect 36553 14527 36598 14555
rect 8194 14493 8222 14527
rect 8176 14441 8182 14493
rect 8234 14441 8240 14493
rect 17266 14481 17294 14527
rect 36592 14515 36598 14527
rect 36650 14555 36656 14567
rect 36787 14558 36845 14564
rect 36787 14555 36799 14558
rect 36650 14527 36799 14555
rect 36650 14515 36656 14527
rect 36787 14524 36799 14527
rect 36833 14524 36845 14558
rect 36787 14518 36845 14524
rect 31312 14481 31318 14493
rect 17266 14453 31318 14481
rect 31312 14441 31318 14453
rect 31370 14441 31376 14493
rect 7600 14407 7606 14419
rect 7561 14379 7606 14407
rect 7600 14367 7606 14379
rect 7658 14367 7664 14419
rect 8176 14145 8182 14197
rect 8234 14145 8240 14197
rect 30832 14145 30838 14197
rect 30890 14185 30896 14197
rect 42832 14185 42838 14197
rect 30890 14157 42838 14185
rect 30890 14145 30896 14157
rect 42832 14145 42838 14157
rect 42890 14145 42896 14197
rect 34384 14071 34390 14123
rect 34442 14111 34448 14123
rect 46672 14111 46678 14123
rect 34442 14083 46678 14111
rect 34442 14071 34448 14083
rect 46672 14071 46678 14083
rect 46730 14071 46736 14123
rect 1152 14012 58848 14034
rect 1152 13960 19654 14012
rect 19706 13960 19718 14012
rect 19770 13960 19782 14012
rect 19834 13960 19846 14012
rect 19898 13960 50374 14012
rect 50426 13960 50438 14012
rect 50490 13960 50502 14012
rect 50554 13960 50566 14012
rect 50618 13960 58848 14012
rect 1152 13938 58848 13960
rect 27568 13849 27574 13901
rect 27626 13889 27632 13901
rect 40912 13889 40918 13901
rect 27626 13861 40918 13889
rect 27626 13849 27632 13861
rect 40912 13849 40918 13861
rect 40970 13849 40976 13901
rect 8176 13775 8182 13827
rect 8234 13815 8240 13827
rect 28816 13815 28822 13827
rect 8234 13787 28822 13815
rect 8234 13775 8240 13787
rect 28816 13775 28822 13787
rect 28874 13775 28880 13827
rect 37744 13775 37750 13827
rect 37802 13815 37808 13827
rect 51856 13815 51862 13827
rect 37802 13787 51862 13815
rect 37802 13775 37808 13787
rect 51856 13775 51862 13787
rect 51914 13775 51920 13827
rect 33808 13701 33814 13753
rect 33866 13741 33872 13753
rect 56944 13741 56950 13753
rect 33866 13713 56950 13741
rect 33866 13701 33872 13713
rect 56944 13701 56950 13713
rect 57002 13701 57008 13753
rect 26032 13627 26038 13679
rect 26090 13667 26096 13679
rect 57040 13667 57046 13679
rect 26090 13639 57046 13667
rect 26090 13627 26096 13639
rect 57040 13627 57046 13639
rect 57098 13627 57104 13679
rect 2995 13596 3053 13602
rect 2995 13562 3007 13596
rect 3041 13593 3053 13596
rect 3283 13596 3341 13602
rect 3283 13593 3295 13596
rect 3041 13565 3295 13593
rect 3041 13562 3053 13565
rect 2995 13556 3053 13562
rect 3283 13562 3295 13565
rect 3329 13593 3341 13596
rect 3329 13565 12974 13593
rect 3329 13562 3341 13565
rect 3283 13556 3341 13562
rect 7507 13522 7565 13528
rect 7507 13488 7519 13522
rect 7553 13519 7565 13522
rect 7795 13522 7853 13528
rect 7795 13519 7807 13522
rect 7553 13491 7807 13519
rect 7553 13488 7565 13491
rect 7507 13482 7565 13488
rect 7795 13488 7807 13491
rect 7841 13519 7853 13522
rect 12946 13519 12974 13565
rect 29584 13519 29590 13531
rect 7841 13491 11582 13519
rect 12946 13491 29590 13519
rect 7841 13488 7853 13491
rect 7795 13482 7853 13488
rect 6835 13448 6893 13454
rect 6835 13414 6847 13448
rect 6881 13445 6893 13448
rect 9904 13445 9910 13457
rect 6881 13417 9910 13445
rect 6881 13414 6893 13417
rect 6835 13408 6893 13414
rect 9904 13405 9910 13417
rect 9962 13405 9968 13457
rect 11440 13445 11446 13457
rect 11401 13417 11446 13445
rect 11440 13405 11446 13417
rect 11498 13405 11504 13457
rect 11554 13445 11582 13491
rect 29584 13479 29590 13491
rect 29642 13479 29648 13531
rect 57712 13445 57718 13457
rect 11554 13417 57718 13445
rect 57712 13405 57718 13417
rect 57770 13405 57776 13457
rect 1152 13346 58848 13368
rect 1152 13294 4294 13346
rect 4346 13294 4358 13346
rect 4410 13294 4422 13346
rect 4474 13294 4486 13346
rect 4538 13294 35014 13346
rect 35066 13294 35078 13346
rect 35130 13294 35142 13346
rect 35194 13294 35206 13346
rect 35258 13294 58848 13346
rect 1152 13272 58848 13294
rect 9904 13183 9910 13235
rect 9962 13223 9968 13235
rect 43696 13223 43702 13235
rect 9962 13195 43702 13223
rect 9962 13183 9968 13195
rect 43696 13183 43702 13195
rect 43754 13183 43760 13235
rect 7603 13152 7661 13158
rect 7603 13118 7615 13152
rect 7649 13149 7661 13152
rect 28144 13149 28150 13161
rect 7649 13121 28150 13149
rect 7649 13118 7661 13121
rect 7603 13112 7661 13118
rect 28144 13109 28150 13121
rect 28202 13109 28208 13161
rect 29008 13109 29014 13161
rect 29066 13149 29072 13161
rect 32656 13149 32662 13161
rect 29066 13121 32662 13149
rect 29066 13109 29072 13121
rect 32656 13109 32662 13121
rect 32714 13109 32720 13161
rect 8560 13035 8566 13087
rect 8618 13075 8624 13087
rect 13744 13075 13750 13087
rect 8618 13047 13750 13075
rect 8618 13035 8624 13047
rect 13744 13035 13750 13047
rect 13802 13035 13808 13087
rect 12880 12961 12886 13013
rect 12938 13001 12944 13013
rect 29011 13004 29069 13010
rect 29011 13001 29023 13004
rect 12938 12973 29023 13001
rect 12938 12961 12944 12973
rect 29011 12970 29023 12973
rect 29057 12970 29069 13004
rect 29011 12964 29069 12970
rect 30160 12961 30166 13013
rect 30218 13001 30224 13013
rect 57907 13004 57965 13010
rect 57907 13001 57919 13004
rect 30218 12973 57919 13001
rect 30218 12961 30224 12973
rect 57907 12970 57919 12973
rect 57953 12970 57965 13004
rect 57907 12964 57965 12970
rect 26320 12853 26326 12865
rect 7968 12825 26326 12853
rect 26320 12813 26326 12825
rect 26378 12813 26384 12865
rect 1152 12680 58848 12702
rect 1152 12628 19654 12680
rect 19706 12628 19718 12680
rect 19770 12628 19782 12680
rect 19834 12628 19846 12680
rect 19898 12628 50374 12680
rect 50426 12628 50438 12680
rect 50490 12628 50502 12680
rect 50554 12628 50566 12680
rect 50618 12628 58848 12680
rect 1152 12606 58848 12628
rect 20272 12517 20278 12569
rect 20330 12557 20336 12569
rect 20848 12557 20854 12569
rect 20330 12529 20854 12557
rect 20330 12517 20336 12529
rect 20848 12517 20854 12529
rect 20906 12517 20912 12569
rect 57232 12517 57238 12569
rect 57290 12557 57296 12569
rect 57331 12560 57389 12566
rect 57331 12557 57343 12560
rect 57290 12529 57343 12557
rect 57290 12517 57296 12529
rect 57331 12526 57343 12529
rect 57377 12526 57389 12560
rect 57331 12520 57389 12526
rect 20656 12369 20662 12421
rect 20714 12409 20720 12421
rect 20848 12409 20854 12421
rect 20714 12381 20854 12409
rect 20714 12369 20720 12381
rect 20848 12369 20854 12381
rect 20906 12369 20912 12421
rect 51088 12369 51094 12421
rect 51146 12409 51152 12421
rect 52816 12409 52822 12421
rect 51146 12381 52822 12409
rect 51146 12369 51152 12381
rect 52816 12369 52822 12381
rect 52874 12369 52880 12421
rect 57346 12409 57374 12520
rect 57619 12412 57677 12418
rect 57619 12409 57631 12412
rect 57346 12381 57631 12409
rect 57619 12378 57631 12381
rect 57665 12409 57677 12412
rect 57907 12412 57965 12418
rect 57907 12409 57919 12412
rect 57665 12381 57919 12409
rect 57665 12378 57677 12381
rect 57619 12372 57677 12378
rect 57907 12378 57919 12381
rect 57953 12378 57965 12412
rect 57907 12372 57965 12378
rect 2320 12295 2326 12347
rect 2378 12335 2384 12347
rect 44176 12335 44182 12347
rect 2378 12307 44182 12335
rect 2378 12295 2384 12307
rect 44176 12295 44182 12307
rect 44234 12295 44240 12347
rect 57715 12264 57773 12270
rect 57715 12230 57727 12264
rect 57761 12230 57773 12264
rect 57715 12224 57773 12230
rect 7792 12147 7798 12199
rect 7850 12187 7856 12199
rect 24976 12187 24982 12199
rect 7850 12159 24982 12187
rect 7850 12147 7856 12159
rect 24976 12147 24982 12159
rect 25034 12147 25040 12199
rect 57520 12147 57526 12199
rect 57578 12187 57584 12199
rect 57730 12187 57758 12224
rect 57578 12159 57758 12187
rect 57578 12147 57584 12159
rect 20368 12113 20374 12125
rect 20329 12085 20374 12113
rect 20368 12073 20374 12085
rect 20426 12073 20432 12125
rect 31024 12113 31030 12125
rect 30985 12085 31030 12113
rect 31024 12073 31030 12085
rect 31082 12073 31088 12125
rect 41776 12073 41782 12125
rect 41834 12113 41840 12125
rect 44563 12116 44621 12122
rect 44563 12113 44575 12116
rect 41834 12085 44575 12113
rect 41834 12073 41840 12085
rect 44563 12082 44575 12085
rect 44609 12082 44621 12116
rect 44563 12076 44621 12082
rect 44752 12073 44758 12125
rect 44810 12113 44816 12125
rect 45328 12113 45334 12125
rect 44810 12085 45334 12113
rect 44810 12073 44816 12085
rect 45328 12073 45334 12085
rect 45386 12073 45392 12125
rect 1152 12014 58848 12036
rect 1152 11962 4294 12014
rect 4346 11962 4358 12014
rect 4410 11962 4422 12014
rect 4474 11962 4486 12014
rect 4538 11962 35014 12014
rect 35066 11962 35078 12014
rect 35130 11962 35142 12014
rect 35194 11962 35206 12014
rect 35258 11962 58848 12014
rect 1152 11940 58848 11962
rect 2035 11894 2093 11900
rect 2035 11860 2047 11894
rect 2081 11891 2093 11894
rect 2320 11891 2326 11903
rect 2081 11863 2326 11891
rect 2081 11860 2093 11863
rect 2035 11854 2093 11860
rect 2320 11851 2326 11863
rect 2378 11851 2384 11903
rect 2704 11851 2710 11903
rect 2762 11891 2768 11903
rect 55507 11894 55565 11900
rect 55507 11891 55519 11894
rect 2762 11863 55519 11891
rect 2762 11851 2768 11863
rect 55507 11860 55519 11863
rect 55553 11891 55565 11894
rect 55553 11863 55742 11891
rect 55553 11860 55565 11863
rect 55507 11854 55565 11860
rect 7603 11820 7661 11826
rect 7603 11786 7615 11820
rect 7649 11817 7661 11820
rect 7792 11817 7798 11829
rect 7649 11789 7798 11817
rect 7649 11786 7661 11789
rect 7603 11780 7661 11786
rect 7792 11777 7798 11789
rect 7850 11777 7856 11829
rect 20368 11777 20374 11829
rect 20426 11817 20432 11829
rect 50800 11817 50806 11829
rect 20426 11789 50806 11817
rect 20426 11777 20432 11789
rect 50800 11777 50806 11789
rect 50858 11777 50864 11829
rect 7968 11715 17294 11743
rect 2512 11629 2518 11681
rect 2570 11669 2576 11681
rect 3568 11669 3574 11681
rect 2570 11641 3574 11669
rect 2570 11629 2576 11641
rect 3568 11629 3574 11641
rect 3626 11629 3632 11681
rect 2992 11595 2998 11607
rect 2953 11567 2998 11595
rect 2992 11555 2998 11567
rect 3050 11555 3056 11607
rect 17266 11595 17294 11715
rect 24496 11703 24502 11755
rect 24554 11743 24560 11755
rect 31024 11743 31030 11755
rect 24554 11715 31030 11743
rect 24554 11703 24560 11715
rect 31024 11703 31030 11715
rect 31082 11703 31088 11755
rect 33907 11746 33965 11752
rect 33907 11712 33919 11746
rect 33953 11743 33965 11746
rect 39763 11746 39821 11752
rect 33953 11715 39326 11743
rect 33953 11712 33965 11715
rect 33907 11706 33965 11712
rect 27952 11629 27958 11681
rect 28010 11669 28016 11681
rect 39298 11669 39326 11715
rect 39763 11712 39775 11746
rect 39809 11743 39821 11746
rect 40051 11746 40109 11752
rect 40051 11743 40063 11746
rect 39809 11715 40063 11743
rect 39809 11712 39821 11715
rect 39763 11706 39821 11712
rect 40051 11712 40063 11715
rect 40097 11743 40109 11746
rect 44752 11743 44758 11755
rect 40097 11715 44758 11743
rect 40097 11712 40109 11715
rect 40051 11706 40109 11712
rect 44752 11703 44758 11715
rect 44810 11703 44816 11755
rect 44848 11703 44854 11755
rect 44906 11743 44912 11755
rect 55714 11752 55742 11863
rect 55699 11746 55757 11752
rect 44906 11715 54878 11743
rect 44906 11703 44912 11715
rect 52624 11669 52630 11681
rect 28010 11641 37454 11669
rect 39298 11641 52630 11669
rect 28010 11629 28016 11641
rect 23344 11595 23350 11607
rect 17266 11567 23350 11595
rect 23344 11555 23350 11567
rect 23402 11555 23408 11607
rect 31504 11555 31510 11607
rect 31562 11595 31568 11607
rect 36496 11595 36502 11607
rect 31562 11567 36502 11595
rect 31562 11555 31568 11567
rect 36496 11555 36502 11567
rect 36554 11555 36560 11607
rect 37426 11595 37454 11641
rect 52624 11629 52630 11641
rect 52682 11629 52688 11681
rect 54850 11669 54878 11715
rect 55699 11712 55711 11746
rect 55745 11712 55757 11746
rect 55699 11706 55757 11712
rect 56563 11746 56621 11752
rect 56563 11712 56575 11746
rect 56609 11743 56621 11746
rect 56609 11715 57614 11743
rect 56609 11712 56621 11715
rect 56563 11706 56621 11712
rect 56947 11672 57005 11678
rect 56947 11669 56959 11672
rect 54850 11641 56959 11669
rect 56947 11638 56959 11641
rect 56993 11669 57005 11672
rect 57235 11672 57293 11678
rect 57235 11669 57247 11672
rect 56993 11641 57247 11669
rect 56993 11638 57005 11641
rect 56947 11632 57005 11638
rect 57235 11638 57247 11641
rect 57281 11638 57293 11672
rect 57235 11632 57293 11638
rect 56179 11598 56237 11604
rect 56179 11595 56191 11598
rect 37426 11567 39998 11595
rect 20848 11481 20854 11533
rect 20906 11521 20912 11533
rect 24112 11521 24118 11533
rect 20906 11493 24118 11521
rect 20906 11481 20912 11493
rect 24112 11481 24118 11493
rect 24170 11481 24176 11533
rect 39970 11521 39998 11567
rect 40162 11567 56191 11595
rect 40162 11521 40190 11567
rect 56179 11564 56191 11567
rect 56225 11595 56237 11598
rect 56467 11598 56525 11604
rect 56467 11595 56479 11598
rect 56225 11567 56479 11595
rect 56225 11564 56237 11567
rect 56179 11558 56237 11564
rect 56467 11564 56479 11567
rect 56513 11595 56525 11598
rect 56755 11598 56813 11604
rect 56755 11595 56767 11598
rect 56513 11567 56767 11595
rect 56513 11564 56525 11567
rect 56467 11558 56525 11564
rect 56755 11564 56767 11567
rect 56801 11564 56813 11598
rect 57586 11595 57614 11715
rect 59728 11595 59734 11607
rect 57586 11567 59734 11595
rect 56755 11558 56813 11564
rect 59728 11555 59734 11567
rect 59786 11555 59792 11607
rect 39970 11493 40190 11521
rect 56272 11407 56278 11459
rect 56330 11447 56336 11459
rect 57331 11450 57389 11456
rect 57331 11447 57343 11450
rect 56330 11419 57343 11447
rect 56330 11407 56336 11419
rect 57331 11416 57343 11419
rect 57377 11416 57389 11450
rect 57331 11410 57389 11416
rect 1152 11348 58848 11370
rect 1152 11296 19654 11348
rect 19706 11296 19718 11348
rect 19770 11296 19782 11348
rect 19834 11296 19846 11348
rect 19898 11296 50374 11348
rect 50426 11296 50438 11348
rect 50490 11296 50502 11348
rect 50554 11296 50566 11348
rect 50618 11296 58848 11348
rect 1152 11274 58848 11296
rect 54640 11037 54646 11089
rect 54698 11077 54704 11089
rect 56083 11080 56141 11086
rect 56083 11077 56095 11080
rect 54698 11049 56095 11077
rect 54698 11037 54704 11049
rect 56083 11046 56095 11049
rect 56129 11046 56141 11080
rect 57904 11077 57910 11089
rect 56083 11040 56141 11046
rect 57586 11049 57910 11077
rect 17008 10963 17014 11015
rect 17066 11003 17072 11015
rect 30160 11003 30166 11015
rect 17066 10975 30166 11003
rect 17066 10963 17072 10975
rect 30160 10963 30166 10975
rect 30218 10963 30224 11015
rect 57043 11006 57101 11012
rect 57043 10972 57055 11006
rect 57089 11003 57101 11006
rect 57331 11006 57389 11012
rect 57331 11003 57343 11006
rect 57089 10975 57343 11003
rect 57089 10972 57101 10975
rect 57043 10966 57101 10972
rect 57331 10972 57343 10975
rect 57377 11003 57389 11006
rect 57586 11003 57614 11049
rect 57904 11037 57910 11049
rect 57962 11037 57968 11089
rect 57377 10975 57614 11003
rect 57377 10972 57389 10975
rect 57331 10966 57389 10972
rect 21520 10889 21526 10941
rect 21578 10929 21584 10941
rect 34576 10929 34582 10941
rect 21578 10901 34582 10929
rect 21578 10889 21584 10901
rect 34576 10889 34582 10901
rect 34634 10889 34640 10941
rect 55987 10932 56045 10938
rect 55987 10898 55999 10932
rect 56033 10898 56045 10932
rect 55987 10892 56045 10898
rect 2992 10815 2998 10867
rect 3050 10855 3056 10867
rect 41200 10855 41206 10867
rect 3050 10827 41206 10855
rect 3050 10815 3056 10827
rect 41200 10815 41206 10827
rect 41258 10815 41264 10867
rect 41875 10858 41933 10864
rect 41875 10824 41887 10858
rect 41921 10855 41933 10858
rect 48784 10855 48790 10867
rect 41921 10827 48790 10855
rect 41921 10824 41933 10827
rect 41875 10818 41933 10824
rect 48784 10815 48790 10827
rect 48842 10815 48848 10867
rect 56002 10855 56030 10892
rect 56752 10889 56758 10941
rect 56810 10929 56816 10941
rect 57235 10932 57293 10938
rect 57235 10929 57247 10932
rect 56810 10901 57247 10929
rect 56810 10889 56816 10901
rect 57235 10898 57247 10901
rect 57281 10898 57293 10932
rect 57235 10892 57293 10898
rect 56848 10855 56854 10867
rect 56002 10827 56854 10855
rect 56848 10815 56854 10827
rect 56906 10815 56912 10867
rect 2899 10784 2957 10790
rect 2899 10750 2911 10784
rect 2945 10781 2957 10784
rect 3187 10784 3245 10790
rect 3187 10781 3199 10784
rect 2945 10753 3199 10781
rect 2945 10750 2957 10753
rect 2899 10744 2957 10750
rect 3187 10750 3199 10753
rect 3233 10781 3245 10784
rect 40432 10781 40438 10793
rect 3233 10753 40438 10781
rect 3233 10750 3245 10753
rect 3187 10744 3245 10750
rect 40432 10741 40438 10753
rect 40490 10741 40496 10793
rect 44752 10781 44758 10793
rect 44713 10753 44758 10781
rect 44752 10741 44758 10753
rect 44810 10741 44816 10793
rect 51856 10741 51862 10793
rect 51914 10781 51920 10793
rect 54739 10784 54797 10790
rect 54739 10781 54751 10784
rect 51914 10753 54751 10781
rect 51914 10741 51920 10753
rect 54739 10750 54751 10753
rect 54785 10750 54797 10784
rect 54739 10744 54797 10750
rect 1152 10682 58848 10704
rect 1152 10630 4294 10682
rect 4346 10630 4358 10682
rect 4410 10630 4422 10682
rect 4474 10630 4486 10682
rect 4538 10630 35014 10682
rect 35066 10630 35078 10682
rect 35130 10630 35142 10682
rect 35194 10630 35206 10682
rect 35258 10630 58848 10682
rect 1152 10608 58848 10630
rect 58576 10559 58582 10571
rect 57586 10531 58582 10559
rect 11440 10445 11446 10497
rect 11498 10485 11504 10497
rect 56947 10488 57005 10494
rect 56947 10485 56959 10488
rect 11498 10457 56959 10485
rect 11498 10445 11504 10457
rect 56947 10454 56959 10457
rect 56993 10485 57005 10488
rect 57043 10488 57101 10494
rect 57043 10485 57055 10488
rect 56993 10457 57055 10485
rect 56993 10454 57005 10457
rect 56947 10448 57005 10454
rect 57043 10454 57055 10457
rect 57089 10454 57101 10488
rect 57043 10448 57101 10454
rect 12304 10411 12310 10423
rect 7968 10383 12310 10411
rect 12304 10371 12310 10383
rect 12362 10371 12368 10423
rect 54835 10414 54893 10420
rect 54835 10380 54847 10414
rect 54881 10411 54893 10414
rect 55024 10411 55030 10423
rect 54881 10383 55030 10411
rect 54881 10380 54893 10383
rect 54835 10374 54893 10380
rect 55024 10371 55030 10383
rect 55082 10371 55088 10423
rect 55123 10414 55181 10420
rect 55123 10380 55135 10414
rect 55169 10411 55181 10414
rect 57586 10411 57614 10531
rect 58576 10519 58582 10531
rect 58634 10519 58640 10571
rect 55169 10383 57614 10411
rect 55169 10380 55181 10383
rect 55123 10374 55181 10380
rect 22384 10297 22390 10349
rect 22442 10337 22448 10349
rect 55507 10340 55565 10346
rect 55507 10337 55519 10340
rect 22442 10309 55519 10337
rect 22442 10297 22448 10309
rect 55507 10306 55519 10309
rect 55553 10337 55565 10340
rect 55795 10340 55853 10346
rect 55795 10337 55807 10340
rect 55553 10309 55807 10337
rect 55553 10306 55565 10309
rect 55507 10300 55565 10306
rect 55795 10306 55807 10309
rect 55841 10337 55853 10340
rect 56083 10340 56141 10346
rect 56083 10337 56095 10340
rect 55841 10309 56095 10337
rect 55841 10306 55853 10309
rect 55795 10300 55853 10306
rect 56083 10306 56095 10309
rect 56129 10306 56141 10340
rect 56083 10300 56141 10306
rect 56947 10340 57005 10346
rect 56947 10306 56959 10340
rect 56993 10337 57005 10340
rect 57331 10340 57389 10346
rect 57331 10337 57343 10340
rect 56993 10309 57343 10337
rect 56993 10306 57005 10309
rect 56947 10300 57005 10306
rect 57331 10306 57343 10309
rect 57377 10306 57389 10340
rect 57331 10300 57389 10306
rect 17584 10223 17590 10275
rect 17642 10263 17648 10275
rect 17683 10266 17741 10272
rect 17683 10263 17695 10266
rect 17642 10235 17695 10263
rect 17642 10223 17648 10235
rect 17683 10232 17695 10235
rect 17729 10232 17741 10266
rect 17683 10226 17741 10232
rect 48688 10223 48694 10275
rect 48746 10263 48752 10275
rect 56659 10266 56717 10272
rect 56659 10263 56671 10266
rect 48746 10235 56671 10263
rect 48746 10223 48752 10235
rect 56659 10232 56671 10235
rect 56705 10232 56717 10266
rect 56659 10226 56717 10232
rect 56464 10149 56470 10201
rect 56522 10189 56528 10201
rect 56522 10161 57470 10189
rect 56522 10149 56528 10161
rect 7603 10118 7661 10124
rect 7603 10084 7615 10118
rect 7649 10115 7661 10118
rect 22096 10115 22102 10127
rect 7649 10087 22102 10115
rect 7649 10084 7661 10087
rect 7603 10078 7661 10084
rect 22096 10075 22102 10087
rect 22154 10075 22160 10127
rect 35536 10075 35542 10127
rect 35594 10115 35600 10127
rect 36112 10115 36118 10127
rect 35594 10087 36118 10115
rect 35594 10075 35600 10087
rect 36112 10075 36118 10087
rect 36170 10075 36176 10127
rect 55696 10075 55702 10127
rect 55754 10115 55760 10127
rect 55891 10118 55949 10124
rect 55891 10115 55903 10118
rect 55754 10087 55903 10115
rect 55754 10075 55760 10087
rect 55891 10084 55903 10087
rect 55937 10084 55949 10118
rect 55891 10078 55949 10084
rect 56080 10075 56086 10127
rect 56138 10115 56144 10127
rect 57442 10124 57470 10161
rect 56563 10118 56621 10124
rect 56563 10115 56575 10118
rect 56138 10087 56575 10115
rect 56138 10075 56144 10087
rect 56563 10084 56575 10087
rect 56609 10084 56621 10118
rect 56563 10078 56621 10084
rect 57427 10118 57485 10124
rect 57427 10084 57439 10118
rect 57473 10084 57485 10118
rect 57427 10078 57485 10084
rect 1152 10016 58848 10038
rect 1152 9964 19654 10016
rect 19706 9964 19718 10016
rect 19770 9964 19782 10016
rect 19834 9964 19846 10016
rect 19898 9964 50374 10016
rect 50426 9964 50438 10016
rect 50490 9964 50502 10016
rect 50554 9964 50566 10016
rect 50618 9964 58848 10016
rect 1152 9942 58848 9964
rect 22960 9853 22966 9905
rect 23018 9893 23024 9905
rect 24016 9893 24022 9905
rect 23018 9865 24022 9893
rect 23018 9853 23024 9865
rect 24016 9853 24022 9865
rect 24074 9853 24080 9905
rect 32368 9853 32374 9905
rect 32426 9893 32432 9905
rect 33136 9893 33142 9905
rect 32426 9865 33142 9893
rect 32426 9853 32432 9865
rect 33136 9853 33142 9865
rect 33194 9853 33200 9905
rect 35632 9853 35638 9905
rect 35690 9893 35696 9905
rect 36208 9893 36214 9905
rect 35690 9865 36214 9893
rect 35690 9853 35696 9865
rect 36208 9853 36214 9865
rect 36266 9853 36272 9905
rect 54064 9853 54070 9905
rect 54122 9893 54128 9905
rect 54835 9896 54893 9902
rect 54835 9893 54847 9896
rect 54122 9865 54847 9893
rect 54122 9853 54128 9865
rect 54835 9862 54847 9865
rect 54881 9893 54893 9896
rect 54881 9865 54974 9893
rect 54881 9862 54893 9865
rect 54835 9856 54893 9862
rect 6064 9779 6070 9831
rect 6122 9819 6128 9831
rect 15856 9819 15862 9831
rect 6122 9791 15862 9819
rect 6122 9779 6128 9791
rect 15856 9779 15862 9791
rect 15914 9779 15920 9831
rect 21904 9779 21910 9831
rect 21962 9819 21968 9831
rect 25168 9819 25174 9831
rect 21962 9791 25174 9819
rect 21962 9779 21968 9791
rect 25168 9779 25174 9791
rect 25226 9779 25232 9831
rect 32752 9779 32758 9831
rect 32810 9819 32816 9831
rect 34000 9819 34006 9831
rect 32810 9791 34006 9819
rect 32810 9779 32816 9791
rect 34000 9779 34006 9791
rect 34058 9779 34064 9831
rect 35440 9779 35446 9831
rect 35498 9819 35504 9831
rect 36976 9819 36982 9831
rect 35498 9791 36982 9819
rect 35498 9779 35504 9791
rect 36976 9779 36982 9791
rect 37034 9779 37040 9831
rect 6256 9705 6262 9757
rect 6314 9745 6320 9757
rect 14704 9745 14710 9757
rect 6314 9717 14710 9745
rect 6314 9705 6320 9717
rect 14704 9705 14710 9717
rect 14762 9705 14768 9757
rect 19216 9705 19222 9757
rect 19274 9745 19280 9757
rect 23728 9745 23734 9757
rect 19274 9717 23734 9745
rect 19274 9705 19280 9717
rect 23728 9705 23734 9717
rect 23786 9705 23792 9757
rect 34288 9705 34294 9757
rect 34346 9745 34352 9757
rect 35728 9745 35734 9757
rect 34346 9717 35734 9745
rect 34346 9705 34352 9717
rect 35728 9705 35734 9717
rect 35786 9705 35792 9757
rect 36784 9705 36790 9757
rect 36842 9745 36848 9757
rect 54448 9745 54454 9757
rect 36842 9717 47534 9745
rect 54409 9717 54454 9745
rect 36842 9705 36848 9717
rect 5680 9631 5686 9683
rect 5738 9671 5744 9683
rect 13840 9671 13846 9683
rect 5738 9643 13846 9671
rect 5738 9631 5744 9643
rect 13840 9631 13846 9643
rect 13898 9631 13904 9683
rect 13936 9631 13942 9683
rect 13994 9671 14000 9683
rect 24496 9671 24502 9683
rect 13994 9643 24502 9671
rect 13994 9631 14000 9643
rect 24496 9631 24502 9643
rect 24554 9631 24560 9683
rect 10672 9557 10678 9609
rect 10730 9597 10736 9609
rect 24304 9597 24310 9609
rect 10730 9569 24310 9597
rect 10730 9557 10736 9569
rect 24304 9557 24310 9569
rect 24362 9557 24368 9609
rect 30352 9557 30358 9609
rect 30410 9597 30416 9609
rect 38416 9597 38422 9609
rect 30410 9569 38422 9597
rect 30410 9557 30416 9569
rect 38416 9557 38422 9569
rect 38474 9557 38480 9609
rect 47506 9597 47534 9717
rect 54448 9705 54454 9717
rect 54506 9705 54512 9757
rect 54946 9745 54974 9865
rect 57808 9819 57814 9831
rect 57586 9791 57814 9819
rect 55123 9748 55181 9754
rect 55123 9745 55135 9748
rect 54946 9717 55135 9745
rect 55123 9714 55135 9717
rect 55169 9714 55181 9748
rect 57586 9745 57614 9791
rect 57808 9779 57814 9791
rect 57866 9779 57872 9831
rect 55123 9708 55181 9714
rect 56098 9717 57614 9745
rect 49648 9631 49654 9683
rect 49706 9671 49712 9683
rect 55987 9674 56045 9680
rect 55987 9671 55999 9674
rect 49706 9643 55999 9671
rect 49706 9631 49712 9643
rect 55987 9640 55999 9643
rect 56033 9640 56045 9674
rect 55987 9634 56045 9640
rect 47506 9569 53918 9597
rect 17680 9483 17686 9535
rect 17738 9523 17744 9535
rect 32560 9523 32566 9535
rect 17738 9495 32566 9523
rect 17738 9483 17744 9495
rect 32560 9483 32566 9495
rect 32618 9483 32624 9535
rect 46675 9526 46733 9532
rect 46675 9492 46687 9526
rect 46721 9523 46733 9526
rect 46963 9526 47021 9532
rect 46963 9523 46975 9526
rect 46721 9495 46975 9523
rect 46721 9492 46733 9495
rect 46675 9486 46733 9492
rect 46963 9492 46975 9495
rect 47009 9523 47021 9526
rect 50224 9523 50230 9535
rect 47009 9495 50230 9523
rect 47009 9492 47021 9495
rect 46963 9486 47021 9492
rect 50224 9483 50230 9495
rect 50282 9483 50288 9535
rect 8272 9409 8278 9461
rect 8330 9449 8336 9461
rect 16144 9449 16150 9461
rect 8330 9421 16150 9449
rect 8330 9409 8336 9421
rect 16144 9409 16150 9421
rect 16202 9409 16208 9461
rect 16240 9409 16246 9461
rect 16298 9449 16304 9461
rect 20272 9449 20278 9461
rect 16298 9421 20278 9449
rect 16298 9409 16304 9421
rect 20272 9409 20278 9421
rect 20330 9409 20336 9461
rect 50992 9409 50998 9461
rect 51050 9449 51056 9461
rect 53107 9452 53165 9458
rect 53107 9449 53119 9452
rect 51050 9421 53119 9449
rect 51050 9409 51056 9421
rect 53107 9418 53119 9421
rect 53153 9418 53165 9452
rect 53776 9449 53782 9461
rect 53737 9421 53782 9449
rect 53107 9412 53165 9418
rect 53776 9409 53782 9421
rect 53834 9409 53840 9461
rect 53890 9449 53918 9569
rect 54256 9557 54262 9609
rect 54314 9597 54320 9609
rect 54355 9600 54413 9606
rect 54355 9597 54367 9600
rect 54314 9569 54367 9597
rect 54314 9557 54320 9569
rect 54355 9566 54367 9569
rect 54401 9566 54413 9600
rect 54355 9560 54413 9566
rect 55219 9600 55277 9606
rect 55219 9566 55231 9600
rect 55265 9566 55277 9600
rect 55219 9560 55277 9566
rect 54928 9483 54934 9535
rect 54986 9523 54992 9535
rect 55234 9523 55262 9560
rect 55312 9557 55318 9609
rect 55370 9597 55376 9609
rect 55891 9600 55949 9606
rect 55891 9597 55903 9600
rect 55370 9569 55903 9597
rect 55370 9557 55376 9569
rect 55891 9566 55903 9569
rect 55937 9566 55949 9600
rect 55891 9560 55949 9566
rect 54986 9495 55262 9523
rect 54986 9483 54992 9495
rect 56098 9449 56126 9717
rect 57616 9631 57622 9683
rect 57674 9671 57680 9683
rect 57674 9643 57719 9671
rect 57674 9631 57680 9643
rect 53890 9421 56126 9449
rect 1152 9350 58848 9372
rect 1152 9298 4294 9350
rect 4346 9298 4358 9350
rect 4410 9298 4422 9350
rect 4474 9298 4486 9350
rect 4538 9298 35014 9350
rect 35066 9298 35078 9350
rect 35130 9298 35142 9350
rect 35194 9298 35206 9350
rect 35258 9298 58848 9350
rect 1152 9276 58848 9298
rect 3091 9230 3149 9236
rect 3091 9196 3103 9230
rect 3137 9227 3149 9230
rect 3137 9199 7982 9227
rect 3137 9196 3149 9199
rect 3091 9190 3149 9196
rect 7603 9156 7661 9162
rect 7603 9122 7615 9156
rect 7649 9153 7661 9156
rect 7699 9156 7757 9162
rect 7699 9153 7711 9156
rect 7649 9125 7711 9153
rect 7649 9122 7661 9125
rect 7603 9116 7661 9122
rect 7699 9122 7711 9125
rect 7745 9122 7757 9156
rect 7954 9153 7982 9199
rect 8242 9199 12974 9227
rect 8242 9153 8270 9199
rect 8467 9156 8525 9162
rect 8467 9153 8479 9156
rect 7954 9125 8270 9153
rect 8352 9125 8479 9153
rect 7699 9116 7757 9122
rect 8467 9122 8479 9125
rect 8513 9153 8525 9156
rect 12496 9153 12502 9165
rect 8513 9125 12502 9153
rect 8513 9122 8525 9125
rect 8467 9116 8525 9122
rect 12496 9113 12502 9125
rect 12554 9113 12560 9165
rect 7942 8943 7994 8949
rect 12946 8931 12974 9199
rect 21520 9187 21526 9239
rect 21578 9227 21584 9239
rect 53776 9227 53782 9239
rect 21578 9199 53782 9227
rect 21578 9187 21584 9199
rect 53776 9187 53782 9199
rect 53834 9187 53840 9239
rect 30928 9113 30934 9165
rect 30986 9153 30992 9165
rect 37459 9156 37517 9162
rect 30986 9125 36926 9153
rect 30986 9113 30992 9125
rect 23920 9039 23926 9091
rect 23978 9079 23984 9091
rect 29680 9079 29686 9091
rect 23978 9051 29686 9079
rect 23978 9039 23984 9051
rect 29680 9039 29686 9051
rect 29738 9039 29744 9091
rect 30067 9082 30125 9088
rect 30067 9048 30079 9082
rect 30113 9079 30125 9082
rect 30352 9079 30358 9091
rect 30113 9051 30358 9079
rect 30113 9048 30125 9051
rect 30067 9042 30125 9048
rect 30352 9039 30358 9051
rect 30410 9039 30416 9091
rect 36499 9082 36557 9088
rect 36499 9048 36511 9082
rect 36545 9079 36557 9082
rect 36784 9079 36790 9091
rect 36545 9051 36790 9079
rect 36545 9048 36557 9051
rect 36499 9042 36557 9048
rect 36784 9039 36790 9051
rect 36842 9039 36848 9091
rect 36898 9079 36926 9125
rect 37459 9122 37471 9156
rect 37505 9153 37517 9156
rect 48688 9153 48694 9165
rect 37505 9125 48694 9153
rect 37505 9122 37517 9125
rect 37459 9116 37517 9122
rect 48688 9113 48694 9125
rect 48746 9113 48752 9165
rect 54643 9082 54701 9088
rect 54643 9079 54655 9082
rect 36898 9051 54655 9079
rect 54643 9048 54655 9051
rect 54689 9048 54701 9082
rect 54643 9042 54701 9048
rect 15184 8965 15190 9017
rect 15242 9005 15248 9017
rect 49363 9008 49421 9014
rect 49363 9005 49375 9008
rect 15242 8977 49375 9005
rect 15242 8965 15248 8977
rect 49363 8974 49375 8977
rect 49409 8974 49421 9008
rect 49363 8968 49421 8974
rect 53315 9008 53373 9014
rect 53315 8974 53327 9008
rect 53361 9005 53373 9008
rect 55888 9005 55894 9017
rect 53361 8977 55894 9005
rect 53361 8974 53373 8977
rect 53315 8968 53373 8974
rect 55888 8965 55894 8977
rect 55946 8965 55952 9017
rect 56563 9008 56621 9014
rect 56563 8974 56575 9008
rect 56609 8974 56621 9008
rect 57232 9005 57238 9017
rect 57193 8977 57238 9005
rect 56563 8968 56621 8974
rect 42739 8934 42797 8940
rect 42739 8931 42751 8934
rect 12946 8903 42751 8931
rect 42739 8900 42751 8903
rect 42785 8900 42797 8934
rect 42739 8894 42797 8900
rect 43024 8891 43030 8943
rect 43082 8931 43088 8943
rect 44083 8934 44141 8940
rect 44083 8931 44095 8934
rect 43082 8903 44095 8931
rect 43082 8891 43088 8903
rect 44083 8900 44095 8903
rect 44129 8900 44141 8934
rect 44083 8894 44141 8900
rect 53200 8891 53206 8943
rect 53258 8931 53264 8943
rect 53395 8934 53453 8940
rect 53395 8931 53407 8934
rect 53258 8903 53407 8931
rect 53258 8891 53264 8903
rect 53395 8900 53407 8903
rect 53441 8900 53453 8934
rect 53395 8894 53453 8900
rect 55411 8934 55469 8940
rect 55411 8900 55423 8934
rect 55457 8900 55469 8934
rect 56578 8931 56606 8968
rect 57232 8965 57238 8977
rect 57290 8965 57296 9017
rect 57328 8931 57334 8943
rect 56578 8903 57334 8931
rect 55411 8894 55469 8900
rect 7942 8885 7994 8891
rect 12592 8817 12598 8869
rect 12650 8857 12656 8869
rect 12650 8829 17294 8857
rect 12650 8817 12656 8829
rect 10192 8743 10198 8795
rect 10250 8783 10256 8795
rect 14896 8783 14902 8795
rect 10250 8755 14902 8783
rect 10250 8743 10256 8755
rect 14896 8743 14902 8755
rect 14954 8743 14960 8795
rect 17266 8783 17294 8829
rect 35056 8817 35062 8869
rect 35114 8857 35120 8869
rect 55426 8857 55454 8894
rect 57328 8891 57334 8903
rect 57386 8891 57392 8943
rect 35114 8829 55454 8857
rect 35114 8817 35120 8829
rect 18832 8783 18838 8795
rect 17266 8755 18838 8783
rect 18832 8743 18838 8755
rect 18890 8743 18896 8795
rect 42739 8786 42797 8792
rect 42739 8752 42751 8786
rect 42785 8783 42797 8786
rect 44944 8783 44950 8795
rect 42785 8755 44950 8783
rect 42785 8752 42797 8755
rect 42739 8746 42797 8752
rect 44944 8743 44950 8755
rect 45002 8743 45008 8795
rect 53872 8743 53878 8795
rect 53930 8783 53936 8795
rect 54547 8786 54605 8792
rect 54547 8783 54559 8786
rect 53930 8755 54559 8783
rect 53930 8743 53936 8755
rect 54547 8752 54559 8755
rect 54593 8752 54605 8786
rect 54547 8746 54605 8752
rect 54640 8743 54646 8795
rect 54698 8783 54704 8795
rect 55315 8786 55373 8792
rect 55315 8783 55327 8786
rect 54698 8755 55327 8783
rect 54698 8743 54704 8755
rect 55315 8752 55327 8755
rect 55361 8752 55373 8786
rect 55315 8746 55373 8752
rect 1152 8684 58848 8706
rect 1152 8632 19654 8684
rect 19706 8632 19718 8684
rect 19770 8632 19782 8684
rect 19834 8632 19846 8684
rect 19898 8632 50374 8684
rect 50426 8632 50438 8684
rect 50490 8632 50502 8684
rect 50554 8632 50566 8684
rect 50618 8632 58848 8684
rect 1152 8610 58848 8632
rect 2035 8564 2093 8570
rect 2035 8561 2047 8564
rect 1762 8533 2047 8561
rect 1762 8422 1790 8533
rect 2035 8530 2047 8533
rect 2081 8561 2093 8564
rect 3664 8561 3670 8573
rect 2081 8533 3670 8561
rect 2081 8530 2093 8533
rect 2035 8524 2093 8530
rect 3664 8521 3670 8533
rect 3722 8521 3728 8573
rect 5584 8521 5590 8573
rect 5642 8561 5648 8573
rect 5642 8533 10046 8561
rect 5642 8521 5648 8533
rect 10018 8487 10046 8533
rect 12784 8521 12790 8573
rect 12842 8561 12848 8573
rect 13555 8564 13613 8570
rect 13555 8561 13567 8564
rect 12842 8533 13567 8561
rect 12842 8521 12848 8533
rect 13555 8530 13567 8533
rect 13601 8530 13613 8564
rect 13555 8524 13613 8530
rect 14515 8564 14573 8570
rect 14515 8530 14527 8564
rect 14561 8561 14573 8564
rect 42067 8564 42125 8570
rect 14561 8533 40958 8561
rect 14561 8530 14573 8533
rect 14515 8524 14573 8530
rect 39475 8490 39533 8496
rect 39475 8487 39487 8490
rect 4546 8459 9950 8487
rect 10018 8459 39487 8487
rect 1747 8416 1805 8422
rect 1747 8382 1759 8416
rect 1793 8382 1805 8416
rect 1747 8376 1805 8382
rect 2995 8416 3053 8422
rect 2995 8382 3007 8416
rect 3041 8413 3053 8416
rect 3280 8413 3286 8425
rect 3041 8385 3286 8413
rect 3041 8382 3053 8385
rect 2995 8376 3053 8382
rect 3280 8373 3286 8385
rect 3338 8373 3344 8425
rect 4546 8422 4574 8459
rect 4243 8416 4301 8422
rect 4243 8382 4255 8416
rect 4289 8413 4301 8416
rect 4531 8416 4589 8422
rect 4531 8413 4543 8416
rect 4289 8385 4543 8413
rect 4289 8382 4301 8385
rect 4243 8376 4301 8382
rect 4531 8382 4543 8385
rect 4577 8382 4589 8416
rect 4531 8376 4589 8382
rect 7216 8299 7222 8351
rect 7274 8339 7280 8351
rect 9424 8339 9430 8351
rect 7274 8311 9430 8339
rect 7274 8299 7280 8311
rect 9424 8299 9430 8311
rect 9482 8299 9488 8351
rect 9811 8342 9869 8348
rect 9811 8339 9823 8342
rect 9634 8311 9823 8339
rect 9634 8277 9662 8311
rect 9811 8308 9823 8311
rect 9857 8308 9869 8342
rect 9922 8339 9950 8459
rect 39475 8456 39487 8459
rect 39521 8487 39533 8490
rect 40930 8487 40958 8533
rect 42067 8530 42079 8564
rect 42113 8561 42125 8564
rect 42160 8561 42166 8573
rect 42113 8533 42166 8561
rect 42113 8530 42125 8533
rect 42067 8524 42125 8530
rect 42160 8521 42166 8533
rect 42218 8521 42224 8573
rect 48592 8561 48598 8573
rect 48553 8533 48598 8561
rect 48592 8521 48598 8533
rect 48650 8521 48656 8573
rect 52435 8564 52493 8570
rect 52435 8530 52447 8564
rect 52481 8561 52493 8564
rect 58960 8561 58966 8573
rect 52481 8533 58966 8561
rect 52481 8530 52493 8533
rect 52435 8524 52493 8530
rect 58960 8521 58966 8533
rect 59018 8521 59024 8573
rect 44368 8487 44374 8499
rect 39521 8459 39710 8487
rect 40930 8459 44374 8487
rect 39521 8456 39533 8459
rect 39475 8450 39533 8456
rect 10576 8413 10582 8425
rect 10537 8385 10582 8413
rect 10576 8373 10582 8385
rect 10634 8373 10640 8425
rect 11059 8416 11117 8422
rect 11059 8382 11071 8416
rect 11105 8413 11117 8416
rect 11344 8413 11350 8425
rect 11105 8385 11350 8413
rect 11105 8382 11117 8385
rect 11059 8376 11117 8382
rect 11344 8373 11350 8385
rect 11402 8373 11408 8425
rect 11827 8416 11885 8422
rect 11827 8382 11839 8416
rect 11873 8413 11885 8416
rect 12112 8413 12118 8425
rect 11873 8385 12118 8413
rect 11873 8382 11885 8385
rect 11827 8376 11885 8382
rect 12112 8373 12118 8385
rect 12170 8373 12176 8425
rect 12880 8413 12886 8425
rect 12841 8385 12886 8413
rect 12880 8373 12886 8385
rect 12938 8373 12944 8425
rect 13648 8413 13654 8425
rect 13609 8385 13654 8413
rect 13648 8373 13654 8385
rect 13706 8373 13712 8425
rect 33904 8413 33910 8425
rect 13762 8385 33910 8413
rect 13762 8339 13790 8385
rect 33904 8373 33910 8385
rect 33962 8373 33968 8425
rect 34099 8416 34157 8422
rect 34099 8382 34111 8416
rect 34145 8413 34157 8416
rect 34384 8413 34390 8425
rect 34145 8385 34390 8413
rect 34145 8382 34157 8385
rect 34099 8376 34157 8382
rect 34384 8373 34390 8385
rect 34442 8373 34448 8425
rect 35056 8413 35062 8425
rect 35017 8385 35062 8413
rect 35056 8373 35062 8385
rect 35114 8373 35120 8425
rect 39682 8422 39710 8459
rect 44368 8447 44374 8459
rect 44426 8447 44432 8499
rect 50704 8487 50710 8499
rect 47506 8459 50710 8487
rect 39667 8416 39725 8422
rect 39667 8382 39679 8416
rect 39713 8382 39725 8416
rect 42160 8413 42166 8425
rect 42121 8385 42166 8413
rect 39667 8376 39725 8382
rect 42160 8373 42166 8385
rect 42218 8373 42224 8425
rect 16240 8339 16246 8351
rect 9922 8311 13790 8339
rect 16201 8311 16246 8339
rect 9811 8302 9869 8308
rect 16240 8299 16246 8311
rect 16298 8299 16304 8351
rect 17008 8339 17014 8351
rect 16969 8311 17014 8339
rect 17008 8299 17014 8311
rect 17066 8299 17072 8351
rect 17104 8299 17110 8351
rect 17162 8339 17168 8351
rect 47506 8339 47534 8459
rect 50704 8447 50710 8459
rect 50762 8447 50768 8499
rect 48211 8416 48269 8422
rect 48211 8382 48223 8416
rect 48257 8413 48269 8416
rect 48880 8413 48886 8425
rect 48257 8385 48886 8413
rect 48257 8382 48269 8385
rect 48211 8376 48269 8382
rect 48880 8373 48886 8385
rect 48938 8373 48944 8425
rect 52528 8413 52534 8425
rect 52489 8385 52534 8413
rect 52528 8373 52534 8385
rect 52586 8373 52592 8425
rect 53296 8413 53302 8425
rect 53257 8385 53302 8413
rect 53296 8373 53302 8385
rect 53354 8373 53360 8425
rect 59824 8413 59830 8425
rect 55234 8385 59830 8413
rect 17162 8311 47534 8339
rect 17162 8299 17168 8311
rect 48784 8299 48790 8351
rect 48842 8339 48848 8351
rect 49747 8342 49805 8348
rect 49747 8339 49759 8342
rect 48842 8311 49759 8339
rect 48842 8299 48848 8311
rect 49747 8308 49759 8311
rect 49793 8308 49805 8342
rect 49747 8302 49805 8308
rect 52912 8299 52918 8351
rect 52970 8339 52976 8351
rect 55234 8348 55262 8385
rect 59824 8373 59830 8385
rect 59882 8373 59888 8425
rect 54067 8342 54125 8348
rect 54067 8339 54079 8342
rect 52970 8311 54079 8339
rect 52970 8299 52976 8311
rect 54067 8308 54079 8311
rect 54113 8308 54125 8342
rect 54067 8302 54125 8308
rect 55219 8342 55277 8348
rect 55219 8308 55231 8342
rect 55265 8308 55277 8342
rect 55219 8302 55277 8308
rect 55987 8342 56045 8348
rect 55987 8308 55999 8342
rect 56033 8308 56045 8342
rect 55987 8302 56045 8308
rect 1648 8265 1654 8277
rect 1609 8237 1654 8265
rect 1648 8225 1654 8237
rect 1706 8225 1712 8277
rect 2128 8225 2134 8277
rect 2186 8265 2192 8277
rect 2419 8268 2477 8274
rect 2419 8265 2431 8268
rect 2186 8237 2431 8265
rect 2186 8225 2192 8237
rect 2419 8234 2431 8237
rect 2465 8234 2477 8268
rect 2419 8228 2477 8234
rect 2515 8268 2573 8274
rect 2515 8234 2527 8268
rect 2561 8265 2573 8268
rect 2704 8265 2710 8277
rect 2561 8237 2710 8265
rect 2561 8234 2573 8237
rect 2515 8228 2573 8234
rect 2704 8225 2710 8237
rect 2762 8225 2768 8277
rect 2992 8225 2998 8277
rect 3050 8265 3056 8277
rect 3187 8268 3245 8274
rect 3187 8265 3199 8268
rect 3050 8237 3199 8265
rect 3050 8225 3056 8237
rect 3187 8234 3199 8237
rect 3233 8234 3245 8268
rect 3187 8228 3245 8234
rect 4435 8268 4493 8274
rect 4435 8234 4447 8268
rect 4481 8234 4493 8268
rect 4435 8228 4493 8234
rect 4450 8191 4478 8228
rect 7696 8225 7702 8277
rect 7754 8265 7760 8277
rect 7795 8268 7853 8274
rect 7795 8265 7807 8268
rect 7754 8237 7807 8265
rect 7754 8225 7760 8237
rect 7795 8234 7807 8237
rect 7841 8234 7853 8268
rect 7795 8228 7853 8234
rect 7891 8268 7949 8274
rect 7891 8234 7903 8268
rect 7937 8234 7949 8268
rect 7891 8228 7949 8234
rect 4816 8191 4822 8203
rect 4450 8163 4822 8191
rect 4816 8151 4822 8163
rect 4874 8151 4880 8203
rect 7906 8191 7934 8228
rect 9616 8225 9622 8277
rect 9674 8225 9680 8277
rect 9712 8225 9718 8277
rect 9770 8274 9776 8277
rect 9770 8268 9789 8274
rect 9777 8234 9789 8268
rect 9770 8228 9789 8234
rect 9770 8225 9776 8228
rect 9904 8225 9910 8277
rect 9962 8265 9968 8277
rect 9962 8237 10094 8265
rect 9962 8225 9968 8237
rect 9808 8191 9814 8203
rect 7906 8163 9814 8191
rect 9808 8151 9814 8163
rect 9866 8151 9872 8203
rect 10066 8191 10094 8237
rect 10288 8225 10294 8277
rect 10346 8265 10352 8277
rect 10483 8268 10541 8274
rect 10483 8265 10495 8268
rect 10346 8237 10495 8265
rect 10346 8225 10352 8237
rect 10483 8234 10495 8237
rect 10529 8234 10541 8268
rect 10483 8228 10541 8234
rect 10576 8225 10582 8277
rect 10634 8265 10640 8277
rect 11251 8268 11309 8274
rect 11251 8265 11263 8268
rect 10634 8237 11263 8265
rect 10634 8225 10640 8237
rect 11251 8234 11263 8237
rect 11297 8234 11309 8268
rect 11251 8228 11309 8234
rect 11344 8225 11350 8277
rect 11402 8265 11408 8277
rect 12019 8268 12077 8274
rect 12019 8265 12031 8268
rect 11402 8237 12031 8265
rect 11402 8225 11408 8237
rect 12019 8234 12031 8237
rect 12065 8234 12077 8268
rect 12019 8228 12077 8234
rect 12112 8225 12118 8277
rect 12170 8265 12176 8277
rect 12787 8268 12845 8274
rect 12787 8265 12799 8268
rect 12170 8237 12799 8265
rect 12170 8225 12176 8237
rect 12787 8234 12799 8237
rect 12833 8234 12845 8268
rect 16144 8265 16150 8277
rect 16105 8237 16150 8265
rect 12787 8228 12845 8234
rect 16144 8225 16150 8237
rect 16202 8225 16208 8277
rect 16336 8225 16342 8277
rect 16394 8265 16400 8277
rect 16915 8268 16973 8274
rect 16915 8265 16927 8268
rect 16394 8237 16927 8265
rect 16394 8225 16400 8237
rect 16915 8234 16927 8237
rect 16961 8234 16973 8268
rect 16915 8228 16973 8234
rect 48016 8225 48022 8277
rect 48074 8265 48080 8277
rect 48115 8268 48173 8274
rect 48115 8265 48127 8268
rect 48074 8237 48127 8265
rect 48074 8225 48080 8237
rect 48115 8234 48127 8237
rect 48161 8234 48173 8268
rect 48115 8228 48173 8234
rect 48592 8225 48598 8277
rect 48650 8265 48656 8277
rect 48883 8268 48941 8274
rect 48883 8265 48895 8268
rect 48650 8237 48895 8265
rect 48650 8225 48656 8237
rect 48883 8234 48895 8237
rect 48929 8234 48941 8268
rect 48883 8228 48941 8234
rect 48979 8268 49037 8274
rect 48979 8234 48991 8268
rect 49025 8234 49037 8268
rect 48979 8228 49037 8234
rect 33619 8194 33677 8200
rect 33619 8191 33631 8194
rect 10066 8163 33631 8191
rect 33619 8160 33631 8163
rect 33665 8160 33677 8194
rect 33619 8154 33677 8160
rect 48688 8151 48694 8203
rect 48746 8191 48752 8203
rect 48994 8191 49022 8228
rect 49456 8225 49462 8277
rect 49514 8265 49520 8277
rect 49651 8268 49709 8274
rect 49651 8265 49663 8268
rect 49514 8237 49663 8265
rect 49514 8225 49520 8237
rect 49651 8234 49663 8237
rect 49697 8234 49709 8268
rect 49651 8228 49709 8234
rect 53104 8225 53110 8277
rect 53162 8265 53168 8277
rect 53203 8268 53261 8274
rect 53203 8265 53215 8268
rect 53162 8237 53215 8265
rect 53162 8225 53168 8237
rect 53203 8234 53215 8237
rect 53249 8234 53261 8268
rect 53203 8228 53261 8234
rect 53488 8225 53494 8277
rect 53546 8265 53552 8277
rect 53971 8268 54029 8274
rect 53971 8265 53983 8268
rect 53546 8237 53983 8265
rect 53546 8225 53552 8237
rect 53971 8234 53983 8237
rect 54017 8234 54029 8268
rect 56002 8265 56030 8302
rect 56944 8299 56950 8351
rect 57002 8339 57008 8351
rect 57139 8342 57197 8348
rect 57139 8339 57151 8342
rect 57002 8311 57151 8339
rect 57002 8299 57008 8311
rect 57139 8308 57151 8311
rect 57185 8308 57197 8342
rect 57139 8302 57197 8308
rect 58384 8265 58390 8277
rect 56002 8237 58390 8265
rect 53971 8228 54029 8234
rect 58384 8225 58390 8237
rect 58442 8225 58448 8277
rect 48746 8163 49022 8191
rect 48746 8151 48752 8163
rect 51184 8151 51190 8203
rect 51242 8191 51248 8203
rect 56656 8191 56662 8203
rect 51242 8163 56662 8191
rect 51242 8151 51248 8163
rect 56656 8151 56662 8163
rect 56714 8151 56720 8203
rect 6160 8117 6166 8129
rect 6121 8089 6166 8117
rect 6160 8077 6166 8089
rect 6218 8077 6224 8129
rect 6931 8120 6989 8126
rect 6931 8086 6943 8120
rect 6977 8117 6989 8120
rect 7600 8117 7606 8129
rect 6977 8089 7606 8117
rect 6977 8086 6989 8089
rect 6931 8080 6989 8086
rect 7600 8077 7606 8089
rect 7658 8077 7664 8129
rect 7792 8077 7798 8129
rect 7850 8117 7856 8129
rect 8560 8117 8566 8129
rect 7850 8089 8566 8117
rect 7850 8077 7856 8089
rect 8560 8077 8566 8089
rect 8618 8077 8624 8129
rect 9523 8120 9581 8126
rect 9523 8086 9535 8120
rect 9569 8117 9581 8120
rect 9616 8117 9622 8129
rect 9569 8089 9622 8117
rect 9569 8086 9581 8089
rect 9523 8080 9581 8086
rect 9616 8077 9622 8089
rect 9674 8117 9680 8129
rect 14515 8120 14573 8126
rect 14515 8117 14527 8120
rect 9674 8089 14527 8117
rect 9674 8077 9680 8089
rect 14515 8086 14527 8089
rect 14561 8086 14573 8120
rect 17776 8117 17782 8129
rect 17737 8089 17782 8117
rect 14515 8080 14573 8086
rect 17776 8077 17782 8089
rect 17834 8077 17840 8129
rect 22096 8117 22102 8129
rect 22057 8089 22102 8117
rect 22096 8077 22102 8089
rect 22154 8077 22160 8129
rect 25939 8120 25997 8126
rect 25939 8086 25951 8120
rect 25985 8117 25997 8120
rect 28048 8117 28054 8129
rect 25985 8089 28054 8117
rect 25985 8086 25997 8089
rect 25939 8080 25997 8086
rect 28048 8077 28054 8089
rect 28106 8077 28112 8129
rect 52528 8077 52534 8129
rect 52586 8117 52592 8129
rect 57712 8117 57718 8129
rect 52586 8089 57718 8117
rect 52586 8077 52592 8089
rect 57712 8077 57718 8089
rect 57770 8077 57776 8129
rect 1152 8018 58848 8040
rect 1152 7966 4294 8018
rect 4346 7966 4358 8018
rect 4410 7966 4422 8018
rect 4474 7966 4486 8018
rect 4538 7966 35014 8018
rect 35066 7966 35078 8018
rect 35130 7966 35142 8018
rect 35194 7966 35206 8018
rect 35258 7966 58848 8018
rect 1152 7944 58848 7966
rect 2896 7855 2902 7907
rect 2954 7895 2960 7907
rect 2954 7867 3326 7895
rect 2954 7855 2960 7867
rect 2512 7747 2518 7759
rect 2473 7719 2518 7747
rect 2512 7707 2518 7719
rect 2570 7707 2576 7759
rect 3298 7756 3326 7867
rect 8560 7855 8566 7907
rect 8618 7895 8624 7907
rect 8618 7867 12974 7895
rect 8618 7855 8624 7867
rect 7603 7824 7661 7830
rect 7603 7790 7615 7824
rect 7649 7821 7661 7824
rect 7792 7821 7798 7833
rect 7649 7793 7798 7821
rect 7649 7790 7661 7793
rect 7603 7784 7661 7790
rect 7792 7781 7798 7793
rect 7850 7781 7856 7833
rect 8755 7824 8813 7830
rect 8755 7790 8767 7824
rect 8801 7821 8813 7824
rect 11248 7821 11254 7833
rect 8801 7793 11254 7821
rect 8801 7790 8813 7793
rect 8755 7784 8813 7790
rect 11248 7781 11254 7793
rect 11306 7781 11312 7833
rect 12946 7821 12974 7867
rect 22096 7855 22102 7907
rect 22154 7895 22160 7907
rect 22154 7867 27374 7895
rect 22154 7855 22160 7867
rect 17104 7821 17110 7833
rect 12946 7793 17110 7821
rect 17104 7781 17110 7793
rect 17162 7781 17168 7833
rect 24304 7821 24310 7833
rect 24265 7793 24310 7821
rect 24304 7781 24310 7793
rect 24362 7821 24368 7833
rect 25072 7821 25078 7833
rect 24362 7793 24638 7821
rect 25033 7793 25078 7821
rect 24362 7781 24368 7793
rect 3283 7750 3341 7756
rect 3283 7716 3295 7750
rect 3329 7716 3341 7750
rect 4048 7747 4054 7759
rect 4009 7719 4054 7747
rect 3283 7710 3341 7716
rect 4048 7707 4054 7719
rect 4106 7707 4112 7759
rect 4819 7750 4877 7756
rect 4819 7716 4831 7750
rect 4865 7747 4877 7750
rect 4912 7747 4918 7759
rect 4865 7719 4918 7747
rect 4865 7716 4877 7719
rect 4819 7710 4877 7716
rect 4912 7707 4918 7719
rect 4970 7707 4976 7759
rect 5299 7750 5357 7756
rect 5299 7716 5311 7750
rect 5345 7747 5357 7750
rect 5584 7747 5590 7759
rect 5345 7719 5590 7747
rect 5345 7716 5357 7719
rect 5299 7710 5357 7716
rect 5584 7707 5590 7719
rect 5642 7707 5648 7759
rect 7936 7707 7942 7759
rect 7994 7707 8000 7759
rect 10192 7747 10198 7759
rect 8386 7719 8544 7747
rect 10153 7719 10198 7747
rect 1456 7633 1462 7685
rect 1514 7673 1520 7685
rect 8386 7682 8414 7719
rect 10192 7707 10198 7719
rect 10250 7707 10256 7759
rect 10960 7747 10966 7759
rect 10921 7719 10966 7747
rect 10960 7707 10966 7719
rect 11018 7707 11024 7759
rect 12400 7747 12406 7759
rect 12361 7719 12406 7747
rect 12400 7707 12406 7719
rect 12458 7707 12464 7759
rect 12496 7707 12502 7759
rect 12554 7747 12560 7759
rect 13843 7750 13901 7756
rect 13843 7747 13855 7750
rect 12554 7719 13855 7747
rect 12554 7707 12560 7719
rect 13843 7716 13855 7719
rect 13889 7716 13901 7750
rect 13843 7710 13901 7716
rect 15571 7750 15629 7756
rect 15571 7716 15583 7750
rect 15617 7747 15629 7750
rect 15859 7750 15917 7756
rect 15859 7747 15871 7750
rect 15617 7719 15871 7747
rect 15617 7716 15629 7719
rect 15571 7710 15629 7716
rect 15859 7716 15871 7719
rect 15905 7747 15917 7750
rect 15952 7747 15958 7759
rect 15905 7719 15958 7747
rect 15905 7716 15917 7719
rect 15859 7710 15917 7716
rect 15952 7707 15958 7719
rect 16010 7707 16016 7759
rect 20944 7747 20950 7759
rect 20905 7719 20950 7747
rect 20944 7707 20950 7719
rect 21002 7707 21008 7759
rect 23635 7750 23693 7756
rect 23635 7716 23647 7750
rect 23681 7747 23693 7750
rect 23920 7747 23926 7759
rect 23681 7719 23926 7747
rect 23681 7716 23693 7719
rect 23635 7710 23693 7716
rect 23920 7707 23926 7719
rect 23978 7707 23984 7759
rect 24610 7756 24638 7793
rect 25072 7781 25078 7793
rect 25130 7821 25136 7833
rect 27346 7821 27374 7867
rect 28912 7855 28918 7907
rect 28970 7895 28976 7907
rect 29011 7898 29069 7904
rect 29011 7895 29023 7898
rect 28970 7867 29023 7895
rect 28970 7855 28976 7867
rect 29011 7864 29023 7867
rect 29057 7864 29069 7898
rect 36496 7895 36502 7907
rect 36457 7867 36502 7895
rect 29011 7858 29069 7864
rect 36496 7855 36502 7867
rect 36554 7855 36560 7907
rect 39088 7855 39094 7907
rect 39146 7895 39152 7907
rect 39187 7898 39245 7904
rect 39187 7895 39199 7898
rect 39146 7867 39199 7895
rect 39146 7855 39152 7867
rect 39187 7864 39199 7867
rect 39233 7864 39245 7898
rect 39187 7858 39245 7864
rect 40051 7898 40109 7904
rect 40051 7864 40063 7898
rect 40097 7895 40109 7898
rect 40240 7895 40246 7907
rect 40097 7867 40246 7895
rect 40097 7864 40109 7867
rect 40051 7858 40109 7864
rect 40240 7855 40246 7867
rect 40298 7855 40304 7907
rect 44752 7895 44758 7907
rect 40354 7867 44758 7895
rect 37456 7821 37462 7833
rect 25130 7793 25502 7821
rect 27346 7793 37462 7821
rect 25130 7781 25136 7793
rect 24595 7750 24653 7756
rect 24595 7716 24607 7750
rect 24641 7716 24653 7750
rect 24595 7710 24653 7716
rect 24784 7707 24790 7759
rect 24842 7747 24848 7759
rect 25474 7756 25502 7793
rect 37456 7781 37462 7793
rect 37514 7781 37520 7833
rect 40354 7821 40382 7867
rect 44752 7855 44758 7867
rect 44810 7855 44816 7907
rect 46099 7898 46157 7904
rect 46099 7864 46111 7898
rect 46145 7895 46157 7898
rect 51184 7895 51190 7907
rect 46145 7867 51190 7895
rect 46145 7864 46157 7867
rect 46099 7858 46157 7864
rect 38722 7793 40382 7821
rect 25363 7750 25421 7756
rect 25363 7747 25375 7750
rect 24842 7719 25375 7747
rect 24842 7707 24848 7719
rect 25363 7716 25375 7719
rect 25409 7716 25421 7750
rect 25363 7710 25421 7716
rect 25459 7750 25517 7756
rect 25459 7716 25471 7750
rect 25505 7716 25517 7750
rect 25459 7710 25517 7716
rect 25939 7750 25997 7756
rect 25939 7716 25951 7750
rect 25985 7747 25997 7750
rect 26128 7747 26134 7759
rect 25985 7719 26134 7747
rect 25985 7716 25997 7719
rect 25939 7710 25997 7716
rect 26128 7707 26134 7719
rect 26186 7707 26192 7759
rect 28912 7707 28918 7759
rect 28970 7747 28976 7759
rect 29299 7750 29357 7756
rect 29299 7747 29311 7750
rect 28970 7719 29311 7747
rect 28970 7707 28976 7719
rect 29299 7716 29311 7719
rect 29345 7716 29357 7750
rect 30160 7747 30166 7759
rect 30121 7719 30166 7747
rect 29299 7710 29357 7716
rect 30160 7707 30166 7719
rect 30218 7707 30224 7759
rect 33808 7747 33814 7759
rect 33769 7719 33814 7747
rect 33808 7707 33814 7719
rect 33866 7707 33872 7759
rect 34576 7747 34582 7759
rect 34537 7719 34582 7747
rect 34576 7707 34582 7719
rect 34634 7707 34640 7759
rect 35344 7747 35350 7759
rect 35305 7719 35350 7747
rect 35344 7707 35350 7719
rect 35402 7707 35408 7759
rect 36112 7747 36118 7759
rect 36073 7719 36118 7747
rect 36112 7707 36118 7719
rect 36170 7707 36176 7759
rect 36496 7707 36502 7759
rect 36554 7747 36560 7759
rect 36787 7750 36845 7756
rect 36787 7747 36799 7750
rect 36554 7719 36799 7747
rect 36554 7707 36560 7719
rect 36787 7716 36799 7719
rect 36833 7716 36845 7750
rect 38722 7747 38750 7793
rect 36787 7710 36845 7716
rect 37426 7719 38750 7747
rect 1555 7676 1613 7682
rect 1555 7673 1567 7676
rect 1514 7645 1567 7673
rect 1514 7633 1520 7645
rect 1555 7642 1567 7645
rect 1601 7642 1613 7676
rect 1555 7636 1613 7642
rect 8371 7676 8429 7682
rect 8371 7642 8383 7676
rect 8417 7642 8429 7676
rect 9424 7673 9430 7685
rect 9385 7645 9430 7673
rect 8371 7636 8429 7642
rect 9424 7633 9430 7645
rect 9482 7633 9488 7685
rect 12883 7676 12941 7682
rect 12883 7642 12895 7676
rect 12929 7673 12941 7676
rect 13171 7676 13229 7682
rect 13171 7673 13183 7676
rect 12929 7645 13183 7673
rect 12929 7642 12941 7645
rect 12883 7636 12941 7642
rect 13171 7642 13183 7645
rect 13217 7673 13229 7676
rect 28339 7676 28397 7682
rect 13217 7645 27374 7673
rect 13217 7642 13229 7645
rect 13171 7636 13229 7642
rect 8230 7611 8282 7617
rect 7024 7559 7030 7611
rect 7082 7599 7088 7611
rect 7123 7602 7181 7608
rect 7123 7599 7135 7602
rect 7082 7571 7135 7599
rect 7082 7559 7088 7571
rect 7123 7568 7135 7571
rect 7169 7568 7181 7602
rect 7123 7562 7181 7568
rect 13939 7602 13997 7608
rect 13939 7568 13951 7602
rect 13985 7599 13997 7602
rect 14224 7599 14230 7611
rect 13985 7571 14230 7599
rect 13985 7568 13997 7571
rect 13939 7562 13997 7568
rect 14224 7559 14230 7571
rect 14282 7559 14288 7611
rect 15187 7602 15245 7608
rect 15187 7568 15199 7602
rect 15233 7568 15245 7602
rect 15187 7562 15245 7568
rect 8230 7553 8282 7559
rect 9136 7485 9142 7537
rect 9194 7525 9200 7537
rect 10115 7528 10173 7534
rect 10115 7525 10127 7528
rect 9194 7497 10127 7525
rect 9194 7485 9200 7497
rect 10115 7494 10127 7497
rect 10161 7494 10173 7528
rect 10115 7488 10173 7494
rect 11728 7485 11734 7537
rect 11786 7525 11792 7537
rect 15202 7525 15230 7562
rect 15952 7559 15958 7611
rect 16010 7599 16016 7611
rect 21715 7602 21773 7608
rect 21715 7599 21727 7602
rect 16010 7571 21727 7599
rect 16010 7559 16016 7571
rect 21715 7568 21727 7571
rect 21761 7568 21773 7602
rect 21715 7562 21773 7568
rect 23251 7602 23309 7608
rect 23251 7568 23263 7602
rect 23297 7568 23309 7602
rect 23251 7562 23309 7568
rect 23152 7525 23158 7537
rect 11786 7497 13118 7525
rect 15202 7497 23158 7525
rect 11786 7485 11792 7497
rect 2416 7451 2422 7463
rect 2377 7423 2422 7451
rect 2416 7411 2422 7423
rect 2474 7411 2480 7463
rect 3187 7454 3245 7460
rect 3187 7420 3199 7454
rect 3233 7451 3245 7454
rect 3280 7451 3286 7463
rect 3233 7423 3286 7451
rect 3233 7420 3245 7423
rect 3187 7414 3245 7420
rect 3280 7411 3286 7423
rect 3338 7411 3344 7463
rect 3376 7411 3382 7463
rect 3434 7451 3440 7463
rect 3955 7454 4013 7460
rect 3955 7451 3967 7454
rect 3434 7423 3967 7451
rect 3434 7411 3440 7423
rect 3955 7420 3967 7423
rect 4001 7420 4013 7454
rect 3955 7414 4013 7420
rect 4048 7411 4054 7463
rect 4106 7451 4112 7463
rect 4723 7454 4781 7460
rect 4723 7451 4735 7454
rect 4106 7423 4735 7451
rect 4106 7411 4112 7423
rect 4723 7420 4735 7423
rect 4769 7420 4781 7454
rect 4723 7414 4781 7420
rect 5296 7411 5302 7463
rect 5354 7451 5360 7463
rect 5491 7454 5549 7460
rect 5491 7451 5503 7454
rect 5354 7423 5503 7451
rect 5354 7411 5360 7423
rect 5491 7420 5503 7423
rect 5537 7420 5549 7454
rect 5491 7414 5549 7420
rect 8752 7411 8758 7463
rect 8810 7451 8816 7463
rect 9331 7454 9389 7460
rect 9331 7451 9343 7454
rect 8810 7423 9343 7451
rect 8810 7411 8816 7423
rect 9331 7420 9343 7423
rect 9377 7420 9389 7454
rect 9331 7414 9389 7420
rect 9904 7411 9910 7463
rect 9962 7451 9968 7463
rect 10867 7454 10925 7460
rect 10867 7451 10879 7454
rect 9962 7423 10879 7451
rect 9962 7411 9968 7423
rect 10867 7420 10879 7423
rect 10913 7420 10925 7454
rect 10867 7414 10925 7420
rect 10960 7411 10966 7463
rect 11018 7451 11024 7463
rect 13090 7460 13118 7497
rect 23152 7485 23158 7497
rect 23210 7485 23216 7537
rect 23266 7525 23294 7562
rect 25456 7559 25462 7611
rect 25514 7599 25520 7611
rect 26995 7602 27053 7608
rect 26995 7599 27007 7602
rect 25514 7571 27007 7599
rect 25514 7559 25520 7571
rect 26995 7568 27007 7571
rect 27041 7568 27053 7602
rect 27346 7599 27374 7645
rect 28339 7642 28351 7676
rect 28385 7673 28397 7676
rect 37426 7673 37454 7719
rect 38800 7707 38806 7759
rect 38858 7747 38864 7759
rect 39571 7750 39629 7756
rect 39571 7747 39583 7750
rect 38858 7719 39583 7747
rect 38858 7707 38864 7719
rect 39571 7716 39583 7719
rect 39617 7716 39629 7750
rect 39571 7710 39629 7716
rect 40240 7707 40246 7759
rect 40298 7747 40304 7759
rect 41011 7750 41069 7756
rect 41011 7747 41023 7750
rect 40298 7719 41023 7747
rect 40298 7707 40304 7719
rect 41011 7716 41023 7719
rect 41057 7716 41069 7750
rect 41011 7710 41069 7716
rect 41107 7750 41165 7756
rect 41107 7716 41119 7750
rect 41153 7747 41165 7750
rect 41776 7747 41782 7759
rect 41153 7719 41782 7747
rect 41153 7716 41165 7719
rect 41107 7710 41165 7716
rect 41776 7707 41782 7719
rect 41834 7707 41840 7759
rect 42643 7750 42701 7756
rect 42643 7716 42655 7750
rect 42689 7747 42701 7750
rect 42736 7747 42742 7759
rect 42689 7719 42742 7747
rect 42689 7716 42701 7719
rect 42643 7710 42701 7716
rect 42736 7707 42742 7719
rect 42794 7707 42800 7759
rect 43984 7707 43990 7759
rect 44042 7747 44048 7759
rect 44083 7750 44141 7756
rect 44083 7747 44095 7750
rect 44042 7719 44095 7747
rect 44042 7707 44048 7719
rect 44083 7716 44095 7719
rect 44129 7716 44141 7750
rect 44083 7710 44141 7716
rect 44851 7750 44909 7756
rect 44851 7716 44863 7750
rect 44897 7747 44909 7750
rect 45040 7747 45046 7759
rect 44897 7719 45046 7747
rect 44897 7716 44909 7719
rect 44851 7710 44909 7716
rect 45040 7707 45046 7719
rect 45098 7707 45104 7759
rect 45616 7747 45622 7759
rect 45577 7719 45622 7747
rect 45616 7707 45622 7719
rect 45674 7707 45680 7759
rect 45808 7707 45814 7759
rect 45866 7747 45872 7759
rect 46402 7756 46430 7867
rect 51184 7855 51190 7867
rect 51242 7855 51248 7907
rect 51472 7895 51478 7907
rect 51433 7867 51478 7895
rect 51472 7855 51478 7867
rect 51530 7895 51536 7907
rect 51530 7867 51806 7895
rect 51530 7855 51536 7867
rect 51664 7821 51670 7833
rect 47170 7793 51670 7821
rect 46291 7750 46349 7756
rect 46291 7747 46303 7750
rect 45866 7719 46303 7747
rect 45866 7707 45872 7719
rect 46291 7716 46303 7719
rect 46337 7716 46349 7750
rect 46291 7710 46349 7716
rect 46387 7750 46445 7756
rect 46387 7716 46399 7750
rect 46433 7716 46445 7750
rect 46387 7710 46445 7716
rect 46480 7707 46486 7759
rect 46538 7747 46544 7759
rect 47059 7750 47117 7756
rect 47059 7747 47071 7750
rect 46538 7719 47071 7747
rect 46538 7707 46544 7719
rect 47059 7716 47071 7719
rect 47105 7716 47117 7750
rect 47059 7710 47117 7716
rect 28385 7645 37454 7673
rect 28385 7642 28397 7645
rect 28339 7636 28397 7642
rect 39088 7633 39094 7685
rect 39146 7673 39152 7685
rect 39475 7676 39533 7682
rect 39475 7673 39487 7676
rect 39146 7645 39487 7673
rect 39146 7633 39152 7645
rect 39475 7642 39487 7645
rect 39521 7642 39533 7676
rect 43888 7673 43894 7685
rect 39475 7636 39533 7642
rect 40066 7645 43894 7673
rect 27346 7571 30302 7599
rect 26995 7562 27053 7568
rect 30160 7525 30166 7537
rect 23266 7497 30166 7525
rect 30160 7485 30166 7497
rect 30218 7485 30224 7537
rect 30274 7525 30302 7571
rect 30640 7559 30646 7611
rect 30698 7599 30704 7611
rect 31219 7602 31277 7608
rect 31219 7599 31231 7602
rect 30698 7571 31231 7599
rect 30698 7559 30704 7571
rect 31219 7568 31231 7571
rect 31265 7568 31277 7602
rect 32368 7599 32374 7611
rect 32329 7571 32374 7599
rect 31219 7562 31277 7568
rect 32368 7559 32374 7571
rect 32426 7559 32432 7611
rect 38803 7602 38861 7608
rect 38803 7568 38815 7602
rect 38849 7599 38861 7602
rect 40066 7599 40094 7645
rect 43888 7633 43894 7645
rect 43946 7633 43952 7685
rect 47170 7673 47198 7793
rect 51664 7781 51670 7793
rect 51722 7781 51728 7833
rect 49360 7747 49366 7759
rect 49321 7719 49366 7747
rect 49360 7707 49366 7719
rect 49418 7707 49424 7759
rect 50131 7750 50189 7756
rect 50131 7716 50143 7750
rect 50177 7747 50189 7750
rect 50992 7747 50998 7759
rect 50177 7719 50998 7747
rect 50177 7716 50189 7719
rect 50131 7710 50189 7716
rect 50992 7707 50998 7719
rect 51050 7707 51056 7759
rect 51778 7756 51806 7867
rect 51763 7750 51821 7756
rect 51763 7716 51775 7750
rect 51809 7716 51821 7750
rect 52624 7747 52630 7759
rect 52585 7719 52630 7747
rect 51763 7710 51821 7716
rect 52624 7707 52630 7719
rect 52682 7707 52688 7759
rect 53392 7747 53398 7759
rect 53353 7719 53398 7747
rect 53392 7707 53398 7719
rect 53450 7707 53456 7759
rect 58768 7747 58774 7759
rect 55138 7719 58774 7747
rect 52528 7673 52534 7685
rect 44674 7645 47198 7673
rect 47506 7645 52534 7673
rect 38849 7571 40094 7599
rect 38849 7568 38861 7571
rect 38803 7562 38861 7568
rect 40144 7559 40150 7611
rect 40202 7599 40208 7611
rect 40243 7602 40301 7608
rect 40243 7599 40255 7602
rect 40202 7571 40255 7599
rect 40202 7559 40208 7571
rect 40243 7568 40255 7571
rect 40289 7568 40301 7602
rect 40243 7562 40301 7568
rect 41875 7602 41933 7608
rect 41875 7568 41887 7602
rect 41921 7599 41933 7602
rect 44674 7599 44702 7645
rect 41921 7571 44702 7599
rect 46867 7602 46925 7608
rect 41921 7568 41933 7571
rect 41875 7562 41933 7568
rect 46867 7568 46879 7602
rect 46913 7599 46925 7602
rect 47155 7602 47213 7608
rect 47155 7599 47167 7602
rect 46913 7571 47167 7599
rect 46913 7568 46925 7571
rect 46867 7562 46925 7568
rect 47155 7568 47167 7571
rect 47201 7599 47213 7602
rect 47506 7599 47534 7645
rect 52528 7633 52534 7645
rect 52586 7633 52592 7685
rect 55138 7682 55166 7719
rect 58768 7707 58774 7719
rect 58826 7707 58832 7759
rect 55123 7676 55181 7682
rect 55123 7642 55135 7676
rect 55169 7642 55181 7676
rect 55792 7673 55798 7685
rect 55753 7645 55798 7673
rect 55123 7636 55181 7642
rect 55792 7633 55798 7645
rect 55850 7633 55856 7685
rect 56176 7633 56182 7685
rect 56234 7673 56240 7685
rect 56563 7676 56621 7682
rect 56563 7673 56575 7676
rect 56234 7645 56575 7673
rect 56234 7633 56240 7645
rect 56563 7642 56575 7645
rect 56609 7642 56621 7676
rect 56563 7636 56621 7642
rect 56656 7633 56662 7685
rect 56714 7673 56720 7685
rect 57331 7676 57389 7682
rect 57331 7673 57343 7676
rect 56714 7645 57343 7673
rect 56714 7633 56720 7645
rect 57331 7642 57343 7645
rect 57377 7642 57389 7676
rect 57331 7636 57389 7642
rect 47920 7599 47926 7611
rect 47201 7571 47534 7599
rect 47881 7571 47926 7599
rect 47201 7568 47213 7571
rect 47155 7562 47213 7568
rect 47920 7559 47926 7571
rect 47978 7559 47984 7611
rect 51091 7602 51149 7608
rect 51091 7568 51103 7602
rect 51137 7599 51149 7602
rect 57136 7599 57142 7611
rect 51137 7571 57142 7599
rect 51137 7568 51149 7571
rect 51091 7562 51149 7568
rect 57136 7559 57142 7571
rect 57194 7559 57200 7611
rect 48112 7525 48118 7537
rect 30274 7497 48118 7525
rect 48112 7485 48118 7497
rect 48170 7485 48176 7537
rect 49168 7485 49174 7537
rect 49226 7525 49232 7537
rect 59344 7525 59350 7537
rect 49226 7497 50078 7525
rect 49226 7485 49232 7497
rect 12307 7454 12365 7460
rect 12307 7451 12319 7454
rect 11018 7423 12319 7451
rect 11018 7411 11024 7423
rect 12307 7420 12319 7423
rect 12353 7420 12365 7454
rect 12307 7414 12365 7420
rect 13075 7454 13133 7460
rect 13075 7420 13087 7454
rect 13121 7420 13133 7454
rect 13075 7414 13133 7420
rect 15664 7411 15670 7463
rect 15722 7451 15728 7463
rect 15763 7454 15821 7460
rect 15763 7451 15775 7454
rect 15722 7423 15775 7451
rect 15722 7411 15728 7423
rect 15763 7420 15775 7423
rect 15809 7420 15821 7454
rect 15763 7414 15821 7420
rect 20752 7411 20758 7463
rect 20810 7451 20816 7463
rect 20851 7454 20909 7460
rect 20851 7451 20863 7454
rect 20810 7423 20863 7451
rect 20810 7411 20816 7423
rect 20851 7420 20863 7423
rect 20897 7420 20909 7454
rect 20851 7414 20909 7420
rect 23728 7411 23734 7463
rect 23786 7451 23792 7463
rect 23827 7454 23885 7460
rect 23827 7451 23839 7454
rect 23786 7423 23839 7451
rect 23786 7411 23792 7423
rect 23827 7420 23839 7423
rect 23873 7420 23885 7454
rect 24688 7451 24694 7463
rect 24649 7423 24694 7451
rect 23827 7414 23885 7420
rect 24688 7411 24694 7423
rect 24746 7411 24752 7463
rect 25936 7411 25942 7463
rect 25994 7451 26000 7463
rect 26227 7454 26285 7460
rect 26227 7451 26239 7454
rect 25994 7423 26239 7451
rect 25994 7411 26000 7423
rect 26227 7420 26239 7423
rect 26273 7420 26285 7454
rect 26227 7414 26285 7420
rect 26704 7411 26710 7463
rect 26762 7451 26768 7463
rect 26899 7454 26957 7460
rect 26899 7451 26911 7454
rect 26762 7423 26911 7451
rect 26762 7411 26768 7423
rect 26899 7420 26911 7423
rect 26945 7420 26957 7454
rect 26899 7414 26957 7420
rect 28144 7411 28150 7463
rect 28202 7451 28208 7463
rect 28243 7454 28301 7460
rect 28243 7451 28255 7454
rect 28202 7423 28255 7451
rect 28202 7411 28208 7423
rect 28243 7420 28255 7423
rect 28289 7420 28301 7454
rect 28243 7414 28301 7420
rect 29200 7411 29206 7463
rect 29258 7451 29264 7463
rect 29395 7454 29453 7460
rect 29395 7451 29407 7454
rect 29258 7423 29407 7451
rect 29258 7411 29264 7423
rect 29395 7420 29407 7423
rect 29441 7420 29453 7454
rect 29395 7414 29453 7420
rect 29584 7411 29590 7463
rect 29642 7451 29648 7463
rect 30067 7454 30125 7460
rect 30067 7451 30079 7454
rect 29642 7423 30079 7451
rect 29642 7411 29648 7423
rect 30067 7420 30079 7423
rect 30113 7420 30125 7454
rect 30067 7414 30125 7420
rect 31024 7411 31030 7463
rect 31082 7451 31088 7463
rect 31123 7454 31181 7460
rect 31123 7451 31135 7454
rect 31082 7423 31135 7451
rect 31082 7411 31088 7423
rect 31123 7420 31135 7423
rect 31169 7420 31181 7454
rect 31123 7414 31181 7420
rect 33616 7411 33622 7463
rect 33674 7451 33680 7463
rect 33715 7454 33773 7460
rect 33715 7451 33727 7454
rect 33674 7423 33727 7451
rect 33674 7411 33680 7423
rect 33715 7420 33727 7423
rect 33761 7420 33773 7454
rect 33715 7414 33773 7420
rect 34384 7411 34390 7463
rect 34442 7451 34448 7463
rect 34483 7454 34541 7460
rect 34483 7451 34495 7454
rect 34442 7423 34495 7451
rect 34442 7411 34448 7423
rect 34483 7420 34495 7423
rect 34529 7420 34541 7454
rect 34483 7414 34541 7420
rect 34768 7411 34774 7463
rect 34826 7451 34832 7463
rect 35251 7454 35309 7460
rect 35251 7451 35263 7454
rect 34826 7423 35263 7451
rect 34826 7411 34832 7423
rect 35251 7420 35263 7423
rect 35297 7420 35309 7454
rect 35251 7414 35309 7420
rect 35824 7411 35830 7463
rect 35882 7451 35888 7463
rect 36019 7454 36077 7460
rect 36019 7451 36031 7454
rect 35882 7423 36031 7451
rect 35882 7411 35888 7423
rect 36019 7420 36031 7423
rect 36065 7420 36077 7454
rect 36019 7414 36077 7420
rect 36592 7411 36598 7463
rect 36650 7451 36656 7463
rect 36883 7454 36941 7460
rect 36883 7451 36895 7454
rect 36650 7423 36895 7451
rect 36650 7411 36656 7423
rect 36883 7420 36895 7423
rect 36929 7420 36941 7454
rect 36883 7414 36941 7420
rect 38032 7411 38038 7463
rect 38090 7451 38096 7463
rect 38707 7454 38765 7460
rect 38707 7451 38719 7454
rect 38090 7423 38719 7451
rect 38090 7411 38096 7423
rect 38707 7420 38719 7423
rect 38753 7420 38765 7454
rect 38707 7414 38765 7420
rect 39472 7411 39478 7463
rect 39530 7451 39536 7463
rect 40339 7454 40397 7460
rect 40339 7451 40351 7454
rect 39530 7423 40351 7451
rect 39530 7411 39536 7423
rect 40339 7420 40351 7423
rect 40385 7420 40397 7454
rect 41776 7451 41782 7463
rect 41737 7423 41782 7451
rect 40339 7414 40397 7420
rect 41776 7411 41782 7423
rect 41834 7411 41840 7463
rect 42448 7411 42454 7463
rect 42506 7451 42512 7463
rect 42547 7454 42605 7460
rect 42547 7451 42559 7454
rect 42506 7423 42559 7451
rect 42506 7411 42512 7423
rect 42547 7420 42559 7423
rect 42593 7420 42605 7454
rect 42547 7414 42605 7420
rect 43888 7411 43894 7463
rect 43946 7451 43952 7463
rect 43987 7454 44045 7460
rect 43987 7451 43999 7454
rect 43946 7423 43999 7451
rect 43946 7411 43952 7423
rect 43987 7420 43999 7423
rect 44033 7420 44045 7454
rect 44752 7451 44758 7463
rect 44713 7423 44758 7451
rect 43987 7414 44045 7420
rect 44752 7411 44758 7423
rect 44810 7411 44816 7463
rect 45040 7411 45046 7463
rect 45098 7451 45104 7463
rect 45523 7454 45581 7460
rect 45523 7451 45535 7454
rect 45098 7423 45535 7451
rect 45098 7411 45104 7423
rect 45523 7420 45535 7423
rect 45569 7420 45581 7454
rect 45523 7414 45581 7420
rect 47248 7411 47254 7463
rect 47306 7451 47312 7463
rect 47827 7454 47885 7460
rect 47827 7451 47839 7454
rect 47306 7423 47839 7451
rect 47306 7411 47312 7423
rect 47827 7420 47839 7423
rect 47873 7420 47885 7454
rect 47827 7414 47885 7420
rect 48400 7411 48406 7463
rect 48458 7451 48464 7463
rect 50050 7460 50078 7497
rect 51010 7497 59350 7525
rect 51010 7460 51038 7497
rect 59344 7485 59350 7497
rect 59402 7485 59408 7537
rect 49267 7454 49325 7460
rect 49267 7451 49279 7454
rect 48458 7423 49279 7451
rect 48458 7411 48464 7423
rect 49267 7420 49279 7423
rect 49313 7420 49325 7454
rect 49267 7414 49325 7420
rect 50035 7454 50093 7460
rect 50035 7420 50047 7454
rect 50081 7420 50093 7454
rect 50035 7414 50093 7420
rect 50995 7454 51053 7460
rect 50995 7420 51007 7454
rect 51041 7420 51053 7454
rect 50995 7414 51053 7420
rect 51664 7411 51670 7463
rect 51722 7451 51728 7463
rect 51859 7454 51917 7460
rect 51859 7451 51871 7454
rect 51722 7423 51871 7451
rect 51722 7411 51728 7423
rect 51859 7420 51871 7423
rect 51905 7420 51917 7454
rect 51859 7414 51917 7420
rect 52336 7411 52342 7463
rect 52394 7451 52400 7463
rect 52531 7454 52589 7460
rect 52531 7451 52543 7454
rect 52394 7423 52543 7451
rect 52394 7411 52400 7423
rect 52531 7420 52543 7423
rect 52577 7420 52589 7454
rect 52531 7414 52589 7420
rect 52720 7411 52726 7463
rect 52778 7451 52784 7463
rect 53299 7454 53357 7460
rect 53299 7451 53311 7454
rect 52778 7423 53311 7451
rect 52778 7411 52784 7423
rect 53299 7420 53311 7423
rect 53345 7420 53357 7454
rect 53299 7414 53357 7420
rect 1152 7352 58848 7374
rect 1152 7300 19654 7352
rect 19706 7300 19718 7352
rect 19770 7300 19782 7352
rect 19834 7300 19846 7352
rect 19898 7300 50374 7352
rect 50426 7300 50438 7352
rect 50490 7300 50502 7352
rect 50554 7300 50566 7352
rect 50618 7300 58848 7352
rect 1152 7278 58848 7300
rect 1840 7189 1846 7241
rect 1898 7229 1904 7241
rect 7792 7229 7798 7241
rect 1898 7201 7798 7229
rect 1898 7189 1904 7201
rect 7792 7189 7798 7201
rect 7850 7189 7856 7241
rect 32368 7189 32374 7241
rect 32426 7229 32432 7241
rect 47920 7229 47926 7241
rect 32426 7201 47926 7229
rect 32426 7189 32432 7201
rect 47920 7189 47926 7201
rect 47978 7189 47984 7241
rect 17779 7158 17837 7164
rect 4546 7127 17726 7155
rect 4546 7090 4574 7127
rect 4243 7084 4301 7090
rect 4243 7050 4255 7084
rect 4289 7081 4301 7084
rect 4531 7084 4589 7090
rect 4531 7081 4543 7084
rect 4289 7053 4543 7081
rect 4289 7050 4301 7053
rect 4243 7044 4301 7050
rect 4531 7050 4543 7053
rect 4577 7050 4589 7084
rect 4531 7044 4589 7050
rect 6547 7084 6605 7090
rect 6547 7050 6559 7084
rect 6593 7081 6605 7084
rect 6832 7081 6838 7093
rect 6593 7053 6838 7081
rect 6593 7050 6605 7053
rect 6547 7044 6605 7050
rect 6832 7041 6838 7053
rect 6890 7041 6896 7093
rect 7600 7081 7606 7093
rect 7561 7053 7606 7081
rect 7600 7041 7606 7053
rect 7658 7041 7664 7093
rect 8368 7081 8374 7093
rect 8329 7053 8374 7081
rect 8368 7041 8374 7053
rect 8426 7041 8432 7093
rect 9811 7084 9869 7090
rect 9811 7050 9823 7084
rect 9857 7081 9869 7084
rect 10000 7081 10006 7093
rect 9857 7053 10006 7081
rect 9857 7050 9869 7053
rect 9811 7044 9869 7050
rect 10000 7041 10006 7053
rect 10058 7041 10064 7093
rect 10291 7084 10349 7090
rect 10291 7050 10303 7084
rect 10337 7081 10349 7084
rect 10579 7084 10637 7090
rect 10579 7081 10591 7084
rect 10337 7053 10591 7081
rect 10337 7050 10349 7053
rect 10291 7044 10349 7050
rect 10579 7050 10591 7053
rect 10625 7081 10637 7084
rect 10864 7081 10870 7093
rect 10625 7053 10870 7081
rect 10625 7050 10637 7053
rect 10579 7044 10637 7050
rect 10864 7041 10870 7053
rect 10922 7041 10928 7093
rect 13456 7041 13462 7093
rect 13514 7081 13520 7093
rect 13651 7084 13709 7090
rect 13651 7081 13663 7084
rect 13514 7053 13663 7081
rect 13514 7041 13520 7053
rect 13651 7050 13663 7053
rect 13697 7050 13709 7084
rect 13651 7044 13709 7050
rect 14803 7084 14861 7090
rect 14803 7050 14815 7084
rect 14849 7081 14861 7084
rect 14992 7081 14998 7093
rect 14849 7053 14998 7081
rect 14849 7050 14861 7053
rect 14803 7044 14861 7050
rect 14992 7041 14998 7053
rect 15050 7041 15056 7093
rect 15859 7084 15917 7090
rect 15859 7050 15871 7084
rect 15905 7081 15917 7084
rect 16048 7081 16054 7093
rect 15905 7053 16054 7081
rect 15905 7050 15917 7053
rect 15859 7044 15917 7050
rect 16048 7041 16054 7053
rect 16106 7041 16112 7093
rect 16339 7084 16397 7090
rect 16339 7050 16351 7084
rect 16385 7081 16397 7084
rect 16624 7081 16630 7093
rect 16385 7053 16630 7081
rect 16385 7050 16397 7053
rect 16339 7044 16397 7050
rect 16624 7041 16630 7053
rect 16682 7041 16688 7093
rect 17296 7041 17302 7093
rect 17354 7081 17360 7093
rect 17354 7053 17399 7081
rect 17354 7041 17360 7053
rect 1648 7007 1654 7019
rect 1609 6979 1654 7007
rect 1648 6967 1654 6979
rect 1706 6967 1712 7019
rect 2512 7007 2518 7019
rect 2473 6979 2518 7007
rect 2512 6967 2518 6979
rect 2570 6967 2576 7019
rect 3664 6967 3670 7019
rect 3722 7007 3728 7019
rect 6067 7010 6125 7016
rect 3722 6979 5246 7007
rect 3722 6967 3728 6979
rect 5218 6942 5246 6979
rect 6067 6976 6079 7010
rect 6113 7007 6125 7010
rect 11248 7007 11254 7019
rect 6113 6979 11006 7007
rect 11209 6979 11254 7007
rect 6113 6976 6125 6979
rect 6067 6970 6125 6976
rect 4435 6936 4493 6942
rect 4435 6902 4447 6936
rect 4481 6902 4493 6936
rect 4435 6896 4493 6902
rect 5203 6936 5261 6942
rect 5203 6902 5215 6936
rect 5249 6902 5261 6936
rect 5203 6896 5261 6902
rect 5299 6936 5357 6942
rect 5299 6902 5311 6936
rect 5345 6933 5357 6936
rect 5776 6933 5782 6945
rect 5345 6905 5782 6933
rect 5345 6902 5357 6905
rect 5299 6896 5357 6902
rect 4450 6785 4478 6896
rect 5776 6893 5782 6905
rect 5834 6893 5840 6945
rect 5872 6893 5878 6945
rect 5930 6933 5936 6945
rect 5971 6936 6029 6942
rect 5971 6933 5983 6936
rect 5930 6905 5983 6933
rect 5930 6893 5936 6905
rect 5971 6902 5983 6905
rect 6017 6902 6029 6936
rect 5971 6896 6029 6902
rect 6544 6893 6550 6945
rect 6602 6933 6608 6945
rect 6739 6936 6797 6942
rect 6739 6933 6751 6936
rect 6602 6905 6751 6933
rect 6602 6893 6608 6905
rect 6739 6902 6751 6905
rect 6785 6902 6797 6936
rect 6739 6896 6797 6902
rect 6928 6893 6934 6945
rect 6986 6933 6992 6945
rect 7507 6936 7565 6942
rect 7507 6933 7519 6936
rect 6986 6905 7519 6933
rect 6986 6893 6992 6905
rect 7507 6902 7519 6905
rect 7553 6902 7565 6936
rect 7507 6896 7565 6902
rect 8275 6936 8333 6942
rect 8275 6902 8287 6936
rect 8321 6902 8333 6936
rect 8275 6896 8333 6902
rect 9715 6936 9773 6942
rect 9715 6902 9727 6936
rect 9761 6902 9773 6936
rect 9715 6896 9773 6902
rect 7312 6819 7318 6871
rect 7370 6859 7376 6871
rect 8290 6859 8318 6896
rect 7370 6831 8318 6859
rect 7370 6819 7376 6831
rect 5200 6785 5206 6797
rect 4450 6757 5206 6785
rect 5200 6745 5206 6757
rect 5258 6745 5264 6797
rect 8176 6745 8182 6797
rect 8234 6785 8240 6797
rect 9730 6785 9758 6896
rect 9808 6893 9814 6945
rect 9866 6933 9872 6945
rect 10483 6936 10541 6942
rect 10483 6933 10495 6936
rect 9866 6905 10495 6933
rect 9866 6893 9872 6905
rect 10483 6902 10495 6905
rect 10529 6902 10541 6936
rect 10978 6933 11006 6979
rect 11248 6967 11254 6979
rect 11306 6967 11312 7019
rect 12688 7007 12694 7019
rect 12649 6979 12694 7007
rect 12688 6967 12694 6979
rect 12746 6967 12752 7019
rect 15952 7007 15958 7019
rect 12946 6979 15958 7007
rect 12946 6933 12974 6979
rect 15952 6967 15958 6979
rect 16010 6967 16016 7019
rect 17698 7007 17726 7127
rect 17779 7124 17791 7158
rect 17825 7155 17837 7158
rect 17872 7155 17878 7167
rect 17825 7127 17878 7155
rect 17825 7124 17837 7127
rect 17779 7118 17837 7124
rect 17872 7115 17878 7127
rect 17930 7155 17936 7167
rect 19984 7155 19990 7167
rect 17930 7127 18110 7155
rect 19945 7127 19990 7155
rect 17930 7115 17936 7127
rect 18082 7090 18110 7127
rect 19984 7115 19990 7127
rect 20042 7155 20048 7167
rect 22288 7155 22294 7167
rect 20042 7127 20318 7155
rect 22249 7127 22294 7155
rect 20042 7115 20048 7127
rect 18067 7084 18125 7090
rect 18067 7050 18079 7084
rect 18113 7050 18125 7084
rect 18832 7081 18838 7093
rect 18793 7053 18838 7081
rect 18067 7044 18125 7050
rect 18832 7041 18838 7053
rect 18890 7041 18896 7093
rect 20290 7090 20318 7127
rect 22288 7115 22294 7127
rect 22346 7155 22352 7167
rect 23155 7158 23213 7164
rect 22346 7127 22718 7155
rect 22346 7115 22352 7127
rect 20275 7084 20333 7090
rect 20275 7050 20287 7084
rect 20321 7050 20333 7084
rect 20275 7044 20333 7050
rect 21139 7084 21197 7090
rect 21139 7050 21151 7084
rect 21185 7081 21197 7084
rect 21232 7081 21238 7093
rect 21185 7053 21238 7081
rect 21185 7050 21197 7053
rect 21139 7044 21197 7050
rect 21232 7041 21238 7053
rect 21290 7041 21296 7093
rect 21619 7084 21677 7090
rect 21619 7050 21631 7084
rect 21665 7081 21677 7084
rect 21904 7081 21910 7093
rect 21665 7053 21910 7081
rect 21665 7050 21677 7053
rect 21619 7044 21677 7050
rect 21904 7041 21910 7053
rect 21962 7041 21968 7093
rect 22690 7090 22718 7127
rect 23155 7124 23167 7158
rect 23201 7155 23213 7158
rect 23248 7155 23254 7167
rect 23201 7127 23254 7155
rect 23201 7124 23213 7127
rect 23155 7118 23213 7124
rect 23248 7115 23254 7127
rect 23306 7155 23312 7167
rect 23824 7155 23830 7167
rect 23306 7127 23390 7155
rect 23785 7127 23830 7155
rect 23306 7115 23312 7127
rect 23362 7090 23390 7127
rect 23824 7115 23830 7127
rect 23882 7155 23888 7167
rect 26032 7155 26038 7167
rect 23882 7127 24158 7155
rect 25993 7127 26038 7155
rect 23882 7115 23888 7127
rect 24130 7090 24158 7127
rect 26032 7115 26038 7127
rect 26090 7155 26096 7167
rect 26800 7155 26806 7167
rect 26090 7127 26462 7155
rect 26761 7127 26806 7155
rect 26090 7115 26096 7127
rect 22675 7084 22733 7090
rect 22675 7050 22687 7084
rect 22721 7050 22733 7084
rect 22675 7044 22733 7050
rect 23347 7084 23405 7090
rect 23347 7050 23359 7084
rect 23393 7050 23405 7084
rect 23347 7044 23405 7050
rect 24115 7084 24173 7090
rect 24115 7050 24127 7084
rect 24161 7050 24173 7084
rect 24115 7044 24173 7050
rect 25363 7084 25421 7090
rect 25363 7050 25375 7084
rect 25409 7081 25421 7084
rect 25648 7081 25654 7093
rect 25409 7053 25654 7081
rect 25409 7050 25421 7053
rect 25363 7044 25421 7050
rect 25648 7041 25654 7053
rect 25706 7041 25712 7093
rect 26434 7090 26462 7127
rect 26800 7115 26806 7127
rect 26858 7155 26864 7167
rect 27568 7155 27574 7167
rect 26858 7127 27134 7155
rect 27529 7127 27574 7155
rect 26858 7115 26864 7127
rect 27106 7090 27134 7127
rect 27568 7115 27574 7127
rect 27626 7155 27632 7167
rect 30544 7155 30550 7167
rect 27626 7127 27998 7155
rect 30505 7127 30550 7155
rect 27626 7115 27632 7127
rect 27970 7090 27998 7127
rect 30544 7115 30550 7127
rect 30602 7155 30608 7167
rect 38128 7155 38134 7167
rect 30602 7127 30878 7155
rect 38089 7127 38134 7155
rect 30602 7115 30608 7127
rect 26419 7084 26477 7090
rect 26419 7050 26431 7084
rect 26465 7050 26477 7084
rect 26419 7044 26477 7050
rect 27091 7084 27149 7090
rect 27091 7050 27103 7084
rect 27137 7050 27149 7084
rect 27091 7044 27149 7050
rect 27955 7084 28013 7090
rect 27955 7050 27967 7084
rect 28001 7050 28013 7084
rect 27955 7044 28013 7050
rect 28048 7041 28054 7093
rect 28106 7081 28112 7093
rect 29488 7081 29494 7093
rect 28106 7053 29342 7081
rect 29449 7053 29494 7081
rect 28106 7041 28112 7053
rect 20656 7007 20662 7019
rect 17698 6979 20662 7007
rect 20656 6967 20662 6979
rect 20714 6967 20720 7019
rect 23152 6967 23158 7019
rect 23210 7007 23216 7019
rect 28723 7010 28781 7016
rect 28723 7007 28735 7010
rect 23210 6979 28735 7007
rect 23210 6967 23216 6979
rect 28723 6976 28735 6979
rect 28769 6976 28781 7010
rect 29314 7007 29342 7053
rect 29488 7041 29494 7053
rect 29546 7041 29552 7093
rect 30850 7090 30878 7127
rect 38128 7115 38134 7127
rect 38186 7155 38192 7167
rect 38186 7127 38462 7155
rect 38186 7115 38192 7127
rect 30835 7084 30893 7090
rect 30835 7050 30847 7084
rect 30881 7050 30893 7084
rect 30835 7044 30893 7050
rect 31411 7084 31469 7090
rect 31411 7050 31423 7084
rect 31457 7081 31469 7084
rect 31600 7081 31606 7093
rect 31457 7053 31606 7081
rect 31457 7050 31469 7053
rect 31411 7044 31469 7050
rect 31600 7041 31606 7053
rect 31658 7041 31664 7093
rect 32464 7081 32470 7093
rect 32425 7053 32470 7081
rect 32464 7041 32470 7053
rect 32522 7041 32528 7093
rect 34000 7081 34006 7093
rect 33961 7053 34006 7081
rect 34000 7041 34006 7053
rect 34058 7041 34064 7093
rect 36208 7081 36214 7093
rect 36169 7053 36214 7081
rect 36208 7041 36214 7053
rect 36266 7041 36272 7093
rect 36976 7081 36982 7093
rect 36937 7053 36982 7081
rect 36976 7041 36982 7053
rect 37034 7041 37040 7093
rect 37744 7081 37750 7093
rect 37705 7053 37750 7081
rect 37744 7041 37750 7053
rect 37802 7041 37808 7093
rect 38434 7090 38462 7127
rect 38512 7115 38518 7167
rect 38570 7155 38576 7167
rect 39475 7158 39533 7164
rect 39475 7155 39487 7158
rect 38570 7127 39487 7155
rect 38570 7115 38576 7127
rect 39475 7124 39487 7127
rect 39521 7124 39533 7158
rect 39664 7155 39670 7167
rect 39625 7127 39670 7155
rect 39475 7118 39533 7124
rect 39664 7115 39670 7127
rect 39722 7155 39728 7167
rect 41872 7155 41878 7167
rect 39722 7127 39998 7155
rect 41833 7127 41878 7155
rect 39722 7115 39728 7127
rect 39970 7090 39998 7127
rect 41872 7115 41878 7127
rect 41930 7115 41936 7167
rect 42256 7164 42262 7167
rect 42243 7158 42262 7164
rect 42243 7124 42255 7158
rect 42243 7118 42262 7124
rect 42256 7115 42262 7118
rect 42314 7115 42320 7167
rect 43504 7155 43510 7167
rect 42850 7127 43510 7155
rect 38419 7084 38477 7090
rect 38419 7050 38431 7084
rect 38465 7050 38477 7084
rect 39955 7084 40013 7090
rect 38419 7044 38477 7050
rect 38914 7053 39902 7081
rect 33235 7010 33293 7016
rect 33235 7007 33247 7010
rect 29314 6979 33247 7007
rect 28723 6970 28781 6976
rect 33235 6976 33247 6979
rect 33281 6976 33293 7010
rect 33235 6970 33293 6976
rect 37456 6967 37462 7019
rect 37514 7007 37520 7019
rect 38914 7007 38942 7053
rect 37514 6979 38942 7007
rect 37514 6967 37520 6979
rect 38992 6967 38998 7019
rect 39050 7007 39056 7019
rect 39283 7010 39341 7016
rect 39283 7007 39295 7010
rect 39050 6979 39295 7007
rect 39050 6967 39056 6979
rect 39283 6976 39295 6979
rect 39329 6976 39341 7010
rect 39874 7007 39902 7053
rect 39955 7050 39967 7084
rect 40001 7050 40013 7084
rect 39955 7044 40013 7050
rect 41491 7084 41549 7090
rect 41491 7050 41503 7084
rect 41537 7081 41549 7084
rect 42850 7081 42878 7127
rect 43504 7115 43510 7127
rect 43562 7115 43568 7167
rect 44944 7155 44950 7167
rect 44905 7127 44950 7155
rect 44944 7115 44950 7127
rect 45002 7155 45008 7167
rect 52240 7155 52246 7167
rect 45002 7127 45278 7155
rect 45002 7115 45008 7127
rect 43024 7081 43030 7093
rect 41537 7053 42878 7081
rect 42985 7053 43030 7081
rect 41537 7050 41549 7053
rect 41491 7044 41549 7050
rect 43024 7041 43030 7053
rect 43082 7041 43088 7093
rect 43408 7041 43414 7093
rect 43466 7081 43472 7093
rect 43699 7084 43757 7090
rect 43699 7081 43711 7084
rect 43466 7053 43711 7081
rect 43466 7041 43472 7053
rect 43699 7050 43711 7053
rect 43745 7050 43757 7084
rect 43699 7044 43757 7050
rect 43792 7041 43798 7093
rect 43850 7081 43856 7093
rect 45250 7090 45278 7127
rect 46786 7127 52246 7155
rect 46786 7090 46814 7127
rect 52240 7115 52246 7127
rect 52298 7115 52304 7167
rect 44179 7084 44237 7090
rect 44179 7081 44191 7084
rect 43850 7053 44191 7081
rect 43850 7041 43856 7053
rect 44179 7050 44191 7053
rect 44225 7081 44237 7084
rect 44467 7084 44525 7090
rect 44467 7081 44479 7084
rect 44225 7053 44479 7081
rect 44225 7050 44237 7053
rect 44179 7044 44237 7050
rect 44467 7050 44479 7053
rect 44513 7050 44525 7084
rect 44467 7044 44525 7050
rect 45235 7084 45293 7090
rect 45235 7050 45247 7084
rect 45281 7050 45293 7084
rect 45235 7044 45293 7050
rect 46771 7084 46829 7090
rect 46771 7050 46783 7084
rect 46817 7050 46829 7084
rect 48304 7081 48310 7093
rect 48265 7053 48310 7081
rect 46771 7044 46829 7050
rect 48304 7041 48310 7053
rect 48362 7041 48368 7093
rect 49072 7081 49078 7093
rect 49033 7053 49078 7081
rect 49072 7041 49078 7053
rect 49130 7041 49136 7093
rect 50128 7041 50134 7093
rect 50186 7081 50192 7093
rect 50323 7084 50381 7090
rect 50323 7081 50335 7084
rect 50186 7053 50335 7081
rect 50186 7041 50192 7053
rect 50323 7050 50335 7053
rect 50369 7050 50381 7084
rect 50323 7044 50381 7050
rect 52051 7084 52109 7090
rect 52051 7050 52063 7084
rect 52097 7081 52109 7084
rect 52144 7081 52150 7093
rect 52097 7053 52150 7081
rect 52097 7050 52109 7053
rect 52051 7044 52109 7050
rect 52144 7041 52150 7053
rect 52202 7041 52208 7093
rect 52816 7081 52822 7093
rect 52777 7053 52822 7081
rect 52816 7041 52822 7053
rect 52874 7041 52880 7093
rect 42163 7010 42221 7016
rect 42163 7007 42175 7010
rect 39874 6979 41822 7007
rect 39283 6970 39341 6976
rect 10978 6905 12974 6933
rect 10483 6896 10541 6902
rect 13456 6893 13462 6945
rect 13514 6933 13520 6945
rect 13555 6936 13613 6942
rect 13555 6933 13567 6936
rect 13514 6905 13567 6933
rect 13514 6893 13520 6905
rect 13555 6902 13567 6905
rect 13601 6902 13613 6936
rect 13555 6896 13613 6902
rect 14608 6893 14614 6945
rect 14666 6933 14672 6945
rect 15091 6936 15149 6942
rect 15091 6933 15103 6936
rect 14666 6905 15103 6933
rect 14666 6893 14672 6905
rect 15091 6902 15103 6905
rect 15137 6902 15149 6936
rect 15091 6896 15149 6902
rect 15376 6893 15382 6945
rect 15434 6933 15440 6945
rect 15763 6936 15821 6942
rect 15763 6933 15775 6936
rect 15434 6905 15775 6933
rect 15434 6893 15440 6905
rect 15763 6902 15775 6905
rect 15809 6902 15821 6936
rect 15763 6896 15821 6902
rect 17104 6893 17110 6945
rect 17162 6933 17168 6945
rect 17203 6936 17261 6942
rect 17203 6933 17215 6936
rect 17162 6905 17215 6933
rect 17162 6893 17168 6905
rect 17203 6902 17215 6905
rect 17249 6902 17261 6936
rect 17203 6896 17261 6902
rect 17872 6893 17878 6945
rect 17930 6933 17936 6945
rect 17971 6936 18029 6942
rect 17971 6933 17983 6936
rect 17930 6905 17983 6933
rect 17930 6893 17936 6905
rect 17971 6902 17983 6905
rect 18017 6902 18029 6936
rect 17971 6896 18029 6902
rect 18544 6893 18550 6945
rect 18602 6933 18608 6945
rect 18739 6936 18797 6942
rect 18739 6933 18751 6936
rect 18602 6905 18751 6933
rect 18602 6893 18608 6905
rect 18739 6902 18751 6905
rect 18785 6902 18797 6936
rect 20368 6933 20374 6945
rect 20329 6905 20374 6933
rect 18739 6896 18797 6902
rect 20368 6893 20374 6905
rect 20426 6893 20432 6945
rect 21043 6936 21101 6942
rect 21043 6902 21055 6936
rect 21089 6902 21101 6936
rect 21043 6896 21101 6902
rect 20656 6819 20662 6871
rect 20714 6859 20720 6871
rect 21058 6859 21086 6896
rect 21136 6893 21142 6945
rect 21194 6933 21200 6945
rect 21811 6936 21869 6942
rect 21811 6933 21823 6936
rect 21194 6905 21823 6933
rect 21194 6893 21200 6905
rect 21811 6902 21823 6905
rect 21857 6902 21869 6936
rect 21811 6896 21869 6902
rect 21904 6893 21910 6945
rect 21962 6933 21968 6945
rect 22579 6936 22637 6942
rect 22579 6933 22591 6936
rect 21962 6905 22591 6933
rect 21962 6893 21968 6905
rect 22579 6902 22591 6905
rect 22625 6902 22637 6936
rect 22579 6896 22637 6902
rect 23344 6893 23350 6945
rect 23402 6933 23408 6945
rect 23443 6936 23501 6942
rect 23443 6933 23455 6936
rect 23402 6905 23455 6933
rect 23402 6893 23408 6905
rect 23443 6902 23455 6905
rect 23489 6902 23501 6936
rect 24208 6933 24214 6945
rect 24169 6905 24214 6933
rect 23443 6896 23501 6902
rect 24208 6893 24214 6905
rect 24266 6893 24272 6945
rect 24496 6893 24502 6945
rect 24554 6933 24560 6945
rect 25555 6936 25613 6942
rect 25555 6933 25567 6936
rect 24554 6905 25567 6933
rect 24554 6893 24560 6905
rect 25555 6902 25567 6905
rect 25601 6902 25613 6936
rect 25555 6896 25613 6902
rect 26323 6936 26381 6942
rect 26323 6902 26335 6936
rect 26369 6902 26381 6936
rect 26323 6896 26381 6902
rect 20714 6831 21086 6859
rect 20714 6819 20720 6831
rect 25168 6819 25174 6871
rect 25226 6859 25232 6871
rect 26338 6859 26366 6896
rect 26896 6893 26902 6945
rect 26954 6933 26960 6945
rect 27187 6936 27245 6942
rect 27187 6933 27199 6936
rect 26954 6905 27199 6933
rect 26954 6893 26960 6905
rect 27187 6902 27199 6905
rect 27233 6902 27245 6936
rect 27859 6936 27917 6942
rect 27859 6933 27871 6936
rect 27187 6896 27245 6902
rect 27346 6905 27871 6933
rect 25226 6831 26366 6859
rect 25226 6819 25232 6831
rect 26992 6819 26998 6871
rect 27050 6859 27056 6871
rect 27346 6859 27374 6905
rect 27859 6902 27871 6905
rect 27905 6902 27917 6936
rect 27859 6896 27917 6902
rect 28627 6936 28685 6942
rect 28627 6902 28639 6936
rect 28673 6902 28685 6936
rect 29392 6933 29398 6945
rect 29353 6905 29398 6933
rect 28627 6896 28685 6902
rect 27050 6831 27374 6859
rect 27050 6819 27056 6831
rect 27760 6819 27766 6871
rect 27818 6859 27824 6871
rect 28642 6859 28670 6896
rect 29392 6893 29398 6905
rect 29450 6893 29456 6945
rect 29968 6893 29974 6945
rect 30026 6933 30032 6945
rect 30931 6936 30989 6942
rect 30931 6933 30943 6936
rect 30026 6905 30943 6933
rect 30026 6893 30032 6905
rect 30931 6902 30943 6905
rect 30977 6902 30989 6936
rect 30931 6896 30989 6902
rect 31699 6936 31757 6942
rect 31699 6902 31711 6936
rect 31745 6933 31757 6936
rect 31792 6933 31798 6945
rect 31745 6905 31798 6933
rect 31745 6902 31757 6905
rect 31699 6896 31757 6902
rect 31792 6893 31798 6905
rect 31850 6893 31856 6945
rect 32368 6933 32374 6945
rect 32329 6905 32374 6933
rect 32368 6893 32374 6905
rect 32426 6893 32432 6945
rect 33139 6936 33197 6942
rect 33139 6902 33151 6936
rect 33185 6902 33197 6936
rect 33139 6896 33197 6902
rect 33907 6936 33965 6942
rect 33907 6902 33919 6936
rect 33953 6902 33965 6936
rect 33907 6896 33965 6902
rect 27818 6831 28670 6859
rect 27818 6819 27824 6831
rect 32176 6819 32182 6871
rect 32234 6859 32240 6871
rect 33154 6859 33182 6896
rect 32234 6831 33182 6859
rect 32234 6819 32240 6831
rect 8234 6757 9758 6785
rect 8234 6745 8240 6757
rect 32944 6745 32950 6797
rect 33002 6785 33008 6797
rect 33922 6785 33950 6896
rect 34576 6893 34582 6945
rect 34634 6933 34640 6945
rect 34675 6936 34733 6942
rect 34675 6933 34687 6936
rect 34634 6905 34687 6933
rect 34634 6893 34640 6905
rect 34675 6902 34687 6905
rect 34721 6902 34733 6936
rect 34675 6896 34733 6902
rect 34771 6936 34829 6942
rect 34771 6902 34783 6936
rect 34817 6933 34829 6936
rect 35728 6933 35734 6945
rect 34817 6905 35734 6933
rect 34817 6902 34829 6905
rect 34771 6896 34829 6902
rect 35728 6893 35734 6905
rect 35786 6893 35792 6945
rect 35920 6893 35926 6945
rect 35978 6933 35984 6945
rect 36115 6936 36173 6942
rect 36115 6933 36127 6936
rect 35978 6905 36127 6933
rect 35978 6893 35984 6905
rect 36115 6902 36127 6905
rect 36161 6902 36173 6936
rect 36115 6896 36173 6902
rect 36400 6893 36406 6945
rect 36458 6933 36464 6945
rect 36883 6936 36941 6942
rect 36883 6933 36895 6936
rect 36458 6905 36895 6933
rect 36458 6893 36464 6905
rect 36883 6902 36895 6905
rect 36929 6902 36941 6936
rect 36883 6896 36941 6902
rect 36976 6893 36982 6945
rect 37034 6933 37040 6945
rect 37651 6936 37709 6942
rect 37651 6933 37663 6936
rect 37034 6905 37663 6933
rect 37034 6893 37040 6905
rect 37651 6902 37663 6905
rect 37697 6902 37709 6936
rect 38512 6933 38518 6945
rect 38473 6905 38518 6933
rect 37651 6896 37709 6902
rect 38512 6893 38518 6905
rect 38570 6893 38576 6945
rect 39187 6936 39245 6942
rect 39187 6902 39199 6936
rect 39233 6902 39245 6936
rect 39187 6896 39245 6902
rect 39475 6936 39533 6942
rect 39475 6902 39487 6936
rect 39521 6933 39533 6936
rect 40051 6936 40109 6942
rect 40051 6933 40063 6936
rect 39521 6905 40063 6933
rect 39521 6902 39533 6905
rect 39475 6896 39533 6902
rect 40051 6902 40063 6905
rect 40097 6902 40109 6936
rect 40051 6896 40109 6902
rect 41395 6936 41453 6942
rect 41395 6902 41407 6936
rect 41441 6902 41453 6936
rect 41395 6896 41453 6902
rect 33002 6757 33950 6785
rect 33002 6745 33008 6757
rect 37648 6745 37654 6797
rect 37706 6785 37712 6797
rect 39202 6785 39230 6896
rect 39856 6819 39862 6871
rect 39914 6859 39920 6871
rect 41410 6859 41438 6896
rect 39914 6831 41438 6859
rect 41794 6859 41822 6979
rect 42082 6979 42175 7007
rect 41872 6893 41878 6945
rect 41930 6933 41936 6945
rect 42082 6933 42110 6979
rect 42163 6976 42175 6979
rect 42209 6976 42221 7010
rect 47539 7010 47597 7016
rect 47539 7007 47551 7010
rect 42163 6970 42221 6976
rect 42370 6979 47551 7007
rect 42370 6933 42398 6979
rect 47539 6976 47551 6979
rect 47585 6976 47597 7010
rect 47539 6970 47597 6976
rect 54067 7010 54125 7016
rect 54067 6976 54079 7010
rect 54113 6976 54125 7010
rect 54736 7007 54742 7019
rect 54697 6979 54742 7007
rect 54067 6970 54125 6976
rect 42931 6936 42989 6942
rect 42931 6933 42943 6936
rect 41930 6905 42110 6933
rect 42274 6905 42398 6933
rect 42466 6905 42943 6933
rect 41930 6893 41936 6905
rect 42274 6859 42302 6905
rect 41794 6831 42302 6859
rect 39914 6819 39920 6831
rect 37706 6757 39230 6785
rect 37706 6745 37712 6757
rect 41104 6745 41110 6797
rect 41162 6785 41168 6797
rect 42466 6785 42494 6905
rect 42931 6902 42943 6905
rect 42977 6902 42989 6936
rect 43792 6933 43798 6945
rect 43753 6905 43798 6933
rect 42931 6896 42989 6902
rect 43792 6893 43798 6905
rect 43850 6893 43856 6945
rect 44563 6936 44621 6942
rect 44563 6902 44575 6936
rect 44609 6902 44621 6936
rect 44563 6896 44621 6902
rect 45331 6936 45389 6942
rect 45331 6902 45343 6936
rect 45377 6902 45389 6936
rect 45331 6896 45389 6902
rect 43600 6819 43606 6871
rect 43658 6859 43664 6871
rect 44578 6859 44606 6896
rect 43658 6831 44606 6859
rect 43658 6819 43664 6831
rect 43408 6785 43414 6797
rect 41162 6757 42494 6785
rect 43369 6757 43414 6785
rect 41162 6745 41168 6757
rect 43408 6745 43414 6757
rect 43466 6745 43472 6797
rect 44272 6745 44278 6797
rect 44330 6785 44336 6797
rect 45346 6785 45374 6896
rect 45424 6893 45430 6945
rect 45482 6933 45488 6945
rect 46675 6936 46733 6942
rect 46675 6933 46687 6936
rect 45482 6905 46687 6933
rect 45482 6893 45488 6905
rect 46675 6902 46687 6905
rect 46721 6902 46733 6936
rect 46675 6896 46733 6902
rect 46768 6893 46774 6945
rect 46826 6933 46832 6945
rect 47443 6936 47501 6942
rect 47443 6933 47455 6936
rect 46826 6905 47455 6933
rect 46826 6893 46832 6905
rect 47443 6902 47455 6905
rect 47489 6902 47501 6936
rect 47443 6896 47501 6902
rect 48211 6936 48269 6942
rect 48211 6902 48223 6936
rect 48257 6902 48269 6936
rect 48211 6896 48269 6902
rect 46864 6819 46870 6871
rect 46922 6859 46928 6871
rect 48226 6859 48254 6896
rect 48304 6893 48310 6945
rect 48362 6933 48368 6945
rect 48979 6936 49037 6942
rect 48979 6933 48991 6936
rect 48362 6905 48991 6933
rect 48362 6893 48368 6905
rect 48979 6902 48991 6905
rect 49025 6902 49037 6936
rect 48979 6896 49037 6902
rect 50128 6893 50134 6945
rect 50186 6933 50192 6945
rect 50227 6936 50285 6942
rect 50227 6933 50239 6936
rect 50186 6905 50239 6933
rect 50186 6893 50192 6905
rect 50227 6902 50239 6905
rect 50273 6902 50285 6936
rect 50227 6896 50285 6902
rect 51376 6893 51382 6945
rect 51434 6933 51440 6945
rect 51955 6936 52013 6942
rect 51955 6933 51967 6936
rect 51434 6905 51967 6933
rect 51434 6893 51440 6905
rect 51955 6902 51967 6905
rect 52001 6902 52013 6936
rect 51955 6896 52013 6902
rect 52432 6893 52438 6945
rect 52490 6933 52496 6945
rect 52723 6936 52781 6942
rect 52723 6933 52735 6936
rect 52490 6905 52735 6933
rect 52490 6893 52496 6905
rect 52723 6902 52735 6905
rect 52769 6902 52781 6936
rect 54082 6933 54110 6970
rect 54736 6967 54742 6979
rect 54794 6967 54800 7019
rect 55408 6967 55414 7019
rect 55466 7007 55472 7019
rect 55507 7010 55565 7016
rect 55507 7007 55519 7010
rect 55466 6979 55519 7007
rect 55466 6967 55472 6979
rect 55507 6976 55519 6979
rect 55553 6976 55565 7010
rect 55507 6970 55565 6976
rect 57811 7010 57869 7016
rect 57811 6976 57823 7010
rect 57857 7007 57869 7010
rect 58480 7007 58486 7019
rect 57857 6979 58486 7007
rect 57857 6976 57869 6979
rect 57811 6970 57869 6976
rect 58480 6967 58486 6979
rect 58538 6967 58544 7019
rect 56368 6933 56374 6945
rect 54082 6905 56374 6933
rect 52723 6896 52781 6902
rect 56368 6893 56374 6905
rect 56426 6893 56432 6945
rect 46922 6831 48254 6859
rect 46922 6819 46928 6831
rect 44330 6757 45374 6785
rect 44330 6745 44336 6757
rect 1152 6686 58848 6708
rect 1152 6634 4294 6686
rect 4346 6634 4358 6686
rect 4410 6634 4422 6686
rect 4474 6634 4486 6686
rect 4538 6634 35014 6686
rect 35066 6634 35078 6686
rect 35130 6634 35142 6686
rect 35194 6634 35206 6686
rect 35258 6634 58848 6686
rect 1152 6612 58848 6634
rect 8467 6566 8525 6572
rect 8467 6532 8479 6566
rect 8513 6563 8525 6566
rect 15088 6563 15094 6575
rect 8513 6535 8654 6563
rect 15049 6535 15094 6563
rect 8513 6532 8525 6535
rect 8467 6526 8525 6532
rect 7603 6492 7661 6498
rect 7603 6458 7615 6492
rect 7649 6489 7661 6492
rect 7699 6492 7757 6498
rect 7699 6489 7711 6492
rect 7649 6461 7711 6489
rect 7649 6458 7661 6461
rect 7603 6452 7661 6458
rect 7699 6458 7711 6461
rect 7745 6458 7757 6492
rect 8626 6489 8654 6535
rect 15088 6523 15094 6535
rect 15146 6563 15152 6575
rect 15856 6563 15862 6575
rect 15146 6535 15518 6563
rect 15817 6535 15862 6563
rect 15146 6523 15152 6535
rect 8944 6489 8950 6501
rect 8626 6475 8950 6489
rect 8640 6461 8950 6475
rect 7699 6452 7757 6458
rect 8944 6449 8950 6461
rect 9002 6449 9008 6501
rect 5395 6418 5453 6424
rect 5395 6384 5407 6418
rect 5441 6415 5453 6418
rect 5680 6415 5686 6427
rect 5441 6387 5686 6415
rect 5441 6384 5453 6387
rect 5395 6378 5453 6384
rect 5680 6375 5686 6387
rect 5738 6375 5744 6427
rect 6835 6418 6893 6424
rect 6835 6384 6847 6418
rect 6881 6415 6893 6418
rect 7120 6415 7126 6427
rect 6881 6387 7126 6415
rect 6881 6384 6893 6387
rect 6835 6378 6893 6384
rect 7120 6375 7126 6387
rect 7178 6375 7184 6427
rect 13936 6415 13942 6427
rect 13897 6387 13942 6415
rect 13936 6375 13942 6387
rect 13994 6375 14000 6427
rect 14704 6415 14710 6427
rect 14665 6387 14710 6415
rect 14704 6375 14710 6387
rect 14762 6375 14768 6427
rect 15490 6424 15518 6535
rect 15856 6523 15862 6535
rect 15914 6563 15920 6575
rect 20467 6566 20525 6572
rect 15914 6535 16190 6563
rect 15914 6523 15920 6535
rect 16162 6424 16190 6535
rect 20467 6532 20479 6566
rect 20513 6563 20525 6566
rect 20560 6563 20566 6575
rect 20513 6535 20566 6563
rect 20513 6532 20525 6535
rect 20467 6526 20525 6532
rect 20560 6523 20566 6535
rect 20618 6563 20624 6575
rect 24112 6563 24118 6575
rect 20618 6535 20798 6563
rect 24073 6535 24118 6563
rect 20618 6523 20624 6535
rect 15475 6418 15533 6424
rect 15475 6384 15487 6418
rect 15521 6384 15533 6418
rect 15475 6378 15533 6384
rect 16147 6418 16205 6424
rect 16147 6384 16159 6418
rect 16193 6384 16205 6418
rect 16147 6378 16205 6384
rect 16243 6418 16301 6424
rect 16243 6384 16255 6418
rect 16289 6384 16301 6418
rect 16243 6378 16301 6384
rect 17395 6418 17453 6424
rect 17395 6384 17407 6418
rect 17441 6415 17453 6418
rect 17680 6415 17686 6427
rect 17441 6387 17686 6415
rect 17441 6384 17453 6387
rect 17395 6378 17453 6384
rect 1552 6341 1558 6353
rect 1513 6313 1558 6341
rect 1552 6301 1558 6313
rect 1610 6301 1616 6353
rect 2032 6301 2038 6353
rect 2090 6341 2096 6353
rect 2323 6344 2381 6350
rect 2323 6341 2335 6344
rect 2090 6313 2335 6341
rect 2090 6301 2096 6313
rect 2323 6310 2335 6313
rect 2369 6310 2381 6344
rect 3184 6341 3190 6353
rect 3145 6313 3190 6341
rect 2323 6304 2381 6310
rect 3184 6301 3190 6313
rect 3242 6301 3248 6353
rect 3856 6301 3862 6353
rect 3914 6341 3920 6353
rect 3955 6344 4013 6350
rect 3955 6341 3967 6344
rect 3914 6313 3967 6341
rect 3914 6301 3920 6313
rect 3955 6310 3967 6313
rect 4001 6310 4013 6344
rect 3955 6304 4013 6310
rect 4624 6301 4630 6353
rect 4682 6341 4688 6353
rect 4723 6344 4781 6350
rect 4723 6341 4735 6344
rect 4682 6313 4735 6341
rect 4682 6301 4688 6313
rect 4723 6310 4735 6313
rect 4769 6310 4781 6344
rect 9424 6341 9430 6353
rect 9385 6313 9430 6341
rect 4723 6304 4781 6310
rect 9424 6301 9430 6313
rect 9482 6301 9488 6353
rect 10096 6301 10102 6353
rect 10154 6341 10160 6353
rect 10195 6344 10253 6350
rect 10195 6341 10207 6344
rect 10154 6313 10207 6341
rect 10154 6301 10160 6313
rect 10195 6310 10207 6313
rect 10241 6310 10253 6344
rect 10195 6304 10253 6310
rect 10864 6301 10870 6353
rect 10922 6341 10928 6353
rect 10963 6344 11021 6350
rect 10963 6341 10975 6344
rect 10922 6313 10975 6341
rect 10922 6301 10928 6313
rect 10963 6310 10975 6313
rect 11009 6310 11021 6344
rect 10963 6304 11021 6310
rect 11632 6301 11638 6353
rect 11690 6341 11696 6353
rect 12211 6344 12269 6350
rect 12211 6341 12223 6344
rect 11690 6313 12223 6341
rect 11690 6301 11696 6313
rect 12211 6310 12223 6313
rect 12257 6310 12269 6344
rect 12211 6304 12269 6310
rect 12304 6301 12310 6353
rect 12362 6341 12368 6353
rect 12979 6344 13037 6350
rect 12979 6341 12991 6344
rect 12362 6313 12991 6341
rect 12362 6301 12368 6313
rect 12979 6310 12991 6313
rect 13025 6310 13037 6344
rect 12979 6304 13037 6310
rect 14896 6301 14902 6353
rect 14954 6341 14960 6353
rect 16258 6341 16286 6378
rect 17680 6375 17686 6387
rect 17738 6375 17744 6427
rect 18163 6418 18221 6424
rect 18163 6384 18175 6418
rect 18209 6415 18221 6418
rect 18448 6415 18454 6427
rect 18209 6387 18454 6415
rect 18209 6384 18221 6387
rect 18163 6378 18221 6384
rect 18448 6375 18454 6387
rect 18506 6375 18512 6427
rect 18931 6418 18989 6424
rect 18931 6384 18943 6418
rect 18977 6415 18989 6418
rect 19216 6415 19222 6427
rect 18977 6387 19222 6415
rect 18977 6384 18989 6387
rect 18931 6378 18989 6384
rect 19216 6375 19222 6387
rect 19274 6375 19280 6427
rect 19987 6418 20045 6424
rect 19987 6384 19999 6418
rect 20033 6415 20045 6418
rect 20464 6415 20470 6427
rect 20033 6387 20470 6415
rect 20033 6384 20045 6387
rect 19987 6378 20045 6384
rect 20464 6375 20470 6387
rect 20522 6375 20528 6427
rect 20770 6424 20798 6535
rect 24112 6523 24118 6535
rect 24170 6563 24176 6575
rect 27856 6563 27862 6575
rect 24170 6535 24446 6563
rect 27817 6535 27862 6563
rect 24170 6523 24176 6535
rect 20659 6418 20717 6424
rect 20659 6384 20671 6418
rect 20705 6384 20717 6418
rect 20659 6378 20717 6384
rect 20755 6418 20813 6424
rect 20755 6384 20767 6418
rect 20801 6384 20813 6418
rect 21520 6415 21526 6427
rect 21481 6387 21526 6415
rect 20755 6378 20813 6384
rect 14954 6313 16286 6341
rect 14954 6301 14960 6313
rect 19312 6301 19318 6353
rect 19370 6341 19376 6353
rect 20674 6341 20702 6378
rect 21520 6375 21526 6387
rect 21578 6375 21584 6427
rect 22960 6415 22966 6427
rect 22921 6387 22966 6415
rect 22960 6375 22966 6387
rect 23018 6375 23024 6427
rect 23443 6418 23501 6424
rect 23443 6384 23455 6418
rect 23489 6415 23501 6418
rect 23632 6415 23638 6427
rect 23489 6387 23638 6415
rect 23489 6384 23501 6387
rect 23443 6378 23501 6384
rect 23632 6375 23638 6387
rect 23690 6375 23696 6427
rect 24418 6424 24446 6535
rect 27856 6523 27862 6535
rect 27914 6563 27920 6575
rect 33136 6563 33142 6575
rect 27914 6535 28190 6563
rect 33097 6535 33142 6563
rect 27914 6523 27920 6535
rect 28162 6424 28190 6535
rect 33136 6523 33142 6535
rect 33194 6563 33200 6575
rect 34672 6563 34678 6575
rect 33194 6535 33470 6563
rect 34633 6535 34678 6563
rect 33194 6523 33200 6535
rect 24403 6418 24461 6424
rect 24403 6384 24415 6418
rect 24449 6384 24461 6418
rect 24403 6378 24461 6384
rect 28147 6418 28205 6424
rect 28147 6384 28159 6418
rect 28193 6384 28205 6418
rect 28147 6378 28205 6384
rect 28723 6418 28781 6424
rect 28723 6384 28735 6418
rect 28769 6415 28781 6418
rect 29008 6415 29014 6427
rect 28769 6387 29014 6415
rect 28769 6384 28781 6387
rect 28723 6378 28781 6384
rect 29008 6375 29014 6387
rect 29066 6375 29072 6427
rect 33442 6424 33470 6535
rect 34672 6523 34678 6535
rect 34730 6563 34736 6575
rect 34730 6535 35006 6563
rect 34730 6523 34736 6535
rect 33427 6418 33485 6424
rect 33427 6384 33439 6418
rect 33473 6384 33485 6418
rect 34288 6415 34294 6427
rect 34249 6387 34294 6415
rect 33427 6378 33485 6384
rect 34288 6375 34294 6387
rect 34346 6375 34352 6427
rect 34978 6424 35006 6535
rect 35728 6523 35734 6575
rect 35786 6563 35792 6575
rect 35827 6566 35885 6572
rect 35827 6563 35839 6566
rect 35786 6535 35839 6563
rect 35786 6523 35792 6535
rect 35827 6532 35839 6535
rect 35873 6532 35885 6566
rect 35827 6526 35885 6532
rect 41296 6523 41302 6575
rect 41354 6563 41360 6575
rect 42256 6563 42262 6575
rect 41354 6535 42262 6563
rect 41354 6523 41360 6535
rect 42256 6523 42262 6535
rect 42314 6523 42320 6575
rect 57040 6449 57046 6501
rect 57098 6449 57104 6501
rect 34963 6418 35021 6424
rect 34963 6384 34975 6418
rect 35009 6384 35021 6418
rect 34963 6378 35021 6384
rect 35059 6418 35117 6424
rect 35059 6384 35071 6418
rect 35105 6384 35117 6418
rect 35059 6378 35117 6384
rect 25648 6341 25654 6353
rect 19370 6313 20702 6341
rect 25609 6313 25654 6341
rect 19370 6301 19376 6313
rect 25648 6301 25654 6313
rect 25706 6301 25712 6353
rect 26800 6341 26806 6353
rect 26761 6313 26806 6341
rect 26800 6301 26806 6313
rect 26858 6301 26864 6353
rect 29680 6341 29686 6353
rect 29641 6313 29686 6341
rect 29680 6301 29686 6313
rect 29738 6301 29744 6353
rect 31216 6341 31222 6353
rect 31177 6313 31222 6341
rect 31216 6301 31222 6313
rect 31274 6301 31280 6353
rect 33808 6301 33814 6353
rect 33866 6341 33872 6353
rect 35074 6341 35102 6378
rect 35440 6375 35446 6427
rect 35498 6415 35504 6427
rect 37267 6418 37325 6424
rect 37267 6415 37279 6418
rect 35498 6387 37279 6415
rect 35498 6375 35504 6387
rect 37267 6384 37279 6387
rect 37313 6384 37325 6418
rect 37267 6378 37325 6384
rect 41011 6418 41069 6424
rect 41011 6384 41023 6418
rect 41057 6415 41069 6418
rect 41200 6415 41206 6427
rect 41057 6387 41206 6415
rect 41057 6384 41069 6387
rect 41011 6378 41069 6384
rect 41200 6375 41206 6387
rect 41258 6375 41264 6427
rect 42832 6415 42838 6427
rect 42793 6387 42838 6415
rect 42832 6375 42838 6387
rect 42890 6375 42896 6427
rect 44080 6415 44086 6427
rect 44041 6387 44086 6415
rect 44080 6375 44086 6387
rect 44138 6375 44144 6427
rect 44656 6375 44662 6427
rect 44714 6415 44720 6427
rect 44851 6418 44909 6424
rect 44851 6415 44863 6418
rect 44714 6387 44863 6415
rect 44714 6375 44720 6387
rect 44851 6384 44863 6387
rect 44897 6384 44909 6418
rect 44851 6378 44909 6384
rect 50611 6418 50669 6424
rect 50611 6384 50623 6418
rect 50657 6415 50669 6418
rect 50800 6415 50806 6427
rect 50657 6387 50806 6415
rect 50657 6384 50669 6387
rect 50611 6378 50669 6384
rect 50800 6375 50806 6387
rect 50858 6375 50864 6427
rect 51379 6418 51437 6424
rect 51379 6384 51391 6418
rect 51425 6415 51437 6418
rect 51568 6415 51574 6427
rect 51425 6387 51574 6415
rect 51425 6384 51437 6387
rect 51379 6378 51437 6384
rect 51568 6375 51574 6387
rect 51626 6375 51632 6427
rect 57058 6415 57086 6449
rect 53314 6387 57086 6415
rect 36304 6341 36310 6353
rect 33866 6313 35102 6341
rect 36265 6313 36310 6341
rect 33866 6301 33872 6313
rect 36304 6301 36310 6313
rect 36362 6301 36368 6353
rect 38896 6341 38902 6353
rect 38857 6313 38902 6341
rect 38896 6301 38902 6313
rect 38954 6301 38960 6353
rect 40336 6341 40342 6353
rect 40297 6313 40342 6341
rect 40336 6301 40342 6313
rect 40394 6301 40400 6353
rect 41872 6341 41878 6353
rect 41833 6313 41878 6341
rect 41872 6301 41878 6313
rect 41930 6301 41936 6353
rect 45520 6341 45526 6353
rect 45481 6313 45526 6341
rect 45520 6301 45526 6313
rect 45578 6301 45584 6353
rect 46960 6341 46966 6353
rect 46921 6313 46966 6341
rect 46960 6301 46966 6313
rect 47018 6301 47024 6353
rect 47728 6341 47734 6353
rect 47689 6313 47734 6341
rect 47728 6301 47734 6313
rect 47786 6301 47792 6353
rect 48784 6301 48790 6353
rect 48842 6341 48848 6353
rect 49171 6344 49229 6350
rect 49171 6341 49183 6344
rect 48842 6313 49183 6341
rect 48842 6301 48848 6313
rect 49171 6310 49183 6313
rect 49217 6310 49229 6344
rect 49171 6304 49229 6310
rect 49552 6301 49558 6353
rect 49610 6341 49616 6353
rect 53314 6350 53342 6387
rect 49939 6344 49997 6350
rect 49939 6341 49951 6344
rect 49610 6313 49951 6341
rect 49610 6301 49616 6313
rect 49939 6310 49951 6313
rect 49985 6310 49997 6344
rect 49939 6304 49997 6310
rect 53299 6344 53357 6350
rect 53299 6310 53311 6344
rect 53345 6310 53357 6344
rect 53299 6304 53357 6310
rect 53968 6301 53974 6353
rect 54026 6341 54032 6353
rect 54451 6344 54509 6350
rect 54451 6341 54463 6344
rect 54026 6313 54463 6341
rect 54026 6301 54032 6313
rect 54451 6310 54463 6313
rect 54497 6310 54509 6344
rect 55216 6341 55222 6353
rect 55177 6313 55222 6341
rect 54451 6304 54509 6310
rect 55216 6301 55222 6313
rect 55274 6301 55280 6353
rect 55987 6344 56045 6350
rect 55987 6310 55999 6344
rect 56033 6310 56045 6344
rect 55987 6304 56045 6310
rect 57043 6344 57101 6350
rect 57043 6310 57055 6344
rect 57089 6310 57101 6344
rect 57043 6304 57101 6310
rect 57811 6344 57869 6350
rect 57811 6310 57823 6344
rect 57857 6341 57869 6344
rect 58096 6341 58102 6353
rect 57857 6313 58102 6341
rect 57857 6310 57869 6313
rect 57811 6304 57869 6310
rect 30640 6267 30646 6279
rect 30601 6239 30646 6267
rect 30640 6227 30646 6239
rect 30698 6227 30704 6279
rect 32179 6270 32237 6276
rect 32179 6236 32191 6270
rect 32225 6236 32237 6270
rect 32179 6230 32237 6236
rect 8080 6193 8086 6205
rect 7968 6165 8086 6193
rect 8080 6153 8086 6165
rect 8138 6153 8144 6205
rect 8368 6193 8374 6205
rect 8256 6165 8374 6193
rect 8368 6153 8374 6165
rect 8426 6153 8432 6205
rect 14128 6153 14134 6205
rect 14186 6193 14192 6205
rect 14186 6165 15422 6193
rect 14186 6153 14192 6165
rect 5488 6079 5494 6131
rect 5546 6119 5552 6131
rect 5587 6122 5645 6128
rect 5587 6119 5599 6122
rect 5546 6091 5599 6119
rect 5546 6079 5552 6091
rect 5587 6088 5599 6091
rect 5633 6088 5645 6122
rect 5587 6082 5645 6088
rect 6256 6079 6262 6131
rect 6314 6119 6320 6131
rect 7027 6122 7085 6128
rect 7027 6119 7039 6122
rect 6314 6091 7039 6119
rect 6314 6079 6320 6091
rect 7027 6088 7039 6091
rect 7073 6088 7085 6122
rect 7027 6082 7085 6088
rect 13072 6079 13078 6131
rect 13130 6119 13136 6131
rect 13843 6122 13901 6128
rect 13843 6119 13855 6122
rect 13130 6091 13855 6119
rect 13130 6079 13136 6091
rect 13843 6088 13855 6091
rect 13889 6088 13901 6122
rect 13843 6082 13901 6088
rect 13936 6079 13942 6131
rect 13994 6119 14000 6131
rect 15394 6128 15422 6165
rect 16816 6153 16822 6205
rect 16874 6193 16880 6205
rect 16874 6165 17630 6193
rect 16874 6153 16880 6165
rect 17602 6128 17630 6165
rect 18256 6153 18262 6205
rect 18314 6193 18320 6205
rect 18314 6165 18494 6193
rect 18314 6153 18320 6165
rect 14611 6122 14669 6128
rect 14611 6119 14623 6122
rect 13994 6091 14623 6119
rect 13994 6079 14000 6091
rect 14611 6088 14623 6091
rect 14657 6088 14669 6122
rect 14611 6082 14669 6088
rect 15379 6122 15437 6128
rect 15379 6088 15391 6122
rect 15425 6088 15437 6122
rect 15379 6082 15437 6088
rect 17587 6122 17645 6128
rect 17587 6088 17599 6122
rect 17633 6088 17645 6122
rect 18352 6119 18358 6131
rect 18313 6091 18358 6119
rect 17587 6082 17645 6088
rect 18352 6079 18358 6091
rect 18410 6079 18416 6131
rect 18466 6119 18494 6165
rect 18928 6153 18934 6205
rect 18986 6193 18992 6205
rect 32194 6193 32222 6230
rect 36880 6227 36886 6279
rect 36938 6267 36944 6279
rect 37171 6270 37229 6276
rect 37171 6267 37183 6270
rect 36938 6239 37183 6267
rect 36938 6227 36944 6239
rect 37171 6236 37183 6239
rect 37217 6236 37229 6270
rect 37171 6230 37229 6236
rect 40624 6227 40630 6279
rect 40682 6267 40688 6279
rect 52435 6270 52493 6276
rect 40682 6239 41438 6267
rect 40682 6227 40688 6239
rect 40816 6193 40822 6205
rect 18986 6165 19934 6193
rect 18986 6153 18992 6165
rect 19906 6128 19934 6165
rect 27346 6165 28286 6193
rect 32194 6165 40822 6193
rect 19123 6122 19181 6128
rect 19123 6119 19135 6122
rect 18466 6091 19135 6119
rect 19123 6088 19135 6091
rect 19169 6088 19181 6122
rect 19123 6082 19181 6088
rect 19891 6122 19949 6128
rect 19891 6088 19903 6122
rect 19937 6088 19949 6122
rect 21424 6119 21430 6131
rect 21385 6091 21430 6119
rect 19891 6082 19949 6088
rect 21424 6079 21430 6091
rect 21482 6079 21488 6131
rect 21520 6079 21526 6131
rect 21578 6119 21584 6131
rect 22867 6122 22925 6128
rect 22867 6119 22879 6122
rect 21578 6091 22879 6119
rect 21578 6079 21584 6091
rect 22867 6088 22879 6091
rect 22913 6088 22925 6122
rect 22867 6082 22925 6088
rect 23632 6079 23638 6131
rect 23690 6119 23696 6131
rect 23731 6122 23789 6128
rect 23731 6119 23743 6122
rect 23690 6091 23743 6119
rect 23690 6079 23696 6091
rect 23731 6088 23743 6091
rect 23777 6088 23789 6122
rect 23731 6082 23789 6088
rect 23920 6079 23926 6131
rect 23978 6119 23984 6131
rect 24499 6122 24557 6128
rect 24499 6119 24511 6122
rect 23978 6091 24511 6119
rect 23978 6079 23984 6091
rect 24499 6088 24511 6091
rect 24545 6088 24557 6122
rect 24499 6082 24557 6088
rect 26320 6079 26326 6131
rect 26378 6119 26384 6131
rect 27346 6119 27374 6165
rect 28258 6128 28286 6165
rect 40816 6153 40822 6165
rect 40874 6153 40880 6205
rect 26378 6091 27374 6119
rect 28243 6122 28301 6128
rect 26378 6079 26384 6091
rect 28243 6088 28255 6122
rect 28289 6088 28301 6122
rect 28243 6082 28301 6088
rect 28432 6079 28438 6131
rect 28490 6119 28496 6131
rect 28915 6122 28973 6128
rect 28915 6119 28927 6122
rect 28490 6091 28927 6119
rect 28490 6079 28496 6091
rect 28915 6088 28927 6091
rect 28961 6088 28973 6122
rect 28915 6082 28973 6088
rect 29776 6079 29782 6131
rect 29834 6119 29840 6131
rect 30547 6122 30605 6128
rect 30547 6119 30559 6122
rect 29834 6091 30559 6119
rect 29834 6079 29840 6091
rect 30547 6088 30559 6091
rect 30593 6088 30605 6122
rect 30547 6082 30605 6088
rect 30736 6079 30742 6131
rect 30794 6119 30800 6131
rect 32083 6122 32141 6128
rect 32083 6119 32095 6122
rect 30794 6091 32095 6119
rect 30794 6079 30800 6091
rect 32083 6088 32095 6091
rect 32129 6088 32141 6122
rect 33520 6119 33526 6131
rect 33481 6091 33526 6119
rect 32083 6082 32141 6088
rect 33520 6079 33526 6091
rect 33578 6079 33584 6131
rect 33712 6079 33718 6131
rect 33770 6119 33776 6131
rect 34195 6122 34253 6128
rect 34195 6119 34207 6122
rect 33770 6091 34207 6119
rect 33770 6079 33776 6091
rect 34195 6088 34207 6091
rect 34241 6088 34253 6122
rect 36880 6119 36886 6131
rect 36841 6091 36886 6119
rect 34195 6082 34253 6088
rect 36880 6079 36886 6091
rect 36938 6079 36944 6131
rect 39952 6079 39958 6131
rect 40010 6119 40016 6131
rect 41299 6122 41357 6128
rect 41299 6119 41311 6122
rect 40010 6091 41311 6119
rect 40010 6079 40016 6091
rect 41299 6088 41311 6091
rect 41345 6088 41357 6122
rect 41410 6119 41438 6239
rect 52435 6236 52447 6270
rect 52481 6267 52493 6270
rect 55120 6267 55126 6279
rect 52481 6239 55126 6267
rect 52481 6236 52493 6239
rect 52435 6230 52493 6236
rect 55120 6227 55126 6239
rect 55178 6227 55184 6279
rect 42640 6153 42646 6205
rect 42698 6193 42704 6205
rect 42698 6165 44030 6193
rect 42698 6153 42704 6165
rect 44002 6128 44030 6165
rect 51568 6153 51574 6205
rect 51626 6193 51632 6205
rect 51626 6165 52382 6193
rect 51626 6153 51632 6165
rect 42739 6122 42797 6128
rect 42739 6119 42751 6122
rect 41410 6091 42751 6119
rect 41299 6082 41357 6088
rect 42739 6088 42751 6091
rect 42785 6088 42797 6122
rect 42739 6082 42797 6088
rect 43987 6122 44045 6128
rect 43987 6088 43999 6122
rect 44033 6088 44045 6122
rect 43987 6082 44045 6088
rect 44080 6079 44086 6131
rect 44138 6119 44144 6131
rect 44755 6122 44813 6128
rect 44755 6119 44767 6122
rect 44138 6091 44767 6119
rect 44138 6079 44144 6091
rect 44755 6088 44767 6091
rect 44801 6088 44813 6122
rect 44755 6082 44813 6088
rect 49744 6079 49750 6131
rect 49802 6119 49808 6131
rect 50899 6122 50957 6128
rect 50899 6119 50911 6122
rect 49802 6091 50911 6119
rect 49802 6079 49808 6091
rect 50899 6088 50911 6091
rect 50945 6088 50957 6122
rect 50899 6082 50957 6088
rect 51088 6079 51094 6131
rect 51146 6119 51152 6131
rect 52354 6128 52382 6165
rect 55024 6153 55030 6205
rect 55082 6193 55088 6205
rect 56002 6193 56030 6304
rect 57058 6267 57086 6304
rect 58096 6301 58102 6313
rect 58154 6301 58160 6353
rect 58864 6267 58870 6279
rect 57058 6239 58870 6267
rect 58864 6227 58870 6239
rect 58922 6227 58928 6279
rect 55082 6165 56030 6193
rect 55082 6153 55088 6165
rect 51667 6122 51725 6128
rect 51667 6119 51679 6122
rect 51146 6091 51679 6119
rect 51146 6079 51152 6091
rect 51667 6088 51679 6091
rect 51713 6088 51725 6122
rect 51667 6082 51725 6088
rect 52339 6122 52397 6128
rect 52339 6088 52351 6122
rect 52385 6088 52397 6122
rect 52339 6082 52397 6088
rect 1152 6020 58848 6042
rect 1152 5968 19654 6020
rect 19706 5968 19718 6020
rect 19770 5968 19782 6020
rect 19834 5968 19846 6020
rect 19898 5968 50374 6020
rect 50426 5968 50438 6020
rect 50490 5968 50502 6020
rect 50554 5968 50566 6020
rect 50618 5968 58848 6020
rect 1152 5946 58848 5968
rect 5776 5857 5782 5909
rect 5834 5897 5840 5909
rect 17584 5897 17590 5909
rect 5834 5869 17590 5897
rect 5834 5857 5840 5869
rect 17584 5857 17590 5869
rect 17642 5857 17648 5909
rect 2608 5783 2614 5835
rect 2666 5823 2672 5835
rect 8368 5823 8374 5835
rect 2666 5795 8374 5823
rect 2666 5783 2672 5795
rect 8368 5783 8374 5795
rect 8426 5783 8432 5835
rect 8848 5783 8854 5835
rect 8906 5823 8912 5835
rect 9808 5823 9814 5835
rect 8906 5795 9814 5823
rect 8906 5783 8912 5795
rect 9808 5783 9814 5795
rect 9866 5783 9872 5835
rect 5008 5709 5014 5761
rect 5066 5749 5072 5761
rect 5779 5752 5837 5758
rect 5779 5749 5791 5752
rect 5066 5721 5791 5749
rect 5066 5709 5072 5721
rect 5779 5718 5791 5721
rect 5825 5749 5837 5752
rect 5971 5752 6029 5758
rect 5971 5749 5983 5752
rect 5825 5721 5983 5749
rect 5825 5718 5837 5721
rect 5779 5712 5837 5718
rect 5971 5718 5983 5721
rect 6017 5718 6029 5752
rect 5971 5712 6029 5718
rect 7024 5709 7030 5761
rect 7082 5749 7088 5761
rect 11539 5752 11597 5758
rect 7082 5721 9950 5749
rect 7082 5709 7088 5721
rect 1072 5635 1078 5687
rect 1130 5675 1136 5687
rect 1555 5678 1613 5684
rect 1555 5675 1567 5678
rect 1130 5647 1567 5675
rect 1130 5635 1136 5647
rect 1555 5644 1567 5647
rect 1601 5644 1613 5678
rect 1555 5638 1613 5644
rect 2896 5635 2902 5687
rect 2954 5675 2960 5687
rect 4435 5678 4493 5684
rect 2954 5647 2999 5675
rect 2954 5635 2960 5647
rect 4435 5644 4447 5678
rect 4481 5675 4493 5678
rect 4912 5675 4918 5687
rect 4481 5647 4918 5675
rect 4481 5644 4493 5647
rect 4435 5638 4493 5644
rect 4912 5635 4918 5647
rect 4970 5635 4976 5687
rect 5104 5675 5110 5687
rect 5065 5647 5110 5675
rect 5104 5635 5110 5647
rect 5162 5635 5168 5687
rect 6832 5675 6838 5687
rect 6793 5647 6838 5675
rect 6832 5635 6838 5647
rect 6890 5635 6896 5687
rect 7216 5635 7222 5687
rect 7274 5675 7280 5687
rect 7603 5678 7661 5684
rect 7603 5675 7615 5678
rect 7274 5647 7615 5675
rect 7274 5635 7280 5647
rect 7603 5644 7615 5647
rect 7649 5644 7661 5678
rect 7603 5638 7661 5644
rect 8371 5678 8429 5684
rect 8371 5644 8383 5678
rect 8417 5644 8429 5678
rect 8371 5638 8429 5644
rect 6067 5604 6125 5610
rect 6067 5570 6079 5604
rect 6113 5570 6125 5604
rect 6067 5564 6125 5570
rect 5776 5487 5782 5539
rect 5834 5527 5840 5539
rect 6082 5527 6110 5564
rect 5834 5499 6110 5527
rect 5834 5487 5840 5499
rect 7600 5487 7606 5539
rect 7658 5527 7664 5539
rect 8386 5527 8414 5638
rect 8752 5635 8758 5687
rect 8810 5675 8816 5687
rect 9619 5678 9677 5684
rect 9619 5675 9631 5678
rect 8810 5647 9631 5675
rect 8810 5635 8816 5647
rect 9619 5644 9631 5647
rect 9665 5644 9677 5678
rect 9619 5638 9677 5644
rect 7658 5499 8414 5527
rect 9922 5527 9950 5721
rect 11539 5718 11551 5752
rect 11585 5749 11597 5752
rect 43408 5749 43414 5761
rect 11585 5721 43414 5749
rect 11585 5718 11597 5721
rect 11539 5712 11597 5718
rect 43408 5709 43414 5721
rect 43466 5709 43472 5761
rect 10192 5635 10198 5687
rect 10250 5675 10256 5687
rect 10387 5678 10445 5684
rect 10387 5675 10399 5678
rect 10250 5647 10399 5675
rect 10250 5635 10256 5647
rect 10387 5644 10399 5647
rect 10433 5644 10445 5678
rect 10387 5638 10445 5644
rect 10480 5635 10486 5687
rect 10538 5675 10544 5687
rect 11155 5678 11213 5684
rect 11155 5675 11167 5678
rect 10538 5647 11167 5675
rect 10538 5635 10544 5647
rect 11155 5644 11167 5647
rect 11201 5644 11213 5678
rect 12592 5675 12598 5687
rect 12553 5647 12598 5675
rect 11155 5638 11213 5644
rect 12592 5635 12598 5647
rect 12650 5635 12656 5687
rect 13360 5675 13366 5687
rect 13321 5647 13366 5675
rect 13360 5635 13366 5647
rect 13418 5635 13424 5687
rect 14992 5675 14998 5687
rect 14953 5647 14998 5675
rect 14992 5635 14998 5647
rect 15050 5635 15056 5687
rect 15856 5675 15862 5687
rect 15817 5647 15862 5675
rect 15856 5635 15862 5647
rect 15914 5635 15920 5687
rect 16240 5635 16246 5687
rect 16298 5675 16304 5687
rect 16531 5678 16589 5684
rect 16531 5675 16543 5678
rect 16298 5647 16543 5675
rect 16298 5635 16304 5647
rect 16531 5644 16543 5647
rect 16577 5644 16589 5678
rect 16531 5638 16589 5644
rect 17296 5635 17302 5687
rect 17354 5675 17360 5687
rect 18736 5675 18742 5687
rect 17354 5647 17399 5675
rect 18697 5647 18742 5675
rect 17354 5635 17360 5647
rect 18736 5635 18742 5647
rect 18794 5635 18800 5687
rect 20176 5675 20182 5687
rect 20137 5647 20182 5675
rect 20176 5635 20182 5647
rect 20234 5635 20240 5687
rect 20560 5635 20566 5687
rect 20618 5675 20624 5687
rect 20947 5678 21005 5684
rect 20947 5675 20959 5678
rect 20618 5647 20959 5675
rect 20618 5635 20624 5647
rect 20947 5644 20959 5647
rect 20993 5644 21005 5678
rect 20947 5638 21005 5644
rect 21619 5678 21677 5684
rect 21619 5644 21631 5678
rect 21665 5675 21677 5678
rect 21715 5678 21773 5684
rect 21715 5675 21727 5678
rect 21665 5647 21727 5675
rect 21665 5644 21677 5647
rect 21619 5638 21677 5644
rect 21715 5644 21727 5647
rect 21761 5644 21773 5678
rect 21715 5638 21773 5644
rect 21808 5635 21814 5687
rect 21866 5675 21872 5687
rect 22483 5678 22541 5684
rect 22483 5675 22495 5678
rect 21866 5647 22495 5675
rect 21866 5635 21872 5647
rect 22483 5644 22495 5647
rect 22529 5644 22541 5678
rect 22483 5638 22541 5644
rect 23056 5635 23062 5687
rect 23114 5675 23120 5687
rect 23251 5678 23309 5684
rect 23251 5675 23263 5678
rect 23114 5647 23263 5675
rect 23114 5635 23120 5647
rect 23251 5644 23263 5647
rect 23297 5644 23309 5678
rect 23251 5638 23309 5644
rect 23440 5635 23446 5687
rect 23498 5675 23504 5687
rect 24019 5678 24077 5684
rect 24019 5675 24031 5678
rect 23498 5647 24031 5675
rect 23498 5635 23504 5647
rect 24019 5644 24031 5647
rect 24065 5644 24077 5678
rect 24019 5638 24077 5644
rect 24592 5635 24598 5687
rect 24650 5675 24656 5687
rect 25459 5678 25517 5684
rect 25459 5675 25471 5678
rect 24650 5647 25471 5675
rect 24650 5635 24656 5647
rect 25459 5644 25471 5647
rect 25505 5644 25517 5678
rect 26224 5675 26230 5687
rect 26185 5647 26230 5675
rect 25459 5638 25517 5644
rect 26224 5635 26230 5647
rect 26282 5635 26288 5687
rect 26611 5678 26669 5684
rect 26611 5644 26623 5678
rect 26657 5675 26669 5678
rect 26995 5678 27053 5684
rect 26995 5675 27007 5678
rect 26657 5647 27007 5675
rect 26657 5644 26669 5647
rect 26611 5638 26669 5644
rect 26995 5644 27007 5647
rect 27041 5644 27053 5678
rect 26995 5638 27053 5644
rect 27376 5635 27382 5687
rect 27434 5675 27440 5687
rect 27763 5678 27821 5684
rect 27763 5675 27775 5678
rect 27434 5647 27775 5675
rect 27434 5635 27440 5647
rect 27763 5644 27775 5647
rect 27809 5644 27821 5678
rect 27763 5638 27821 5644
rect 27856 5635 27862 5687
rect 27914 5675 27920 5687
rect 28531 5678 28589 5684
rect 28531 5675 28543 5678
rect 27914 5647 28543 5675
rect 27914 5635 27920 5647
rect 28531 5644 28543 5647
rect 28577 5644 28589 5678
rect 28531 5638 28589 5644
rect 28816 5635 28822 5687
rect 28874 5675 28880 5687
rect 29299 5678 29357 5684
rect 29299 5675 29311 5678
rect 28874 5647 29311 5675
rect 28874 5635 28880 5647
rect 29299 5644 29311 5647
rect 29345 5644 29357 5678
rect 29299 5638 29357 5644
rect 30256 5635 30262 5687
rect 30314 5675 30320 5687
rect 30739 5678 30797 5684
rect 30739 5675 30751 5678
rect 30314 5647 30751 5675
rect 30314 5635 30320 5647
rect 30739 5644 30751 5647
rect 30785 5644 30797 5678
rect 30739 5638 30797 5644
rect 30832 5635 30838 5687
rect 30890 5675 30896 5687
rect 31507 5678 31565 5684
rect 31507 5675 31519 5678
rect 30890 5647 31519 5675
rect 30890 5635 30896 5647
rect 31507 5644 31519 5647
rect 31553 5644 31565 5678
rect 31507 5638 31565 5644
rect 31696 5635 31702 5687
rect 31754 5675 31760 5687
rect 32275 5678 32333 5684
rect 32275 5675 32287 5678
rect 31754 5647 32287 5675
rect 31754 5635 31760 5647
rect 32275 5644 32287 5647
rect 32321 5644 32333 5678
rect 33136 5675 33142 5687
rect 33097 5647 33142 5675
rect 32275 5638 32333 5644
rect 33136 5635 33142 5647
rect 33194 5635 33200 5687
rect 33232 5635 33238 5687
rect 33290 5675 33296 5687
rect 33811 5678 33869 5684
rect 33811 5675 33823 5678
rect 33290 5647 33823 5675
rect 33290 5635 33296 5647
rect 33811 5644 33823 5647
rect 33857 5644 33869 5678
rect 34672 5675 34678 5687
rect 34633 5647 34678 5675
rect 33811 5638 33869 5644
rect 34672 5635 34678 5647
rect 34730 5635 34736 5687
rect 36016 5675 36022 5687
rect 35977 5647 36022 5675
rect 36016 5635 36022 5647
rect 36074 5635 36080 5687
rect 36208 5635 36214 5687
rect 36266 5675 36272 5687
rect 36787 5678 36845 5684
rect 36787 5675 36799 5678
rect 36266 5647 36799 5675
rect 36266 5635 36272 5647
rect 36787 5644 36799 5647
rect 36833 5644 36845 5678
rect 37552 5675 37558 5687
rect 37513 5647 37558 5675
rect 36787 5638 36845 5644
rect 37552 5635 37558 5647
rect 37610 5635 37616 5687
rect 38323 5678 38381 5684
rect 38323 5644 38335 5678
rect 38369 5644 38381 5678
rect 39088 5675 39094 5687
rect 39049 5647 39094 5675
rect 38323 5638 38381 5644
rect 36880 5601 36886 5613
rect 12946 5573 36886 5601
rect 12946 5527 12974 5573
rect 36880 5561 36886 5573
rect 36938 5561 36944 5613
rect 37456 5561 37462 5613
rect 37514 5601 37520 5613
rect 38338 5601 38366 5638
rect 39088 5635 39094 5647
rect 39146 5635 39152 5687
rect 39280 5635 39286 5687
rect 39338 5675 39344 5687
rect 39859 5678 39917 5684
rect 39859 5675 39871 5678
rect 39338 5647 39871 5675
rect 39338 5635 39344 5647
rect 39859 5644 39871 5647
rect 39905 5644 39917 5678
rect 39859 5638 39917 5644
rect 40720 5635 40726 5687
rect 40778 5675 40784 5687
rect 41299 5678 41357 5684
rect 41299 5675 41311 5678
rect 40778 5647 41311 5675
rect 40778 5635 40784 5647
rect 41299 5644 41311 5647
rect 41345 5644 41357 5678
rect 42064 5675 42070 5687
rect 42025 5647 42070 5675
rect 41299 5638 41357 5644
rect 42064 5635 42070 5647
rect 42122 5635 42128 5687
rect 42256 5635 42262 5687
rect 42314 5675 42320 5687
rect 42835 5678 42893 5684
rect 42835 5675 42847 5678
rect 42314 5647 42847 5675
rect 42314 5635 42320 5647
rect 42835 5644 42847 5647
rect 42881 5644 42893 5678
rect 42835 5638 42893 5644
rect 43216 5635 43222 5687
rect 43274 5675 43280 5687
rect 43603 5678 43661 5684
rect 43603 5675 43615 5678
rect 43274 5647 43615 5675
rect 43274 5635 43280 5647
rect 43603 5644 43615 5647
rect 43649 5644 43661 5678
rect 43603 5638 43661 5644
rect 43696 5635 43702 5687
rect 43754 5675 43760 5687
rect 44371 5678 44429 5684
rect 44371 5675 44383 5678
rect 43754 5647 44383 5675
rect 43754 5635 43760 5647
rect 44371 5644 44383 5647
rect 44417 5644 44429 5678
rect 44371 5638 44429 5644
rect 44656 5635 44662 5687
rect 44714 5675 44720 5687
rect 45139 5678 45197 5684
rect 45139 5675 45151 5678
rect 44714 5647 45151 5675
rect 44714 5635 44720 5647
rect 45139 5644 45151 5647
rect 45185 5644 45197 5678
rect 45139 5638 45197 5644
rect 46096 5635 46102 5687
rect 46154 5675 46160 5687
rect 46579 5678 46637 5684
rect 46579 5675 46591 5678
rect 46154 5647 46591 5675
rect 46154 5635 46160 5647
rect 46579 5644 46591 5647
rect 46625 5644 46637 5678
rect 46579 5638 46637 5644
rect 46672 5635 46678 5687
rect 46730 5675 46736 5687
rect 47347 5678 47405 5684
rect 47347 5675 47359 5678
rect 46730 5647 47359 5675
rect 46730 5635 46736 5647
rect 47347 5644 47359 5647
rect 47393 5644 47405 5678
rect 47347 5638 47405 5644
rect 47536 5635 47542 5687
rect 47594 5675 47600 5687
rect 48115 5678 48173 5684
rect 48115 5675 48127 5678
rect 47594 5647 48127 5675
rect 47594 5635 47600 5647
rect 48115 5644 48127 5647
rect 48161 5644 48173 5678
rect 48976 5675 48982 5687
rect 48937 5647 48982 5675
rect 48115 5638 48173 5644
rect 48976 5635 48982 5647
rect 49034 5635 49040 5687
rect 49648 5675 49654 5687
rect 49609 5647 49654 5675
rect 49648 5635 49654 5647
rect 49706 5635 49712 5687
rect 50515 5678 50573 5684
rect 50515 5644 50527 5678
rect 50561 5675 50573 5678
rect 50704 5675 50710 5687
rect 50561 5647 50710 5675
rect 50561 5644 50573 5647
rect 50515 5638 50573 5644
rect 50704 5635 50710 5647
rect 50762 5635 50768 5687
rect 52144 5675 52150 5687
rect 52105 5647 52150 5675
rect 52144 5635 52150 5647
rect 52202 5635 52208 5687
rect 52528 5635 52534 5687
rect 52586 5675 52592 5687
rect 52915 5678 52973 5684
rect 52915 5675 52927 5678
rect 52586 5647 52927 5675
rect 52586 5635 52592 5647
rect 52915 5644 52927 5647
rect 52961 5644 52973 5678
rect 53680 5675 53686 5687
rect 53641 5647 53686 5675
rect 52915 5638 52973 5644
rect 53680 5635 53686 5647
rect 53738 5635 53744 5687
rect 54451 5678 54509 5684
rect 54451 5644 54463 5678
rect 54497 5644 54509 5678
rect 54451 5638 54509 5644
rect 55987 5678 56045 5684
rect 55987 5644 55999 5678
rect 56033 5644 56045 5678
rect 57424 5675 57430 5687
rect 57385 5647 57430 5675
rect 55987 5638 56045 5644
rect 37514 5573 38366 5601
rect 37514 5561 37520 5573
rect 53584 5561 53590 5613
rect 53642 5601 53648 5613
rect 54466 5601 54494 5638
rect 53642 5573 54494 5601
rect 56002 5601 56030 5638
rect 57424 5635 57430 5647
rect 57482 5635 57488 5687
rect 59632 5601 59638 5613
rect 56002 5573 59638 5601
rect 53642 5561 53648 5573
rect 59632 5561 59638 5573
rect 59690 5561 59696 5613
rect 9922 5499 12974 5527
rect 21619 5530 21677 5536
rect 7658 5487 7664 5499
rect 21619 5496 21631 5530
rect 21665 5527 21677 5530
rect 21712 5527 21718 5539
rect 21665 5499 21718 5527
rect 21665 5496 21677 5499
rect 21619 5490 21677 5496
rect 21712 5487 21718 5499
rect 21770 5487 21776 5539
rect 26032 5487 26038 5539
rect 26090 5527 26096 5539
rect 26611 5530 26669 5536
rect 26611 5527 26623 5530
rect 26090 5499 26623 5527
rect 26090 5487 26096 5499
rect 26611 5496 26623 5499
rect 26657 5496 26669 5530
rect 38992 5527 38998 5539
rect 26611 5490 26669 5496
rect 27346 5499 38998 5527
rect 6160 5413 6166 5465
rect 6218 5453 6224 5465
rect 11539 5456 11597 5462
rect 11539 5453 11551 5456
rect 6218 5425 11551 5453
rect 6218 5413 6224 5425
rect 11539 5422 11551 5425
rect 11585 5422 11597 5456
rect 11539 5416 11597 5422
rect 17776 5413 17782 5465
rect 17834 5453 17840 5465
rect 27346 5453 27374 5499
rect 38992 5487 38998 5499
rect 39050 5487 39056 5539
rect 17834 5425 27374 5453
rect 17834 5413 17840 5425
rect 30640 5413 30646 5465
rect 30698 5453 30704 5465
rect 55411 5456 55469 5462
rect 55411 5453 55423 5456
rect 30698 5425 55423 5453
rect 30698 5413 30704 5425
rect 55411 5422 55423 5425
rect 55457 5422 55469 5456
rect 55411 5416 55469 5422
rect 1152 5354 58848 5376
rect 1152 5302 4294 5354
rect 4346 5302 4358 5354
rect 4410 5302 4422 5354
rect 4474 5302 4486 5354
rect 4538 5302 35014 5354
rect 35066 5302 35078 5354
rect 35130 5302 35142 5354
rect 35194 5302 35206 5354
rect 35258 5302 58848 5354
rect 1152 5280 58848 5302
rect 4720 5191 4726 5243
rect 4778 5231 4784 5243
rect 7507 5234 7565 5240
rect 7507 5231 7519 5234
rect 4778 5203 7519 5231
rect 4778 5191 4784 5203
rect 7507 5200 7519 5203
rect 7553 5231 7565 5234
rect 7699 5234 7757 5240
rect 7699 5231 7711 5234
rect 7553 5203 7711 5231
rect 7553 5200 7565 5203
rect 7507 5194 7565 5200
rect 7699 5200 7711 5203
rect 7745 5200 7757 5234
rect 7699 5194 7757 5200
rect 8467 5234 8525 5240
rect 8467 5200 8479 5234
rect 8513 5231 8525 5234
rect 8513 5203 8654 5231
rect 8513 5200 8525 5203
rect 8467 5194 8525 5200
rect 8626 5143 8654 5203
rect 57136 5191 57142 5243
rect 57194 5231 57200 5243
rect 58003 5234 58061 5240
rect 58003 5231 58015 5234
rect 57194 5203 58015 5231
rect 57194 5191 57200 5203
rect 58003 5200 58015 5203
rect 58049 5200 58061 5234
rect 58003 5194 58061 5200
rect 304 4969 310 5021
rect 362 5009 368 5021
rect 1555 5012 1613 5018
rect 1555 5009 1567 5012
rect 362 4981 1567 5009
rect 362 4969 368 4981
rect 1555 4978 1567 4981
rect 1601 4978 1613 5012
rect 1555 4972 1613 4978
rect 1840 4969 1846 5021
rect 1898 5009 1904 5021
rect 2323 5012 2381 5018
rect 2323 5009 2335 5012
rect 1898 4981 2335 5009
rect 1898 4969 1904 4981
rect 2323 4978 2335 4981
rect 2369 4978 2381 5012
rect 3088 5009 3094 5021
rect 3049 4981 3094 5009
rect 2323 4972 2381 4978
rect 3088 4969 3094 4981
rect 3146 4969 3152 5021
rect 4144 5009 4150 5021
rect 4105 4981 4150 5009
rect 4144 4969 4150 4981
rect 4202 4969 4208 5021
rect 5392 5009 5398 5021
rect 5353 4981 5398 5009
rect 5392 4969 5398 4981
rect 5450 4969 5456 5021
rect 6064 4969 6070 5021
rect 6122 5009 6128 5021
rect 6931 5012 6989 5018
rect 6931 5009 6943 5012
rect 6122 4981 6943 5009
rect 6122 4969 6128 4981
rect 6931 4978 6943 4981
rect 6977 4978 6989 5012
rect 9232 5009 9238 5021
rect 9193 4981 9238 5009
rect 6931 4972 6989 4978
rect 9232 4969 9238 4981
rect 9290 4969 9296 5021
rect 10000 5009 10006 5021
rect 9961 4981 10006 5009
rect 10000 4969 10006 4981
rect 10058 4969 10064 5021
rect 10672 4969 10678 5021
rect 10730 5009 10736 5021
rect 10771 5012 10829 5018
rect 10771 5009 10783 5012
rect 10730 4981 10783 5009
rect 10730 4969 10736 4981
rect 10771 4978 10783 4981
rect 10817 4978 10829 5012
rect 10771 4972 10829 4978
rect 11824 4969 11830 5021
rect 11882 5009 11888 5021
rect 12211 5012 12269 5018
rect 12211 5009 12223 5012
rect 11882 4981 12223 5009
rect 11882 4969 11888 4981
rect 12211 4978 12223 4981
rect 12257 4978 12269 5012
rect 12976 5009 12982 5021
rect 12937 4981 12982 5009
rect 12211 4972 12269 4978
rect 12976 4969 12982 4981
rect 13034 4969 13040 5021
rect 13936 5009 13942 5021
rect 13897 4981 13942 5009
rect 13936 4969 13942 4981
rect 13994 4969 14000 5021
rect 14416 4969 14422 5021
rect 14474 5009 14480 5021
rect 14707 5012 14765 5018
rect 14707 5009 14719 5012
rect 14474 4981 14719 5009
rect 14474 4969 14480 4981
rect 14707 4978 14719 4981
rect 14753 4978 14765 5012
rect 14707 4972 14765 4978
rect 14800 4969 14806 5021
rect 14858 5009 14864 5021
rect 15475 5012 15533 5018
rect 15475 5009 15487 5012
rect 14858 4981 15487 5009
rect 14858 4969 14864 4981
rect 15475 4978 15487 4981
rect 15521 4978 15533 5012
rect 15475 4972 15533 4978
rect 16339 5012 16397 5018
rect 16339 4978 16351 5012
rect 16385 5009 16397 5012
rect 16528 5009 16534 5021
rect 16385 4981 16534 5009
rect 16385 4978 16397 4981
rect 16339 4972 16397 4978
rect 16528 4969 16534 4981
rect 16586 4969 16592 5021
rect 17488 5009 17494 5021
rect 17449 4981 17494 5009
rect 17488 4969 17494 4981
rect 17546 4969 17552 5021
rect 17968 4969 17974 5021
rect 18026 5009 18032 5021
rect 18259 5012 18317 5018
rect 18259 5009 18271 5012
rect 18026 4981 18271 5009
rect 18026 4969 18032 4981
rect 18259 4978 18271 4981
rect 18305 4978 18317 5012
rect 19024 5009 19030 5021
rect 18985 4981 19030 5009
rect 18259 4972 18317 4978
rect 19024 4969 19030 4981
rect 19082 4969 19088 5021
rect 19120 4969 19126 5021
rect 19178 5009 19184 5021
rect 19795 5012 19853 5018
rect 19795 5009 19807 5012
rect 19178 4981 19807 5009
rect 19178 4969 19184 4981
rect 19795 4978 19807 4981
rect 19841 4978 19853 5012
rect 20656 5009 20662 5021
rect 20617 4981 20662 5009
rect 19795 4972 19853 4978
rect 20656 4969 20662 4981
rect 20714 4969 20720 5021
rect 20848 4969 20854 5021
rect 20906 5009 20912 5021
rect 21331 5012 21389 5018
rect 21331 5009 21343 5012
rect 20906 4981 21343 5009
rect 20906 4969 20912 4981
rect 21331 4978 21343 4981
rect 21377 4978 21389 5012
rect 22768 5009 22774 5021
rect 22729 4981 22774 5009
rect 21331 4972 21389 4978
rect 22768 4969 22774 4981
rect 22826 4969 22832 5021
rect 23536 5009 23542 5021
rect 23497 4981 23542 5009
rect 23536 4969 23542 4981
rect 23594 4969 23600 5021
rect 24307 5012 24365 5018
rect 24307 4978 24319 5012
rect 24353 4978 24365 5012
rect 25072 5009 25078 5021
rect 25033 4981 25078 5009
rect 24307 4972 24365 4978
rect 7942 4947 7994 4953
rect 23152 4895 23158 4947
rect 23210 4935 23216 4947
rect 24322 4935 24350 4972
rect 25072 4969 25078 4981
rect 25130 4969 25136 5021
rect 25843 5012 25901 5018
rect 25843 4978 25855 5012
rect 25889 4978 25901 5012
rect 26608 5009 26614 5021
rect 26569 4981 26614 5009
rect 25843 4972 25901 4978
rect 23210 4907 24350 4935
rect 23210 4895 23216 4907
rect 24880 4895 24886 4947
rect 24938 4935 24944 4947
rect 25858 4935 25886 4972
rect 26608 4969 26614 4981
rect 26666 4969 26672 5021
rect 28048 5009 28054 5021
rect 28009 4981 28054 5009
rect 28048 4969 28054 4981
rect 28106 4969 28112 5021
rect 28912 5009 28918 5021
rect 28873 4981 28918 5009
rect 28912 4969 28918 4981
rect 28970 4969 28976 5021
rect 29296 4969 29302 5021
rect 29354 5009 29360 5021
rect 29587 5012 29645 5018
rect 29587 5009 29599 5012
rect 29354 4981 29599 5009
rect 29354 4969 29360 4981
rect 29587 4978 29599 4981
rect 29633 4978 29645 5012
rect 30352 5009 30358 5021
rect 30313 4981 30358 5009
rect 29587 4972 29645 4978
rect 30352 4969 30358 4981
rect 30410 4969 30416 5021
rect 31120 5009 31126 5021
rect 31081 4981 31126 5009
rect 31120 4969 31126 4981
rect 31178 4969 31184 5021
rect 31888 5009 31894 5021
rect 31849 4981 31894 5009
rect 31888 4969 31894 4981
rect 31946 4969 31952 5021
rect 33328 5009 33334 5021
rect 33289 4981 33334 5009
rect 33328 4969 33334 4981
rect 33386 4969 33392 5021
rect 34096 5009 34102 5021
rect 34057 4981 34102 5009
rect 34096 4969 34102 4981
rect 34154 4969 34160 5021
rect 34864 5009 34870 5021
rect 34825 4981 34870 5009
rect 34864 4969 34870 4981
rect 34922 4969 34928 5021
rect 35344 4969 35350 5021
rect 35402 5009 35408 5021
rect 35635 5012 35693 5018
rect 35635 5009 35647 5012
rect 35402 4981 35647 5009
rect 35402 4969 35408 4981
rect 35635 4978 35647 4981
rect 35681 4978 35693 5012
rect 35635 4972 35693 4978
rect 36112 4969 36118 5021
rect 36170 5009 36176 5021
rect 36403 5012 36461 5018
rect 36403 5009 36415 5012
rect 36170 4981 36415 5009
rect 36170 4969 36176 4981
rect 36403 4978 36415 4981
rect 36449 4978 36461 5012
rect 36403 4972 36461 4978
rect 36880 4969 36886 5021
rect 36938 5009 36944 5021
rect 37171 5012 37229 5018
rect 37171 5009 37183 5012
rect 36938 4981 37183 5009
rect 36938 4969 36944 4981
rect 37171 4978 37183 4981
rect 37217 4978 37229 5012
rect 38608 5009 38614 5021
rect 38569 4981 38614 5009
rect 37171 4972 37229 4978
rect 38608 4969 38614 4981
rect 38666 4969 38672 5021
rect 39376 5009 39382 5021
rect 39337 4981 39382 5009
rect 39376 4969 39382 4981
rect 39434 4969 39440 5021
rect 39568 4969 39574 5021
rect 39626 5009 39632 5021
rect 40147 5012 40205 5018
rect 40147 5009 40159 5012
rect 39626 4981 40159 5009
rect 39626 4969 39632 4981
rect 40147 4978 40159 4981
rect 40193 4978 40205 5012
rect 40912 5009 40918 5021
rect 40873 4981 40918 5009
rect 40147 4972 40205 4978
rect 40912 4969 40918 4981
rect 40970 4969 40976 5021
rect 41680 5009 41686 5021
rect 41641 4981 41686 5009
rect 41680 4969 41686 4981
rect 41738 4969 41744 5021
rect 42160 4969 42166 5021
rect 42218 5009 42224 5021
rect 42451 5012 42509 5018
rect 42451 5009 42463 5012
rect 42218 4981 42463 5009
rect 42218 4969 42224 4981
rect 42451 4978 42463 4981
rect 42497 4978 42509 5012
rect 42451 4972 42509 4978
rect 43312 4969 43318 5021
rect 43370 5009 43376 5021
rect 43891 5012 43949 5018
rect 43891 5009 43903 5012
rect 43370 4981 43903 5009
rect 43370 4969 43376 4981
rect 43891 4978 43903 4981
rect 43937 4978 43949 5012
rect 43891 4972 43949 4978
rect 44755 5012 44813 5018
rect 44755 4978 44767 5012
rect 44801 5009 44813 5012
rect 44848 5009 44854 5021
rect 44801 4981 44854 5009
rect 44801 4978 44813 4981
rect 44755 4972 44813 4978
rect 44848 4969 44854 4981
rect 44906 4969 44912 5021
rect 45424 5009 45430 5021
rect 45385 4981 45430 5009
rect 45424 4969 45430 4981
rect 45482 4969 45488 5021
rect 46192 5009 46198 5021
rect 46153 4981 46198 5009
rect 46192 4969 46198 4981
rect 46250 4969 46256 5021
rect 46288 4969 46294 5021
rect 46346 5009 46352 5021
rect 46963 5012 47021 5018
rect 46963 5009 46975 5012
rect 46346 4981 46975 5009
rect 46346 4969 46352 4981
rect 46963 4978 46975 4981
rect 47009 4978 47021 5012
rect 46963 4972 47021 4978
rect 47632 4969 47638 5021
rect 47690 5009 47696 5021
rect 47731 5012 47789 5018
rect 47731 5009 47743 5012
rect 47690 4981 47743 5009
rect 47690 4969 47696 4981
rect 47731 4978 47743 4981
rect 47777 4978 47789 5012
rect 49360 5009 49366 5021
rect 49321 4981 49366 5009
rect 47731 4972 47789 4978
rect 49360 4969 49366 4981
rect 49418 4969 49424 5021
rect 50416 5009 50422 5021
rect 50377 4981 50422 5009
rect 50416 4969 50422 4981
rect 50474 4969 50480 5021
rect 50896 4969 50902 5021
rect 50954 5009 50960 5021
rect 51091 5012 51149 5018
rect 51091 5009 51103 5012
rect 50954 4981 51103 5009
rect 50954 4969 50960 4981
rect 51091 4978 51103 4981
rect 51137 4978 51149 5012
rect 51856 5009 51862 5021
rect 51817 4981 51862 5009
rect 51091 4972 51149 4978
rect 51856 4969 51862 4981
rect 51914 4969 51920 5021
rect 52240 4969 52246 5021
rect 52298 5009 52304 5021
rect 52627 5012 52685 5018
rect 52627 5009 52639 5012
rect 52298 4981 52639 5009
rect 52298 4969 52304 4981
rect 52627 4978 52639 4981
rect 52673 4978 52685 5012
rect 52627 4972 52685 4978
rect 53296 4969 53302 5021
rect 53354 5009 53360 5021
rect 54451 5012 54509 5018
rect 54451 5009 54463 5012
rect 53354 4981 54463 5009
rect 53354 4969 53360 4981
rect 54451 4978 54463 4981
rect 54497 4978 54509 5012
rect 54451 4972 54509 4978
rect 55603 5012 55661 5018
rect 55603 4978 55615 5012
rect 55649 4978 55661 5012
rect 55603 4972 55661 4978
rect 56371 5012 56429 5018
rect 56371 4978 56383 5012
rect 56417 4978 56429 5012
rect 57040 5009 57046 5021
rect 57001 4981 57046 5009
rect 56371 4972 56429 4978
rect 24938 4907 25886 4935
rect 24938 4895 24944 4907
rect 7942 4889 7994 4895
rect 8368 4861 8374 4873
rect 8256 4833 8374 4861
rect 8368 4821 8374 4833
rect 8426 4821 8432 4873
rect 55618 4861 55646 4972
rect 56386 4935 56414 4972
rect 57040 4969 57046 4981
rect 57098 4969 57104 5021
rect 57808 4935 57814 4947
rect 56386 4907 57814 4935
rect 57808 4895 57814 4907
rect 57866 4895 57872 4947
rect 59248 4861 59254 4873
rect 55618 4833 59254 4861
rect 59248 4821 59254 4833
rect 59306 4821 59312 4873
rect 1152 4688 58848 4710
rect 1152 4636 19654 4688
rect 19706 4636 19718 4688
rect 19770 4636 19782 4688
rect 19834 4636 19846 4688
rect 19898 4636 50374 4688
rect 50426 4636 50438 4688
rect 50490 4636 50502 4688
rect 50554 4636 50566 4688
rect 50618 4636 58848 4688
rect 1152 4614 58848 4636
rect 784 4377 790 4429
rect 842 4417 848 4429
rect 842 4389 2366 4417
rect 842 4377 848 4389
rect 1168 4303 1174 4355
rect 1226 4343 1232 4355
rect 2338 4352 2366 4389
rect 14032 4377 14038 4429
rect 14090 4417 14096 4429
rect 41107 4420 41165 4426
rect 41107 4417 41119 4420
rect 14090 4389 41119 4417
rect 14090 4377 14096 4389
rect 41107 4386 41119 4389
rect 41153 4417 41165 4420
rect 41299 4420 41357 4426
rect 41299 4417 41311 4420
rect 41153 4389 41311 4417
rect 41153 4386 41165 4389
rect 41107 4380 41165 4386
rect 41299 4386 41311 4389
rect 41345 4386 41357 4420
rect 41299 4380 41357 4386
rect 1555 4346 1613 4352
rect 1555 4343 1567 4346
rect 1226 4315 1567 4343
rect 1226 4303 1232 4315
rect 1555 4312 1567 4315
rect 1601 4312 1613 4346
rect 1555 4306 1613 4312
rect 2323 4346 2381 4352
rect 2323 4312 2335 4346
rect 2369 4312 2381 4346
rect 3091 4346 3149 4352
rect 3091 4343 3103 4346
rect 2323 4306 2381 4312
rect 2866 4315 3103 4343
rect 1360 4229 1366 4281
rect 1418 4269 1424 4281
rect 2866 4269 2894 4315
rect 3091 4312 3103 4315
rect 3137 4312 3149 4346
rect 3091 4306 3149 4312
rect 4339 4346 4397 4352
rect 4339 4312 4351 4346
rect 4385 4312 4397 4346
rect 4339 4306 4397 4312
rect 1418 4241 2894 4269
rect 1418 4229 1424 4241
rect 3760 4229 3766 4281
rect 3818 4269 3824 4281
rect 4354 4269 4382 4306
rect 4720 4303 4726 4355
rect 4778 4343 4784 4355
rect 5107 4346 5165 4352
rect 5107 4343 5119 4346
rect 4778 4315 5119 4343
rect 4778 4303 4784 4315
rect 5107 4312 5119 4315
rect 5153 4312 5165 4346
rect 5875 4346 5933 4352
rect 5875 4343 5887 4346
rect 5107 4306 5165 4312
rect 5602 4315 5887 4343
rect 3818 4241 4382 4269
rect 3818 4229 3824 4241
rect 5008 4229 5014 4281
rect 5066 4269 5072 4281
rect 5602 4269 5630 4315
rect 5875 4312 5887 4315
rect 5921 4312 5933 4346
rect 5875 4306 5933 4312
rect 6643 4346 6701 4352
rect 6643 4312 6655 4346
rect 6689 4312 6701 4346
rect 7408 4343 7414 4355
rect 7369 4315 7414 4343
rect 6643 4306 6701 4312
rect 5066 4241 5630 4269
rect 5066 4229 5072 4241
rect 5680 4229 5686 4281
rect 5738 4269 5744 4281
rect 6658 4269 6686 4306
rect 7408 4303 7414 4315
rect 7466 4303 7472 4355
rect 8179 4346 8237 4352
rect 8179 4312 8191 4346
rect 8225 4312 8237 4346
rect 9616 4343 9622 4355
rect 9577 4315 9622 4343
rect 8179 4306 8237 4312
rect 5738 4241 6686 4269
rect 5738 4229 5744 4241
rect 3472 4155 3478 4207
rect 3530 4195 3536 4207
rect 4912 4195 4918 4207
rect 3530 4167 4918 4195
rect 3530 4155 3536 4167
rect 4912 4155 4918 4167
rect 4970 4155 4976 4207
rect 6448 4155 6454 4207
rect 6506 4195 6512 4207
rect 8194 4195 8222 4306
rect 9616 4303 9622 4315
rect 9674 4303 9680 4355
rect 10384 4343 10390 4355
rect 10345 4315 10390 4343
rect 10384 4303 10390 4315
rect 10442 4303 10448 4355
rect 10768 4303 10774 4355
rect 10826 4343 10832 4355
rect 11155 4346 11213 4352
rect 11155 4343 11167 4346
rect 10826 4315 11167 4343
rect 10826 4303 10832 4315
rect 11155 4312 11167 4315
rect 11201 4312 11213 4346
rect 11155 4306 11213 4312
rect 11923 4346 11981 4352
rect 11923 4312 11935 4346
rect 11969 4312 11981 4346
rect 11923 4306 11981 4312
rect 12691 4346 12749 4352
rect 12691 4312 12703 4346
rect 12737 4312 12749 4346
rect 13552 4343 13558 4355
rect 13513 4315 13558 4343
rect 12691 4306 12749 4312
rect 9808 4229 9814 4281
rect 9866 4269 9872 4281
rect 10192 4269 10198 4281
rect 9866 4241 10198 4269
rect 9866 4229 9872 4241
rect 10192 4229 10198 4241
rect 10250 4229 10256 4281
rect 6506 4167 8222 4195
rect 6506 4155 6512 4167
rect 11152 4155 11158 4207
rect 11210 4195 11216 4207
rect 11938 4195 11966 4306
rect 11210 4167 11966 4195
rect 11210 4155 11216 4167
rect 3952 4081 3958 4133
rect 4010 4121 4016 4133
rect 5104 4121 5110 4133
rect 4010 4093 5110 4121
rect 4010 4081 4016 4093
rect 5104 4081 5110 4093
rect 5162 4081 5168 4133
rect 9040 4081 9046 4133
rect 9098 4121 9104 4133
rect 10672 4121 10678 4133
rect 9098 4093 10678 4121
rect 9098 4081 9104 4093
rect 10672 4081 10678 4093
rect 10730 4081 10736 4133
rect 11440 4081 11446 4133
rect 11498 4121 11504 4133
rect 12706 4121 12734 4306
rect 13552 4303 13558 4315
rect 13610 4303 13616 4355
rect 15472 4343 15478 4355
rect 15433 4315 15478 4343
rect 15472 4303 15478 4315
rect 15530 4303 15536 4355
rect 15952 4303 15958 4355
rect 16010 4343 16016 4355
rect 16243 4346 16301 4352
rect 16243 4343 16255 4346
rect 16010 4315 16255 4343
rect 16010 4303 16016 4315
rect 16243 4312 16255 4315
rect 16289 4312 16301 4346
rect 16243 4306 16301 4312
rect 16432 4303 16438 4355
rect 16490 4343 16496 4355
rect 17011 4346 17069 4352
rect 17011 4343 17023 4346
rect 16490 4315 17023 4343
rect 16490 4303 16496 4315
rect 17011 4312 17023 4315
rect 17057 4312 17069 4346
rect 17779 4346 17837 4352
rect 17779 4343 17791 4346
rect 17011 4306 17069 4312
rect 17266 4315 17791 4343
rect 16912 4229 16918 4281
rect 16970 4269 16976 4281
rect 17266 4269 17294 4315
rect 17779 4312 17791 4315
rect 17825 4312 17837 4346
rect 17779 4306 17837 4312
rect 18547 4346 18605 4352
rect 18547 4312 18559 4346
rect 18593 4312 18605 4346
rect 20272 4343 20278 4355
rect 20233 4315 20278 4343
rect 18547 4306 18605 4312
rect 16970 4241 17294 4269
rect 16970 4229 16976 4241
rect 17584 4229 17590 4281
rect 17642 4269 17648 4281
rect 18562 4269 18590 4306
rect 20272 4303 20278 4315
rect 20330 4303 20336 4355
rect 21040 4343 21046 4355
rect 21001 4315 21046 4343
rect 21040 4303 21046 4315
rect 21098 4303 21104 4355
rect 21808 4343 21814 4355
rect 21769 4315 21814 4343
rect 21808 4303 21814 4315
rect 21866 4303 21872 4355
rect 23248 4343 23254 4355
rect 23209 4315 23254 4343
rect 23248 4303 23254 4315
rect 23306 4303 23312 4355
rect 24019 4346 24077 4352
rect 24019 4312 24031 4346
rect 24065 4312 24077 4346
rect 25456 4343 25462 4355
rect 25417 4315 25462 4343
rect 24019 4306 24077 4312
rect 17642 4241 18590 4269
rect 17642 4229 17648 4241
rect 22000 4229 22006 4281
rect 22058 4269 22064 4281
rect 24034 4269 24062 4306
rect 25456 4303 25462 4315
rect 25514 4303 25520 4355
rect 26128 4303 26134 4355
rect 26186 4343 26192 4355
rect 26227 4346 26285 4352
rect 26227 4343 26239 4346
rect 26186 4315 26239 4343
rect 26186 4303 26192 4315
rect 26227 4312 26239 4315
rect 26273 4312 26285 4346
rect 26227 4306 26285 4312
rect 26512 4303 26518 4355
rect 26570 4343 26576 4355
rect 26995 4346 27053 4352
rect 26995 4343 27007 4346
rect 26570 4315 27007 4343
rect 26570 4303 26576 4315
rect 26995 4312 27007 4315
rect 27041 4312 27053 4346
rect 28336 4343 28342 4355
rect 28297 4315 28342 4343
rect 26995 4306 27053 4312
rect 28336 4303 28342 4315
rect 28394 4303 28400 4355
rect 29104 4343 29110 4355
rect 29065 4315 29110 4343
rect 29104 4303 29110 4315
rect 29162 4303 29168 4355
rect 30928 4343 30934 4355
rect 30889 4315 30934 4343
rect 30928 4303 30934 4315
rect 30986 4303 30992 4355
rect 31696 4343 31702 4355
rect 31657 4315 31702 4343
rect 31696 4303 31702 4315
rect 31754 4303 31760 4355
rect 32752 4343 32758 4355
rect 32713 4315 32758 4343
rect 32752 4303 32758 4315
rect 32810 4303 32816 4355
rect 33904 4343 33910 4355
rect 33865 4315 33910 4343
rect 33904 4303 33910 4315
rect 33962 4303 33968 4355
rect 34576 4303 34582 4355
rect 34634 4343 34640 4355
rect 34675 4346 34733 4352
rect 34675 4343 34687 4346
rect 34634 4315 34687 4343
rect 34634 4303 34640 4315
rect 34675 4312 34687 4315
rect 34721 4312 34733 4346
rect 36019 4346 36077 4352
rect 36019 4343 36031 4346
rect 34675 4306 34733 4312
rect 34786 4315 36031 4343
rect 22058 4241 24062 4269
rect 22058 4229 22064 4241
rect 34192 4229 34198 4281
rect 34250 4269 34256 4281
rect 34786 4269 34814 4315
rect 36019 4312 36031 4315
rect 36065 4312 36077 4346
rect 36784 4343 36790 4355
rect 36745 4315 36790 4343
rect 36019 4306 36077 4312
rect 36784 4303 36790 4315
rect 36842 4303 36848 4355
rect 37555 4346 37613 4352
rect 37555 4343 37567 4346
rect 37426 4315 37567 4343
rect 34250 4241 34814 4269
rect 34250 4229 34256 4241
rect 37168 4229 37174 4281
rect 37226 4269 37232 4281
rect 37426 4269 37454 4315
rect 37555 4312 37567 4315
rect 37601 4312 37613 4346
rect 38992 4343 38998 4355
rect 38953 4315 38998 4343
rect 37555 4306 37613 4312
rect 38992 4303 38998 4315
rect 39050 4303 39056 4355
rect 39760 4343 39766 4355
rect 39721 4315 39766 4343
rect 39760 4303 39766 4315
rect 39818 4303 39824 4355
rect 41968 4343 41974 4355
rect 41929 4315 41974 4343
rect 41968 4303 41974 4315
rect 42026 4303 42032 4355
rect 42352 4303 42358 4355
rect 42410 4343 42416 4355
rect 42739 4346 42797 4352
rect 42739 4343 42751 4346
rect 42410 4315 42751 4343
rect 42410 4303 42416 4315
rect 42739 4312 42751 4315
rect 42785 4312 42797 4346
rect 42739 4306 42797 4312
rect 43408 4303 43414 4355
rect 43466 4343 43472 4355
rect 43507 4346 43565 4352
rect 43507 4343 43519 4346
rect 43466 4315 43519 4343
rect 43466 4303 43472 4315
rect 43507 4312 43519 4315
rect 43553 4312 43565 4346
rect 44944 4343 44950 4355
rect 44905 4315 44950 4343
rect 43507 4306 43565 4312
rect 44944 4303 44950 4315
rect 45002 4303 45008 4355
rect 46768 4343 46774 4355
rect 46729 4315 46774 4343
rect 46768 4303 46774 4315
rect 46826 4303 46832 4355
rect 47539 4346 47597 4352
rect 47539 4312 47551 4346
rect 47585 4312 47597 4346
rect 47539 4306 47597 4312
rect 37226 4241 37454 4269
rect 37226 4229 37232 4241
rect 47440 4229 47446 4281
rect 47498 4269 47504 4281
rect 47554 4269 47582 4306
rect 47824 4303 47830 4355
rect 47882 4343 47888 4355
rect 48307 4346 48365 4352
rect 48307 4343 48319 4346
rect 47882 4315 48319 4343
rect 47882 4303 47888 4315
rect 48307 4312 48319 4315
rect 48353 4312 48365 4346
rect 48307 4306 48365 4312
rect 49075 4346 49133 4352
rect 49075 4312 49087 4346
rect 49121 4312 49133 4346
rect 49840 4343 49846 4355
rect 49801 4315 49846 4343
rect 49075 4306 49133 4312
rect 47498 4241 47582 4269
rect 47498 4229 47504 4241
rect 48592 4229 48598 4281
rect 48650 4269 48656 4281
rect 49090 4269 49118 4306
rect 49840 4303 49846 4315
rect 49898 4303 49904 4355
rect 50611 4346 50669 4352
rect 50611 4312 50623 4346
rect 50657 4312 50669 4346
rect 50611 4306 50669 4312
rect 51859 4346 51917 4352
rect 51859 4312 51871 4346
rect 51905 4312 51917 4346
rect 52624 4343 52630 4355
rect 52585 4315 52630 4343
rect 51859 4306 51917 4312
rect 48650 4241 49118 4269
rect 48650 4229 48656 4241
rect 49936 4229 49942 4281
rect 49994 4269 50000 4281
rect 50626 4269 50654 4306
rect 49994 4241 50654 4269
rect 49994 4229 50000 4241
rect 50992 4229 50998 4281
rect 51050 4269 51056 4281
rect 51874 4269 51902 4306
rect 52624 4303 52630 4315
rect 52682 4303 52688 4355
rect 53395 4346 53453 4352
rect 53395 4312 53407 4346
rect 53441 4312 53453 4346
rect 53395 4306 53453 4312
rect 51050 4241 51902 4269
rect 51050 4229 51056 4241
rect 53008 4229 53014 4281
rect 53066 4269 53072 4281
rect 53410 4269 53438 4306
rect 54064 4303 54070 4355
rect 54122 4343 54128 4355
rect 54163 4346 54221 4352
rect 54163 4343 54175 4346
rect 54122 4315 54175 4343
rect 54122 4303 54128 4315
rect 54163 4312 54175 4315
rect 54209 4312 54221 4346
rect 55600 4343 55606 4355
rect 55561 4315 55606 4343
rect 54163 4306 54221 4312
rect 55600 4303 55606 4315
rect 55658 4303 55664 4355
rect 56656 4303 56662 4355
rect 56714 4343 56720 4355
rect 57139 4346 57197 4352
rect 57139 4343 57151 4346
rect 56714 4315 57151 4343
rect 56714 4303 56720 4315
rect 57139 4312 57151 4315
rect 57185 4312 57197 4346
rect 57139 4306 57197 4312
rect 55120 4269 55126 4281
rect 53066 4241 53438 4269
rect 55081 4241 55126 4269
rect 53066 4229 53072 4241
rect 55120 4229 55126 4241
rect 55178 4229 55184 4281
rect 56368 4229 56374 4281
rect 56426 4269 56432 4281
rect 59440 4269 59446 4281
rect 56426 4241 59446 4269
rect 56426 4229 56432 4241
rect 59440 4229 59446 4241
rect 59498 4229 59504 4281
rect 43504 4155 43510 4207
rect 43562 4195 43568 4207
rect 44467 4198 44525 4204
rect 44467 4195 44479 4198
rect 43562 4167 44479 4195
rect 43562 4155 43568 4167
rect 44467 4164 44479 4167
rect 44513 4164 44525 4198
rect 44467 4158 44525 4164
rect 11498 4093 12734 4121
rect 11498 4081 11504 4093
rect 55888 4081 55894 4133
rect 55946 4121 55952 4133
rect 57904 4121 57910 4133
rect 55946 4093 57910 4121
rect 55946 4081 55952 4093
rect 57904 4081 57910 4093
rect 57962 4081 57968 4133
rect 1152 4022 58848 4044
rect 1152 3970 4294 4022
rect 4346 3970 4358 4022
rect 4410 3970 4422 4022
rect 4474 3970 4486 4022
rect 4538 3970 35014 4022
rect 35066 3970 35078 4022
rect 35130 3970 35142 4022
rect 35194 3970 35206 4022
rect 35258 3970 58848 4022
rect 1152 3948 58848 3970
rect 1936 3859 1942 3911
rect 1994 3899 2000 3911
rect 3280 3899 3286 3911
rect 1994 3871 3286 3899
rect 1994 3859 2000 3871
rect 3280 3859 3286 3871
rect 3338 3859 3344 3911
rect 7888 3859 7894 3911
rect 7946 3899 7952 3911
rect 9232 3899 9238 3911
rect 7946 3871 9238 3899
rect 7946 3859 7952 3871
rect 9232 3859 9238 3871
rect 9290 3859 9296 3911
rect 21232 3859 21238 3911
rect 21290 3899 21296 3911
rect 22768 3899 22774 3911
rect 21290 3871 22774 3899
rect 21290 3859 21296 3871
rect 22768 3859 22774 3871
rect 22826 3859 22832 3911
rect 29776 3899 29782 3911
rect 28834 3871 29782 3899
rect 28834 3837 28862 3871
rect 29776 3859 29782 3871
rect 29834 3859 29840 3911
rect 31984 3859 31990 3911
rect 32042 3899 32048 3911
rect 33520 3899 33526 3911
rect 32042 3871 33526 3899
rect 32042 3859 32048 3871
rect 33520 3859 33526 3871
rect 33578 3859 33584 3911
rect 35536 3859 35542 3911
rect 35594 3899 35600 3911
rect 39184 3899 39190 3911
rect 35594 3871 39190 3899
rect 35594 3859 35600 3871
rect 39184 3859 39190 3871
rect 39242 3859 39248 3911
rect 57328 3859 57334 3911
rect 57386 3899 57392 3911
rect 59152 3899 59158 3911
rect 57386 3871 59158 3899
rect 57386 3859 57392 3871
rect 59152 3859 59158 3871
rect 59210 3859 59216 3911
rect 496 3785 502 3837
rect 554 3825 560 3837
rect 1648 3825 1654 3837
rect 554 3797 1654 3825
rect 554 3785 560 3797
rect 1648 3785 1654 3797
rect 1706 3785 1712 3837
rect 2320 3785 2326 3837
rect 2378 3825 2384 3837
rect 3088 3825 3094 3837
rect 2378 3797 3094 3825
rect 2378 3785 2384 3797
rect 3088 3785 3094 3797
rect 3146 3785 3152 3837
rect 8272 3785 8278 3837
rect 8330 3825 8336 3837
rect 10000 3825 10006 3837
rect 8330 3797 10006 3825
rect 8330 3785 8336 3797
rect 10000 3785 10006 3797
rect 10058 3785 10064 3837
rect 16720 3785 16726 3837
rect 16778 3825 16784 3837
rect 17296 3825 17302 3837
rect 16778 3797 17302 3825
rect 16778 3785 16784 3797
rect 17296 3785 17302 3797
rect 17354 3785 17360 3837
rect 19408 3785 19414 3837
rect 19466 3825 19472 3837
rect 20656 3825 20662 3837
rect 19466 3797 20662 3825
rect 19466 3785 19472 3797
rect 20656 3785 20662 3797
rect 20714 3785 20720 3837
rect 22288 3785 22294 3837
rect 22346 3825 22352 3837
rect 23632 3825 23638 3837
rect 22346 3797 23638 3825
rect 22346 3785 22352 3797
rect 23632 3785 23638 3797
rect 23690 3785 23696 3837
rect 26416 3785 26422 3837
rect 26474 3825 26480 3837
rect 28048 3825 28054 3837
rect 26474 3797 28054 3825
rect 26474 3785 26480 3797
rect 28048 3785 28054 3797
rect 28106 3785 28112 3837
rect 28816 3785 28822 3837
rect 28874 3785 28880 3837
rect 29008 3785 29014 3837
rect 29066 3825 29072 3837
rect 30352 3825 30358 3837
rect 29066 3797 30358 3825
rect 29066 3785 29072 3797
rect 30352 3785 30358 3797
rect 30410 3785 30416 3837
rect 33424 3785 33430 3837
rect 33482 3825 33488 3837
rect 34864 3825 34870 3837
rect 33482 3797 34870 3825
rect 33482 3785 33488 3797
rect 34864 3785 34870 3797
rect 34922 3785 34928 3837
rect 37840 3785 37846 3837
rect 37898 3825 37904 3837
rect 39376 3825 39382 3837
rect 37898 3797 39382 3825
rect 37898 3785 37904 3797
rect 39376 3785 39382 3797
rect 39434 3785 39440 3837
rect 40048 3785 40054 3837
rect 40106 3825 40112 3837
rect 41680 3825 41686 3837
rect 40106 3797 41686 3825
rect 40106 3785 40112 3797
rect 41680 3785 41686 3797
rect 41738 3785 41744 3837
rect 49264 3785 49270 3837
rect 49322 3825 49328 3837
rect 50704 3825 50710 3837
rect 49322 3797 50710 3825
rect 49322 3785 49328 3797
rect 50704 3785 50710 3797
rect 50762 3785 50768 3837
rect 51280 3785 51286 3837
rect 51338 3785 51344 3837
rect 54352 3785 54358 3837
rect 54410 3825 54416 3837
rect 55216 3825 55222 3837
rect 54410 3797 55222 3825
rect 54410 3785 54416 3797
rect 55216 3785 55222 3797
rect 55274 3785 55280 3837
rect 57136 3785 57142 3837
rect 57194 3825 57200 3837
rect 57194 3797 57374 3825
rect 57194 3785 57200 3797
rect 5200 3751 5206 3763
rect 3202 3723 5206 3751
rect 112 3637 118 3689
rect 170 3677 176 3689
rect 1555 3680 1613 3686
rect 1555 3677 1567 3680
rect 170 3649 1567 3677
rect 170 3637 176 3649
rect 1555 3646 1567 3649
rect 1601 3646 1613 3680
rect 1555 3640 1613 3646
rect 1648 3637 1654 3689
rect 1706 3677 1712 3689
rect 2323 3680 2381 3686
rect 2323 3677 2335 3680
rect 1706 3649 2335 3677
rect 1706 3637 1712 3649
rect 2323 3646 2335 3649
rect 2369 3646 2381 3680
rect 2323 3640 2381 3646
rect 2704 3637 2710 3689
rect 2762 3677 2768 3689
rect 3091 3680 3149 3686
rect 3091 3677 3103 3680
rect 2762 3649 3103 3677
rect 2762 3637 2768 3649
rect 3091 3646 3103 3649
rect 3137 3646 3149 3680
rect 3091 3640 3149 3646
rect 976 3563 982 3615
rect 1034 3603 1040 3615
rect 2416 3603 2422 3615
rect 1034 3575 2422 3603
rect 1034 3563 1040 3575
rect 2416 3563 2422 3575
rect 2474 3563 2480 3615
rect 3202 3603 3230 3723
rect 5200 3711 5206 3723
rect 5258 3711 5264 3763
rect 24112 3711 24118 3763
rect 24170 3751 24176 3763
rect 24688 3751 24694 3763
rect 24170 3723 24694 3751
rect 24170 3711 24176 3723
rect 24688 3711 24694 3723
rect 24746 3711 24752 3763
rect 28720 3711 28726 3763
rect 28778 3751 28784 3763
rect 28778 3723 29630 3751
rect 28778 3711 28784 3723
rect 3859 3680 3917 3686
rect 3859 3646 3871 3680
rect 3905 3646 3917 3680
rect 3859 3640 3917 3646
rect 4627 3680 4685 3686
rect 4627 3646 4639 3680
rect 4673 3646 4685 3680
rect 5584 3677 5590 3689
rect 5545 3649 5590 3677
rect 4627 3640 4685 3646
rect 2866 3575 3230 3603
rect 592 3415 598 3467
rect 650 3455 656 3467
rect 1456 3455 1462 3467
rect 650 3427 1462 3455
rect 650 3415 656 3427
rect 1456 3415 1462 3427
rect 1514 3415 1520 3467
rect 2416 3415 2422 3467
rect 2474 3455 2480 3467
rect 2866 3455 2894 3575
rect 3088 3489 3094 3541
rect 3146 3529 3152 3541
rect 3874 3529 3902 3640
rect 3146 3501 3902 3529
rect 3146 3489 3152 3501
rect 2474 3427 2894 3455
rect 2474 3415 2480 3427
rect 3376 3415 3382 3467
rect 3434 3455 3440 3467
rect 4642 3455 4670 3640
rect 5584 3637 5590 3649
rect 5642 3637 5648 3689
rect 6352 3637 6358 3689
rect 6410 3677 6416 3689
rect 6931 3680 6989 3686
rect 6931 3677 6943 3680
rect 6410 3649 6943 3677
rect 6410 3637 6416 3649
rect 6931 3646 6943 3649
rect 6977 3646 6989 3680
rect 6931 3640 6989 3646
rect 7024 3637 7030 3689
rect 7082 3677 7088 3689
rect 7699 3680 7757 3686
rect 7699 3677 7711 3680
rect 7082 3649 7711 3677
rect 7082 3637 7088 3649
rect 7699 3646 7711 3649
rect 7745 3646 7757 3680
rect 7699 3640 7757 3646
rect 7792 3637 7798 3689
rect 7850 3677 7856 3689
rect 8467 3680 8525 3686
rect 8467 3677 8479 3680
rect 7850 3649 8479 3677
rect 7850 3637 7856 3649
rect 8467 3646 8479 3649
rect 8513 3646 8525 3680
rect 8467 3640 8525 3646
rect 8560 3637 8566 3689
rect 8618 3677 8624 3689
rect 9235 3680 9293 3686
rect 9235 3677 9247 3680
rect 8618 3649 9247 3677
rect 8618 3637 8624 3649
rect 9235 3646 9247 3649
rect 9281 3646 9293 3680
rect 9235 3640 9293 3646
rect 9328 3637 9334 3689
rect 9386 3677 9392 3689
rect 10003 3680 10061 3686
rect 10003 3677 10015 3680
rect 9386 3649 10015 3677
rect 9386 3637 9392 3649
rect 10003 3646 10015 3649
rect 10049 3646 10061 3680
rect 10003 3640 10061 3646
rect 10771 3680 10829 3686
rect 10771 3646 10783 3680
rect 10817 3646 10829 3680
rect 10771 3640 10829 3646
rect 12979 3680 13037 3686
rect 12979 3646 12991 3680
rect 13025 3677 13037 3680
rect 13168 3677 13174 3689
rect 13025 3649 13174 3677
rect 13025 3646 13037 3649
rect 12979 3640 13037 3646
rect 10000 3489 10006 3541
rect 10058 3529 10064 3541
rect 10786 3529 10814 3640
rect 13168 3637 13174 3649
rect 13226 3637 13232 3689
rect 13648 3677 13654 3689
rect 13609 3649 13654 3677
rect 13648 3637 13654 3649
rect 13706 3637 13712 3689
rect 14032 3637 14038 3689
rect 14090 3677 14096 3689
rect 14419 3680 14477 3686
rect 14419 3677 14431 3680
rect 14090 3649 14431 3677
rect 14090 3637 14096 3649
rect 14419 3646 14431 3649
rect 14465 3646 14477 3680
rect 14419 3640 14477 3646
rect 14800 3637 14806 3689
rect 14858 3677 14864 3689
rect 15187 3680 15245 3686
rect 15187 3677 15199 3680
rect 14858 3649 15199 3677
rect 14858 3637 14864 3649
rect 15187 3646 15199 3649
rect 15233 3646 15245 3680
rect 15187 3640 15245 3646
rect 15280 3637 15286 3689
rect 15338 3677 15344 3689
rect 15955 3680 16013 3686
rect 15955 3677 15967 3680
rect 15338 3649 15967 3677
rect 15338 3637 15344 3649
rect 15955 3646 15967 3649
rect 16001 3646 16013 3680
rect 15955 3640 16013 3646
rect 17392 3637 17398 3689
rect 17450 3677 17456 3689
rect 17491 3680 17549 3686
rect 17491 3677 17503 3680
rect 17450 3649 17503 3677
rect 17450 3637 17456 3649
rect 17491 3646 17503 3649
rect 17537 3646 17549 3680
rect 17491 3640 17549 3646
rect 18064 3637 18070 3689
rect 18122 3677 18128 3689
rect 18259 3680 18317 3686
rect 18259 3677 18271 3680
rect 18122 3649 18271 3677
rect 18122 3637 18128 3649
rect 18259 3646 18271 3649
rect 18305 3646 18317 3680
rect 18259 3640 18317 3646
rect 18448 3637 18454 3689
rect 18506 3677 18512 3689
rect 19027 3680 19085 3686
rect 19027 3677 19039 3680
rect 18506 3649 19039 3677
rect 18506 3637 18512 3649
rect 19027 3646 19039 3649
rect 19073 3646 19085 3680
rect 19027 3640 19085 3646
rect 19216 3637 19222 3689
rect 19274 3677 19280 3689
rect 19795 3680 19853 3686
rect 19795 3677 19807 3680
rect 19274 3649 19807 3677
rect 19274 3637 19280 3649
rect 19795 3646 19807 3649
rect 19841 3646 19853 3680
rect 19795 3640 19853 3646
rect 19984 3637 19990 3689
rect 20042 3677 20048 3689
rect 20563 3680 20621 3686
rect 20563 3677 20575 3680
rect 20042 3649 20575 3677
rect 20042 3637 20048 3649
rect 20563 3646 20575 3649
rect 20609 3646 20621 3680
rect 20563 3640 20621 3646
rect 20656 3637 20662 3689
rect 20714 3677 20720 3689
rect 21331 3680 21389 3686
rect 21331 3677 21343 3680
rect 20714 3649 21343 3677
rect 20714 3637 20720 3649
rect 21331 3646 21343 3649
rect 21377 3646 21389 3680
rect 21331 3640 21389 3646
rect 22096 3637 22102 3689
rect 22154 3677 22160 3689
rect 22771 3680 22829 3686
rect 22771 3677 22783 3680
rect 22154 3649 22783 3677
rect 22154 3637 22160 3649
rect 22771 3646 22783 3649
rect 22817 3646 22829 3680
rect 22771 3640 22829 3646
rect 22864 3637 22870 3689
rect 22922 3677 22928 3689
rect 23539 3680 23597 3686
rect 23539 3677 23551 3680
rect 22922 3649 23551 3677
rect 22922 3637 22928 3649
rect 23539 3646 23551 3649
rect 23585 3646 23597 3680
rect 23539 3640 23597 3646
rect 23632 3637 23638 3689
rect 23690 3677 23696 3689
rect 24307 3680 24365 3686
rect 24307 3677 24319 3680
rect 23690 3649 24319 3677
rect 23690 3637 23696 3649
rect 24307 3646 24319 3649
rect 24353 3646 24365 3680
rect 24307 3640 24365 3646
rect 24400 3637 24406 3689
rect 24458 3677 24464 3689
rect 25075 3680 25133 3686
rect 25075 3677 25087 3680
rect 24458 3649 25087 3677
rect 24458 3637 24464 3649
rect 25075 3646 25087 3649
rect 25121 3646 25133 3680
rect 25843 3680 25901 3686
rect 25843 3677 25855 3680
rect 25075 3640 25133 3646
rect 25186 3649 25855 3677
rect 24688 3563 24694 3615
rect 24746 3603 24752 3615
rect 25186 3603 25214 3649
rect 25843 3646 25855 3649
rect 25889 3646 25901 3680
rect 25843 3640 25901 3646
rect 26611 3680 26669 3686
rect 26611 3646 26623 3680
rect 26657 3646 26669 3680
rect 26611 3640 26669 3646
rect 24746 3575 25214 3603
rect 24746 3563 24752 3575
rect 25552 3563 25558 3615
rect 25610 3603 25616 3615
rect 25936 3603 25942 3615
rect 25610 3575 25942 3603
rect 25610 3563 25616 3575
rect 25936 3563 25942 3575
rect 25994 3563 26000 3615
rect 10058 3501 10814 3529
rect 10058 3489 10064 3501
rect 17296 3489 17302 3541
rect 17354 3529 17360 3541
rect 17488 3529 17494 3541
rect 17354 3501 17494 3529
rect 17354 3489 17360 3501
rect 17488 3489 17494 3501
rect 17546 3489 17552 3541
rect 22576 3489 22582 3541
rect 22634 3529 22640 3541
rect 23344 3529 23350 3541
rect 22634 3501 23350 3529
rect 22634 3489 22640 3501
rect 23344 3489 23350 3501
rect 23402 3489 23408 3541
rect 25840 3489 25846 3541
rect 25898 3529 25904 3541
rect 26626 3529 26654 3640
rect 27280 3637 27286 3689
rect 27338 3677 27344 3689
rect 29602 3686 29630 3723
rect 42832 3711 42838 3763
rect 42890 3751 42896 3763
rect 43792 3751 43798 3763
rect 42890 3723 43798 3751
rect 42890 3711 42896 3723
rect 43792 3711 43798 3723
rect 43850 3711 43856 3763
rect 44560 3711 44566 3763
rect 44618 3751 44624 3763
rect 51298 3751 51326 3785
rect 57346 3763 57374 3797
rect 44618 3723 45470 3751
rect 44618 3711 44624 3723
rect 28051 3680 28109 3686
rect 28051 3677 28063 3680
rect 27338 3649 28063 3677
rect 27338 3637 27344 3649
rect 28051 3646 28063 3649
rect 28097 3646 28109 3680
rect 28051 3640 28109 3646
rect 28819 3680 28877 3686
rect 28819 3646 28831 3680
rect 28865 3646 28877 3680
rect 28819 3640 28877 3646
rect 29587 3680 29645 3686
rect 29587 3646 29599 3680
rect 29633 3646 29645 3680
rect 29587 3640 29645 3646
rect 30355 3680 30413 3686
rect 30355 3646 30367 3680
rect 30401 3646 30413 3680
rect 30355 3640 30413 3646
rect 25898 3501 26654 3529
rect 25898 3489 25904 3501
rect 28048 3489 28054 3541
rect 28106 3529 28112 3541
rect 28834 3529 28862 3640
rect 29488 3563 29494 3615
rect 29546 3603 29552 3615
rect 30370 3603 30398 3640
rect 30448 3637 30454 3689
rect 30506 3677 30512 3689
rect 31123 3680 31181 3686
rect 31123 3677 31135 3680
rect 30506 3649 31135 3677
rect 30506 3637 30512 3649
rect 31123 3646 31135 3649
rect 31169 3646 31181 3680
rect 31123 3640 31181 3646
rect 31312 3637 31318 3689
rect 31370 3677 31376 3689
rect 31891 3680 31949 3686
rect 31891 3677 31903 3680
rect 31370 3649 31903 3677
rect 31370 3637 31376 3649
rect 31891 3646 31903 3649
rect 31937 3646 31949 3680
rect 31891 3640 31949 3646
rect 32464 3637 32470 3689
rect 32522 3677 32528 3689
rect 33331 3680 33389 3686
rect 33331 3677 33343 3680
rect 32522 3649 33343 3677
rect 32522 3637 32528 3649
rect 33331 3646 33343 3649
rect 33377 3646 33389 3680
rect 33331 3640 33389 3646
rect 33520 3637 33526 3689
rect 33578 3677 33584 3689
rect 34099 3680 34157 3686
rect 34099 3677 34111 3680
rect 33578 3649 34111 3677
rect 33578 3637 33584 3649
rect 34099 3646 34111 3649
rect 34145 3646 34157 3680
rect 34099 3640 34157 3646
rect 34288 3637 34294 3689
rect 34346 3677 34352 3689
rect 34867 3680 34925 3686
rect 34867 3677 34879 3680
rect 34346 3649 34879 3677
rect 34346 3637 34352 3649
rect 34867 3646 34879 3649
rect 34913 3646 34925 3680
rect 34867 3640 34925 3646
rect 34960 3637 34966 3689
rect 35018 3677 35024 3689
rect 35635 3680 35693 3686
rect 35635 3677 35647 3680
rect 35018 3649 35647 3677
rect 35018 3637 35024 3649
rect 35635 3646 35647 3649
rect 35681 3646 35693 3680
rect 35635 3640 35693 3646
rect 35728 3637 35734 3689
rect 35786 3677 35792 3689
rect 36403 3680 36461 3686
rect 36403 3677 36415 3680
rect 35786 3649 36415 3677
rect 35786 3637 35792 3649
rect 36403 3646 36415 3649
rect 36449 3646 36461 3680
rect 36403 3640 36461 3646
rect 36496 3637 36502 3689
rect 36554 3677 36560 3689
rect 37171 3680 37229 3686
rect 37171 3677 37183 3680
rect 36554 3649 37183 3677
rect 36554 3637 36560 3649
rect 37171 3646 37183 3649
rect 37217 3646 37229 3680
rect 37171 3640 37229 3646
rect 37936 3637 37942 3689
rect 37994 3677 38000 3689
rect 38611 3680 38669 3686
rect 38611 3677 38623 3680
rect 37994 3649 38623 3677
rect 37994 3637 38000 3649
rect 38611 3646 38623 3649
rect 38657 3646 38669 3680
rect 38611 3640 38669 3646
rect 38704 3637 38710 3689
rect 38762 3677 38768 3689
rect 39379 3680 39437 3686
rect 39379 3677 39391 3680
rect 38762 3649 39391 3677
rect 38762 3637 38768 3649
rect 39379 3646 39391 3649
rect 39425 3646 39437 3680
rect 39379 3640 39437 3646
rect 40147 3680 40205 3686
rect 40147 3646 40159 3680
rect 40193 3646 40205 3680
rect 40147 3640 40205 3646
rect 40915 3680 40973 3686
rect 40915 3646 40927 3680
rect 40961 3646 40973 3680
rect 40915 3640 40973 3646
rect 29546 3575 30398 3603
rect 29546 3563 29552 3575
rect 30736 3563 30742 3615
rect 30794 3603 30800 3615
rect 31792 3603 31798 3615
rect 30794 3575 31798 3603
rect 30794 3563 30800 3575
rect 31792 3563 31798 3575
rect 31850 3563 31856 3615
rect 40162 3603 40190 3640
rect 39394 3575 40190 3603
rect 39394 3541 39422 3575
rect 28106 3501 28862 3529
rect 28106 3489 28112 3501
rect 31408 3489 31414 3541
rect 31466 3529 31472 3541
rect 32368 3529 32374 3541
rect 31466 3501 32374 3529
rect 31466 3489 31472 3501
rect 32368 3489 32374 3501
rect 32426 3489 32432 3541
rect 37360 3489 37366 3541
rect 37418 3529 37424 3541
rect 38512 3529 38518 3541
rect 37418 3501 38518 3529
rect 37418 3489 37424 3501
rect 38512 3489 38518 3501
rect 38570 3489 38576 3541
rect 39376 3489 39382 3541
rect 39434 3489 39440 3541
rect 40144 3489 40150 3541
rect 40202 3529 40208 3541
rect 40930 3529 40958 3640
rect 41008 3637 41014 3689
rect 41066 3677 41072 3689
rect 41683 3680 41741 3686
rect 41683 3677 41695 3680
rect 41066 3649 41695 3677
rect 41066 3637 41072 3649
rect 41683 3646 41695 3649
rect 41729 3646 41741 3680
rect 41683 3640 41741 3646
rect 42451 3680 42509 3686
rect 42451 3646 42463 3680
rect 42497 3646 42509 3680
rect 42451 3640 42509 3646
rect 40202 3501 40958 3529
rect 40202 3489 40208 3501
rect 41584 3489 41590 3541
rect 41642 3529 41648 3541
rect 42466 3529 42494 3640
rect 42736 3637 42742 3689
rect 42794 3677 42800 3689
rect 45442 3686 45470 3723
rect 49378 3723 51326 3751
rect 43891 3680 43949 3686
rect 43891 3677 43903 3680
rect 42794 3649 43903 3677
rect 42794 3637 42800 3649
rect 43891 3646 43903 3649
rect 43937 3646 43949 3680
rect 43891 3640 43949 3646
rect 44659 3680 44717 3686
rect 44659 3646 44671 3680
rect 44705 3646 44717 3680
rect 44659 3640 44717 3646
rect 45427 3680 45485 3686
rect 45427 3646 45439 3680
rect 45473 3646 45485 3680
rect 45427 3640 45485 3646
rect 46195 3680 46253 3686
rect 46195 3646 46207 3680
rect 46241 3646 46253 3680
rect 46195 3640 46253 3646
rect 46963 3680 47021 3686
rect 46963 3646 46975 3680
rect 47009 3646 47021 3680
rect 46963 3640 47021 3646
rect 43792 3563 43798 3615
rect 43850 3603 43856 3615
rect 44674 3603 44702 3640
rect 43850 3575 44702 3603
rect 43850 3563 43856 3575
rect 45232 3563 45238 3615
rect 45290 3603 45296 3615
rect 46210 3603 46238 3640
rect 45290 3575 46238 3603
rect 45290 3563 45296 3575
rect 41642 3501 42494 3529
rect 41642 3489 41648 3501
rect 46000 3489 46006 3541
rect 46058 3529 46064 3541
rect 46978 3529 47006 3640
rect 47152 3637 47158 3689
rect 47210 3677 47216 3689
rect 47731 3680 47789 3686
rect 47731 3677 47743 3680
rect 47210 3649 47743 3677
rect 47210 3637 47216 3649
rect 47731 3646 47743 3649
rect 47777 3646 47789 3680
rect 47731 3640 47789 3646
rect 48208 3637 48214 3689
rect 48266 3677 48272 3689
rect 49171 3680 49229 3686
rect 49171 3677 49183 3680
rect 48266 3649 49183 3677
rect 48266 3637 48272 3649
rect 49171 3646 49183 3649
rect 49217 3646 49229 3680
rect 49171 3640 49229 3646
rect 46058 3501 47006 3529
rect 46058 3489 46064 3501
rect 47536 3489 47542 3541
rect 47594 3529 47600 3541
rect 48304 3529 48310 3541
rect 47594 3501 48310 3529
rect 47594 3489 47600 3501
rect 48304 3489 48310 3501
rect 48362 3489 48368 3541
rect 3434 3427 4670 3455
rect 12115 3458 12173 3464
rect 3434 3415 3440 3427
rect 12115 3424 12127 3458
rect 12161 3455 12173 3458
rect 12403 3458 12461 3464
rect 12403 3455 12415 3458
rect 12161 3427 12415 3455
rect 12161 3424 12173 3427
rect 12115 3418 12173 3424
rect 12403 3424 12415 3427
rect 12449 3455 12461 3458
rect 49378 3455 49406 3723
rect 55888 3711 55894 3763
rect 55946 3751 55952 3763
rect 55946 3723 56798 3751
rect 55946 3711 55952 3723
rect 50515 3680 50573 3686
rect 50515 3646 50527 3680
rect 50561 3677 50573 3680
rect 50704 3677 50710 3689
rect 50561 3649 50710 3677
rect 50561 3646 50573 3649
rect 50515 3640 50573 3646
rect 50704 3637 50710 3649
rect 50762 3637 50768 3689
rect 50800 3637 50806 3689
rect 50858 3677 50864 3689
rect 51187 3680 51245 3686
rect 51187 3677 51199 3680
rect 50858 3649 51199 3677
rect 50858 3637 50864 3649
rect 51187 3646 51199 3649
rect 51233 3646 51245 3680
rect 51187 3640 51245 3646
rect 51280 3637 51286 3689
rect 51338 3677 51344 3689
rect 51955 3680 52013 3686
rect 51955 3677 51967 3680
rect 51338 3649 51967 3677
rect 51338 3637 51344 3649
rect 51955 3646 51967 3649
rect 52001 3646 52013 3680
rect 51955 3640 52013 3646
rect 52048 3637 52054 3689
rect 52106 3677 52112 3689
rect 52723 3680 52781 3686
rect 52723 3677 52735 3680
rect 52106 3649 52735 3677
rect 52106 3637 52112 3649
rect 52723 3646 52735 3649
rect 52769 3646 52781 3680
rect 52723 3640 52781 3646
rect 53392 3637 53398 3689
rect 53450 3677 53456 3689
rect 56770 3686 56798 3723
rect 57328 3711 57334 3763
rect 57386 3711 57392 3763
rect 54451 3680 54509 3686
rect 54451 3677 54463 3680
rect 53450 3649 54463 3677
rect 53450 3637 53456 3649
rect 54451 3646 54463 3649
rect 54497 3646 54509 3680
rect 54451 3640 54509 3646
rect 55219 3680 55277 3686
rect 55219 3646 55231 3680
rect 55265 3646 55277 3680
rect 55219 3640 55277 3646
rect 55987 3680 56045 3686
rect 55987 3646 55999 3680
rect 56033 3646 56045 3680
rect 55987 3640 56045 3646
rect 56755 3680 56813 3686
rect 56755 3646 56767 3680
rect 56801 3646 56813 3680
rect 56755 3640 56813 3646
rect 57523 3680 57581 3686
rect 57523 3646 57535 3680
rect 57569 3646 57581 3680
rect 57523 3640 57581 3646
rect 54448 3489 54454 3541
rect 54506 3529 54512 3541
rect 55234 3529 55262 3640
rect 54506 3501 55262 3529
rect 54506 3489 54512 3501
rect 12449 3427 49406 3455
rect 12449 3424 12461 3427
rect 12403 3418 12461 3424
rect 55216 3415 55222 3467
rect 55274 3455 55280 3467
rect 56002 3455 56030 3640
rect 56272 3563 56278 3615
rect 56330 3603 56336 3615
rect 57538 3603 57566 3640
rect 56330 3575 57566 3603
rect 56330 3563 56336 3575
rect 56368 3489 56374 3541
rect 56426 3529 56432 3541
rect 57136 3529 57142 3541
rect 56426 3501 57142 3529
rect 56426 3489 56432 3501
rect 57136 3489 57142 3501
rect 57194 3489 57200 3541
rect 55274 3427 56030 3455
rect 55274 3415 55280 3427
rect 1152 3356 58848 3378
rect 1152 3304 19654 3356
rect 19706 3304 19718 3356
rect 19770 3304 19782 3356
rect 19834 3304 19846 3356
rect 19898 3304 50374 3356
rect 50426 3304 50438 3356
rect 50490 3304 50502 3356
rect 50554 3304 50566 3356
rect 50618 3304 58848 3356
rect 1152 3282 58848 3304
rect 1456 3193 1462 3245
rect 1514 3233 1520 3245
rect 2128 3233 2134 3245
rect 1514 3205 2134 3233
rect 1514 3193 1520 3205
rect 2128 3193 2134 3205
rect 2186 3193 2192 3245
rect 12016 3193 12022 3245
rect 12074 3233 12080 3245
rect 13360 3233 13366 3245
rect 12074 3205 13366 3233
rect 12074 3193 12080 3205
rect 13360 3193 13366 3205
rect 13418 3193 13424 3245
rect 17488 3193 17494 3245
rect 17546 3233 17552 3245
rect 18352 3233 18358 3245
rect 17546 3205 18358 3233
rect 17546 3193 17552 3205
rect 18352 3193 18358 3205
rect 18410 3193 18416 3245
rect 19696 3193 19702 3245
rect 19754 3233 19760 3245
rect 20368 3233 20374 3245
rect 19754 3205 20374 3233
rect 19754 3193 19760 3205
rect 20368 3193 20374 3205
rect 20426 3193 20432 3245
rect 23344 3193 23350 3245
rect 23402 3233 23408 3245
rect 24208 3233 24214 3245
rect 23402 3205 24214 3233
rect 23402 3193 23408 3205
rect 24208 3193 24214 3205
rect 24266 3193 24272 3245
rect 25936 3193 25942 3245
rect 25994 3233 26000 3245
rect 26896 3233 26902 3245
rect 25994 3205 26902 3233
rect 25994 3193 26000 3205
rect 26896 3193 26902 3205
rect 26954 3193 26960 3245
rect 27376 3193 27382 3245
rect 27434 3233 27440 3245
rect 28432 3233 28438 3245
rect 27434 3205 28438 3233
rect 27434 3193 27440 3205
rect 28432 3193 28438 3205
rect 28490 3193 28496 3245
rect 28528 3193 28534 3245
rect 28586 3233 28592 3245
rect 29392 3233 29398 3245
rect 28586 3205 29398 3233
rect 28586 3193 28592 3205
rect 29392 3193 29398 3205
rect 29450 3193 29456 3245
rect 30448 3193 30454 3245
rect 30506 3233 30512 3245
rect 31888 3233 31894 3245
rect 30506 3205 31894 3233
rect 30506 3193 30512 3205
rect 31888 3193 31894 3205
rect 31946 3193 31952 3245
rect 32656 3193 32662 3245
rect 32714 3233 32720 3245
rect 34096 3233 34102 3245
rect 32714 3205 34102 3233
rect 32714 3193 32720 3205
rect 34096 3193 34102 3205
rect 34154 3193 34160 3245
rect 38512 3193 38518 3245
rect 38570 3233 38576 3245
rect 39568 3233 39574 3245
rect 38570 3205 39574 3233
rect 38570 3193 38576 3205
rect 39568 3193 39574 3205
rect 39626 3193 39632 3245
rect 41200 3193 41206 3245
rect 41258 3233 41264 3245
rect 41680 3233 41686 3245
rect 41258 3205 41686 3233
rect 41258 3193 41264 3205
rect 41680 3193 41686 3205
rect 41738 3193 41744 3245
rect 44080 3193 44086 3245
rect 44138 3233 44144 3245
rect 45424 3233 45430 3245
rect 44138 3205 45430 3233
rect 44138 3193 44144 3205
rect 45424 3193 45430 3205
rect 45482 3193 45488 3245
rect 48496 3193 48502 3245
rect 48554 3233 48560 3245
rect 49648 3233 49654 3245
rect 48554 3205 49654 3233
rect 48554 3193 48560 3205
rect 49648 3193 49654 3205
rect 49706 3193 49712 3245
rect 52048 3193 52054 3245
rect 52106 3233 52112 3245
rect 52432 3233 52438 3245
rect 52106 3205 52438 3233
rect 52106 3193 52112 3205
rect 52432 3193 52438 3205
rect 52490 3193 52496 3245
rect 56848 3193 56854 3245
rect 56906 3233 56912 3245
rect 58288 3233 58294 3245
rect 56906 3205 58294 3233
rect 56906 3193 56912 3205
rect 58288 3193 58294 3205
rect 58346 3193 58352 3245
rect 208 3119 214 3171
rect 266 3159 272 3171
rect 1744 3159 1750 3171
rect 266 3131 1750 3159
rect 266 3119 272 3131
rect 1744 3119 1750 3131
rect 1802 3119 1808 3171
rect 12208 3119 12214 3171
rect 12266 3159 12272 3171
rect 12976 3159 12982 3171
rect 12266 3131 12982 3159
rect 12266 3119 12272 3131
rect 12976 3119 12982 3131
rect 13034 3119 13040 3171
rect 20080 3119 20086 3171
rect 20138 3159 20144 3171
rect 21424 3159 21430 3171
rect 20138 3131 21430 3159
rect 20138 3119 20144 3131
rect 21424 3119 21430 3131
rect 21482 3119 21488 3171
rect 22960 3119 22966 3171
rect 23018 3159 23024 3171
rect 23920 3159 23926 3171
rect 23018 3131 23926 3159
rect 23018 3119 23024 3131
rect 23920 3119 23926 3131
rect 23978 3119 23984 3171
rect 24976 3119 24982 3171
rect 25034 3159 25040 3171
rect 26608 3159 26614 3171
rect 25034 3131 26614 3159
rect 25034 3119 25040 3131
rect 26608 3119 26614 3131
rect 26666 3119 26672 3171
rect 28240 3119 28246 3171
rect 28298 3159 28304 3171
rect 29296 3159 29302 3171
rect 28298 3131 29302 3159
rect 28298 3119 28304 3131
rect 29296 3119 29302 3131
rect 29354 3119 29360 3171
rect 29776 3119 29782 3171
rect 29834 3159 29840 3171
rect 30544 3159 30550 3171
rect 29834 3131 30550 3159
rect 29834 3119 29840 3131
rect 30544 3119 30550 3131
rect 30602 3119 30608 3171
rect 31792 3119 31798 3171
rect 31850 3159 31856 3171
rect 31984 3159 31990 3171
rect 31850 3131 31990 3159
rect 31850 3119 31856 3131
rect 31984 3119 31990 3131
rect 32042 3119 32048 3171
rect 32560 3119 32566 3171
rect 32618 3159 32624 3171
rect 33712 3159 33718 3171
rect 32618 3131 33718 3159
rect 32618 3119 32624 3131
rect 33712 3119 33718 3131
rect 33770 3119 33776 3171
rect 35347 3162 35405 3168
rect 35347 3128 35359 3162
rect 35393 3159 35405 3162
rect 35536 3159 35542 3171
rect 35393 3131 35542 3159
rect 35393 3128 35405 3131
rect 35347 3122 35405 3128
rect 35536 3119 35542 3131
rect 35594 3159 35600 3171
rect 35594 3131 35678 3159
rect 35594 3119 35600 3131
rect 8944 3045 8950 3097
rect 9002 3085 9008 3097
rect 13267 3088 13325 3094
rect 13267 3085 13279 3088
rect 9002 3057 13279 3085
rect 9002 3045 9008 3057
rect 13267 3054 13279 3057
rect 13313 3054 13325 3088
rect 13267 3048 13325 3054
rect 18352 3045 18358 3097
rect 18410 3085 18416 3097
rect 19024 3085 19030 3097
rect 18410 3057 19030 3085
rect 18410 3045 18416 3057
rect 19024 3045 19030 3057
rect 19082 3045 19088 3097
rect 19792 3045 19798 3097
rect 19850 3085 19856 3097
rect 20176 3085 20182 3097
rect 19850 3057 20182 3085
rect 19850 3045 19856 3057
rect 20176 3045 20182 3057
rect 20234 3045 20240 3097
rect 22384 3045 22390 3097
rect 22442 3085 22448 3097
rect 23536 3085 23542 3097
rect 22442 3057 23542 3085
rect 22442 3045 22448 3057
rect 23536 3045 23542 3057
rect 23594 3045 23600 3097
rect 23824 3045 23830 3097
rect 23882 3085 23888 3097
rect 25072 3085 25078 3097
rect 23882 3057 25078 3085
rect 23882 3045 23888 3057
rect 25072 3045 25078 3057
rect 25130 3045 25136 3097
rect 25360 3045 25366 3097
rect 25418 3085 25424 3097
rect 26224 3085 26230 3097
rect 25418 3057 26230 3085
rect 25418 3045 25424 3057
rect 26224 3045 26230 3057
rect 26282 3045 26288 3097
rect 27472 3045 27478 3097
rect 27530 3085 27536 3097
rect 28912 3085 28918 3097
rect 27530 3057 28918 3085
rect 27530 3045 27536 3057
rect 28912 3045 28918 3057
rect 28970 3045 28976 3097
rect 29392 3045 29398 3097
rect 29450 3085 29456 3097
rect 31120 3085 31126 3097
rect 29450 3057 31126 3085
rect 29450 3045 29456 3057
rect 31120 3045 31126 3057
rect 31178 3045 31184 3097
rect 31888 3045 31894 3097
rect 31946 3085 31952 3097
rect 33328 3085 33334 3097
rect 31946 3057 33334 3085
rect 31946 3045 31952 3057
rect 33328 3045 33334 3057
rect 33386 3045 33392 3097
rect 34000 3045 34006 3097
rect 34058 3085 34064 3097
rect 34480 3085 34486 3097
rect 34058 3057 34486 3085
rect 34058 3045 34064 3057
rect 34480 3045 34486 3057
rect 34538 3045 34544 3097
rect 35650 3094 35678 3131
rect 37072 3119 37078 3171
rect 37130 3159 37136 3171
rect 38608 3159 38614 3171
rect 37130 3131 38614 3159
rect 37130 3119 37136 3131
rect 38608 3119 38614 3131
rect 38666 3119 38672 3171
rect 39664 3119 39670 3171
rect 39722 3159 39728 3171
rect 40912 3159 40918 3171
rect 39722 3131 40918 3159
rect 39722 3119 39728 3131
rect 40912 3119 40918 3131
rect 40970 3119 40976 3171
rect 41104 3119 41110 3171
rect 41162 3159 41168 3171
rect 42160 3159 42166 3171
rect 41162 3131 42166 3159
rect 41162 3119 41168 3131
rect 42160 3119 42166 3131
rect 42218 3119 42224 3171
rect 44848 3159 44854 3171
rect 43234 3131 44854 3159
rect 43234 3097 43262 3131
rect 44848 3119 44854 3131
rect 44906 3119 44912 3171
rect 45136 3119 45142 3171
rect 45194 3159 45200 3171
rect 46288 3159 46294 3171
rect 45194 3131 46294 3159
rect 45194 3119 45200 3131
rect 46288 3119 46294 3131
rect 46346 3119 46352 3171
rect 48112 3119 48118 3171
rect 48170 3159 48176 3171
rect 48976 3159 48982 3171
rect 48170 3131 48982 3159
rect 48170 3119 48176 3131
rect 48976 3119 48982 3131
rect 49034 3119 49040 3171
rect 57328 3119 57334 3171
rect 57386 3159 57392 3171
rect 58000 3159 58006 3171
rect 57386 3131 58006 3159
rect 57386 3119 57392 3131
rect 58000 3119 58006 3131
rect 58058 3119 58064 3171
rect 35635 3088 35693 3094
rect 35635 3054 35647 3088
rect 35681 3054 35693 3088
rect 35635 3048 35693 3054
rect 35920 3045 35926 3097
rect 35978 3085 35984 3097
rect 36112 3085 36118 3097
rect 35978 3057 36118 3085
rect 35978 3045 35984 3057
rect 36112 3045 36118 3057
rect 36170 3045 36176 3097
rect 36688 3045 36694 3097
rect 36746 3085 36752 3097
rect 37552 3085 37558 3097
rect 36746 3057 37558 3085
rect 36746 3045 36752 3057
rect 37552 3045 37558 3057
rect 37610 3045 37616 3097
rect 38320 3045 38326 3097
rect 38378 3085 38384 3097
rect 38378 3057 40094 3085
rect 38378 3045 38384 3057
rect 16 2971 22 3023
rect 74 3011 80 3023
rect 1555 3014 1613 3020
rect 1555 3011 1567 3014
rect 74 2983 1567 3011
rect 74 2971 80 2983
rect 1555 2980 1567 2983
rect 1601 2980 1613 3014
rect 2323 3014 2381 3020
rect 2323 3011 2335 3014
rect 1555 2974 1613 2980
rect 1666 2983 2335 3011
rect 688 2897 694 2949
rect 746 2937 752 2949
rect 1666 2937 1694 2983
rect 2323 2980 2335 2983
rect 2369 2980 2381 3014
rect 3091 3014 3149 3020
rect 3091 3011 3103 3014
rect 2323 2974 2381 2980
rect 2866 2983 3103 3011
rect 746 2909 1694 2937
rect 746 2897 752 2909
rect 2128 2897 2134 2949
rect 2186 2937 2192 2949
rect 2866 2937 2894 2983
rect 3091 2980 3103 2983
rect 3137 2980 3149 3014
rect 4912 3011 4918 3023
rect 4873 2983 4918 3011
rect 3091 2974 3149 2980
rect 4912 2971 4918 2983
rect 4970 2971 4976 3023
rect 5200 2971 5206 3023
rect 5258 3011 5264 3023
rect 5683 3014 5741 3020
rect 5683 3011 5695 3014
rect 5258 2983 5695 3011
rect 5258 2971 5264 2983
rect 5683 2980 5695 2983
rect 5729 2980 5741 3014
rect 5683 2974 5741 2980
rect 5968 2971 5974 3023
rect 6026 3011 6032 3023
rect 7027 3014 7085 3020
rect 7027 3011 7039 3014
rect 6026 2983 7039 3011
rect 6026 2971 6032 2983
rect 7027 2980 7039 2983
rect 7073 2980 7085 3014
rect 7027 2974 7085 2980
rect 7795 3014 7853 3020
rect 7795 2980 7807 3014
rect 7841 2980 7853 3014
rect 7795 2974 7853 2980
rect 2186 2909 2894 2937
rect 2186 2897 2192 2909
rect 6736 2897 6742 2949
rect 6794 2937 6800 2949
rect 7810 2937 7838 2974
rect 8176 2971 8182 3023
rect 8234 3011 8240 3023
rect 9715 3014 9773 3020
rect 9715 3011 9727 3014
rect 8234 2983 9727 3011
rect 8234 2971 8240 2983
rect 9715 2980 9727 2983
rect 9761 2980 9773 3014
rect 9715 2974 9773 2980
rect 10483 3014 10541 3020
rect 10483 2980 10495 3014
rect 10529 2980 10541 3014
rect 12976 3011 12982 3023
rect 12937 2983 12982 3011
rect 10483 2974 10541 2980
rect 6794 2909 7838 2937
rect 6794 2897 6800 2909
rect 8944 2897 8950 2949
rect 9002 2937 9008 2949
rect 10498 2937 10526 2974
rect 12976 2971 12982 2983
rect 13034 2971 13040 3023
rect 13360 2971 13366 3023
rect 13418 3011 13424 3023
rect 13747 3014 13805 3020
rect 13747 3011 13759 3014
rect 13418 2983 13759 3011
rect 13418 2971 13424 2983
rect 13747 2980 13759 2983
rect 13793 2980 13805 3014
rect 13747 2974 13805 2980
rect 14512 2971 14518 3023
rect 14570 3011 14576 3023
rect 15091 3014 15149 3020
rect 15091 3011 15103 3014
rect 14570 2983 15103 3011
rect 14570 2971 14576 2983
rect 15091 2980 15103 2983
rect 15137 2980 15149 3014
rect 16624 3011 16630 3023
rect 16585 2983 16630 3011
rect 15091 2974 15149 2980
rect 16624 2971 16630 2983
rect 16682 2971 16688 3023
rect 17008 2971 17014 3023
rect 17066 3011 17072 3023
rect 17779 3014 17837 3020
rect 17779 3011 17791 3014
rect 17066 2983 17791 3011
rect 17066 2971 17072 2983
rect 17779 2980 17791 2983
rect 17825 2980 17837 3014
rect 17779 2974 17837 2980
rect 18547 3014 18605 3020
rect 18547 2980 18559 3014
rect 18593 2980 18605 3014
rect 18547 2974 18605 2980
rect 9002 2909 10526 2937
rect 9002 2897 9008 2909
rect 15376 2897 15382 2949
rect 15434 2937 15440 2949
rect 16528 2937 16534 2949
rect 15434 2909 16534 2937
rect 15434 2897 15440 2909
rect 16528 2897 16534 2909
rect 16586 2897 16592 2949
rect 17680 2897 17686 2949
rect 17738 2937 17744 2949
rect 18562 2937 18590 2974
rect 18832 2971 18838 3023
rect 18890 3011 18896 3023
rect 20467 3014 20525 3020
rect 20467 3011 20479 3014
rect 18890 2983 20479 3011
rect 18890 2971 18896 2983
rect 20467 2980 20479 2983
rect 20513 2980 20525 3014
rect 21235 3014 21293 3020
rect 21235 3011 21247 3014
rect 20467 2974 20525 2980
rect 20578 2983 21247 3011
rect 17738 2909 18590 2937
rect 17738 2897 17744 2909
rect 19600 2897 19606 2949
rect 19658 2937 19664 2949
rect 20578 2937 20606 2983
rect 21235 2980 21247 2983
rect 21281 2980 21293 3014
rect 21235 2974 21293 2980
rect 21424 2971 21430 3023
rect 21482 3011 21488 3023
rect 23155 3014 23213 3020
rect 23155 3011 23167 3014
rect 21482 2983 23167 3011
rect 21482 2971 21488 2983
rect 23155 2980 23167 2983
rect 23201 2980 23213 3014
rect 23155 2974 23213 2980
rect 23923 3014 23981 3020
rect 23923 2980 23935 3014
rect 23969 2980 23981 3014
rect 23923 2974 23981 2980
rect 19658 2909 20606 2937
rect 19658 2897 19664 2909
rect 20944 2897 20950 2949
rect 21002 2937 21008 2949
rect 21712 2937 21718 2949
rect 21002 2909 21718 2937
rect 21002 2897 21008 2909
rect 21712 2897 21718 2909
rect 21770 2897 21776 2949
rect 22480 2897 22486 2949
rect 22538 2937 22544 2949
rect 23938 2937 23966 2974
rect 24016 2971 24022 3023
rect 24074 3011 24080 3023
rect 25843 3014 25901 3020
rect 25843 3011 25855 3014
rect 24074 2983 25855 3011
rect 24074 2971 24080 2983
rect 25843 2980 25855 2983
rect 25889 2980 25901 3014
rect 25843 2974 25901 2980
rect 26611 3014 26669 3020
rect 26611 2980 26623 3014
rect 26657 2980 26669 3014
rect 26611 2974 26669 2980
rect 22538 2909 23966 2937
rect 22538 2897 22544 2909
rect 24208 2897 24214 2949
rect 24266 2937 24272 2949
rect 24880 2937 24886 2949
rect 24266 2909 24886 2937
rect 24266 2897 24272 2909
rect 24880 2897 24886 2909
rect 24938 2897 24944 2949
rect 25072 2897 25078 2949
rect 25130 2937 25136 2949
rect 26626 2937 26654 2974
rect 26896 2971 26902 3023
rect 26954 3011 26960 3023
rect 28531 3014 28589 3020
rect 28531 3011 28543 3014
rect 26954 2983 28543 3011
rect 26954 2971 26960 2983
rect 28531 2980 28543 2983
rect 28577 2980 28589 3014
rect 28531 2974 28589 2980
rect 29299 3014 29357 3020
rect 29299 2980 29311 3014
rect 29345 2980 29357 3014
rect 29299 2974 29357 2980
rect 25130 2909 26654 2937
rect 25130 2897 25136 2909
rect 27664 2897 27670 2949
rect 27722 2937 27728 2949
rect 29314 2937 29342 2974
rect 29872 2971 29878 3023
rect 29930 3011 29936 3023
rect 31219 3014 31277 3020
rect 31219 3011 31231 3014
rect 29930 2983 31231 3011
rect 29930 2971 29936 2983
rect 31219 2980 31231 2983
rect 31265 2980 31277 3014
rect 31219 2974 31277 2980
rect 31987 3014 32045 3020
rect 31987 2980 31999 3014
rect 32033 2980 32045 3014
rect 31987 2974 32045 2980
rect 27722 2909 29342 2937
rect 27722 2897 27728 2909
rect 30544 2897 30550 2949
rect 30602 2937 30608 2949
rect 32002 2937 32030 2974
rect 32080 2971 32086 3023
rect 32138 3011 32144 3023
rect 33907 3014 33965 3020
rect 33907 3011 33919 3014
rect 32138 2983 33919 3011
rect 32138 2971 32144 2983
rect 33907 2980 33919 2983
rect 33953 2980 33965 3014
rect 33907 2974 33965 2980
rect 34675 3014 34733 3020
rect 34675 2980 34687 3014
rect 34721 2980 34733 3014
rect 34675 2974 34733 2980
rect 30602 2909 32030 2937
rect 30602 2897 30608 2909
rect 32272 2897 32278 2949
rect 32330 2937 32336 2949
rect 33136 2937 33142 2949
rect 32330 2909 33142 2937
rect 32330 2897 32336 2909
rect 33136 2897 33142 2909
rect 33194 2897 33200 2949
rect 33328 2897 33334 2949
rect 33386 2937 33392 2949
rect 34690 2937 34718 2974
rect 35344 2971 35350 3023
rect 35402 3011 35408 3023
rect 36595 3014 36653 3020
rect 36595 3011 36607 3014
rect 35402 2983 36607 3011
rect 35402 2971 35408 2983
rect 36595 2980 36607 2983
rect 36641 2980 36653 3014
rect 36595 2974 36653 2980
rect 37264 2971 37270 3023
rect 37322 3011 37328 3023
rect 40066 3020 40094 3057
rect 40816 3045 40822 3097
rect 40874 3085 40880 3097
rect 41011 3088 41069 3094
rect 41011 3085 41023 3088
rect 40874 3057 41023 3085
rect 40874 3045 40880 3057
rect 41011 3054 41023 3057
rect 41057 3054 41069 3088
rect 41011 3048 41069 3054
rect 41200 3045 41206 3097
rect 41258 3085 41264 3097
rect 41258 3057 42782 3085
rect 41258 3045 41264 3057
rect 37363 3014 37421 3020
rect 37363 3011 37375 3014
rect 37322 2983 37375 3011
rect 37322 2971 37328 2983
rect 37363 2980 37375 2983
rect 37409 2980 37421 3014
rect 39283 3014 39341 3020
rect 39283 3011 39295 3014
rect 37363 2974 37421 2980
rect 37570 2983 39295 3011
rect 37570 2949 37598 2983
rect 39283 2980 39295 2983
rect 39329 2980 39341 3014
rect 39283 2974 39341 2980
rect 40051 3014 40109 3020
rect 40051 2980 40063 3014
rect 40097 2980 40109 3014
rect 40051 2974 40109 2980
rect 40528 2971 40534 3023
rect 40586 3011 40592 3023
rect 41971 3014 42029 3020
rect 41971 3011 41983 3014
rect 40586 2983 41983 3011
rect 40586 2971 40592 2983
rect 41971 2980 41983 2983
rect 42017 2980 42029 3014
rect 41971 2974 42029 2980
rect 42160 2971 42166 3023
rect 42218 3011 42224 3023
rect 42640 3011 42646 3023
rect 42218 2983 42646 3011
rect 42218 2971 42224 2983
rect 42640 2971 42646 2983
rect 42698 2971 42704 3023
rect 42754 3020 42782 3057
rect 43216 3045 43222 3097
rect 43274 3045 43280 3097
rect 44752 3045 44758 3097
rect 44810 3085 44816 3097
rect 46192 3085 46198 3097
rect 44810 3057 46198 3085
rect 44810 3045 44816 3057
rect 46192 3045 46198 3057
rect 46250 3045 46256 3097
rect 46384 3045 46390 3097
rect 46442 3085 46448 3097
rect 46442 3057 47534 3085
rect 46442 3045 46448 3057
rect 42739 3014 42797 3020
rect 42739 2980 42751 3014
rect 42785 2980 42797 3014
rect 42739 2974 42797 2980
rect 43024 2971 43030 3023
rect 43082 3011 43088 3023
rect 44659 3014 44717 3020
rect 44659 3011 44671 3014
rect 43082 2983 44671 3011
rect 43082 2971 43088 2983
rect 44659 2980 44671 2983
rect 44705 2980 44717 3014
rect 44659 2974 44717 2980
rect 45427 3014 45485 3020
rect 45427 2980 45439 3014
rect 45473 2980 45485 3014
rect 45427 2974 45485 2980
rect 33386 2909 34718 2937
rect 33386 2897 33392 2909
rect 35440 2897 35446 2949
rect 35498 2937 35504 2949
rect 36016 2937 36022 2949
rect 35498 2909 36022 2937
rect 35498 2897 35504 2909
rect 36016 2897 36022 2909
rect 36074 2897 36080 2949
rect 37552 2897 37558 2949
rect 37610 2897 37616 2949
rect 38128 2897 38134 2949
rect 38186 2937 38192 2949
rect 39088 2937 39094 2949
rect 38186 2909 39094 2937
rect 38186 2897 38192 2909
rect 39088 2897 39094 2909
rect 39146 2897 39152 2949
rect 39184 2897 39190 2949
rect 39242 2937 39248 2949
rect 39952 2937 39958 2949
rect 39242 2909 39958 2937
rect 39242 2897 39248 2909
rect 39952 2897 39958 2909
rect 40010 2897 40016 2949
rect 40834 2909 41246 2937
rect 40834 2875 40862 2909
rect 2608 2823 2614 2875
rect 2666 2863 2672 2875
rect 2666 2835 13406 2863
rect 2666 2823 2672 2835
rect 5104 2749 5110 2801
rect 5162 2789 5168 2801
rect 5776 2789 5782 2801
rect 5162 2761 5782 2789
rect 5162 2749 5168 2761
rect 5776 2749 5782 2761
rect 5834 2749 5840 2801
rect 8752 2789 8758 2801
rect 8713 2761 8758 2789
rect 8752 2749 8758 2761
rect 8810 2749 8816 2801
rect 13378 2789 13406 2835
rect 14224 2823 14230 2875
rect 14282 2863 14288 2875
rect 14282 2835 34622 2863
rect 14282 2823 14288 2835
rect 33808 2789 33814 2801
rect 13378 2761 33814 2789
rect 33808 2749 33814 2761
rect 33866 2749 33872 2801
rect 34594 2789 34622 2835
rect 40816 2823 40822 2875
rect 40874 2823 40880 2875
rect 41218 2863 41246 2909
rect 41488 2897 41494 2949
rect 41546 2937 41552 2949
rect 42064 2937 42070 2949
rect 41546 2909 42070 2937
rect 41546 2897 41552 2909
rect 42064 2897 42070 2909
rect 42122 2897 42128 2949
rect 42544 2897 42550 2949
rect 42602 2937 42608 2949
rect 43312 2937 43318 2949
rect 42602 2909 43318 2937
rect 42602 2897 42608 2909
rect 43312 2897 43318 2909
rect 43370 2897 43376 2949
rect 44176 2897 44182 2949
rect 44234 2937 44240 2949
rect 45442 2937 45470 2974
rect 45616 2971 45622 3023
rect 45674 3011 45680 3023
rect 47347 3014 47405 3020
rect 47347 3011 47359 3014
rect 45674 2983 47359 3011
rect 45674 2971 45680 2983
rect 47347 2980 47359 2983
rect 47393 2980 47405 3014
rect 47506 3011 47534 3057
rect 51760 3045 51766 3097
rect 51818 3085 51824 3097
rect 52240 3085 52246 3097
rect 51818 3057 52246 3085
rect 51818 3045 51824 3057
rect 52240 3045 52246 3057
rect 52298 3045 52304 3097
rect 53107 3088 53165 3094
rect 53107 3054 53119 3088
rect 53153 3085 53165 3088
rect 53200 3085 53206 3097
rect 53153 3057 53206 3085
rect 53153 3054 53165 3057
rect 53107 3048 53165 3054
rect 53200 3045 53206 3057
rect 53258 3045 53264 3097
rect 48115 3014 48173 3020
rect 48115 3011 48127 3014
rect 47506 2983 48127 3011
rect 47347 2974 47405 2980
rect 48115 2980 48127 2983
rect 48161 2980 48173 3014
rect 48115 2974 48173 2980
rect 49648 2971 49654 3023
rect 49706 3011 49712 3023
rect 50035 3014 50093 3020
rect 50035 3011 50047 3014
rect 49706 2983 50047 3011
rect 49706 2971 49712 2983
rect 50035 2980 50047 2983
rect 50081 2980 50093 3014
rect 50035 2974 50093 2980
rect 50803 3014 50861 3020
rect 50803 2980 50815 3014
rect 50849 2980 50861 3014
rect 50803 2974 50861 2980
rect 44234 2909 45470 2937
rect 44234 2897 44240 2909
rect 46288 2897 46294 2949
rect 46346 2937 46352 2949
rect 47632 2937 47638 2949
rect 46346 2909 47638 2937
rect 46346 2897 46352 2909
rect 47632 2897 47638 2909
rect 47690 2897 47696 2949
rect 48976 2897 48982 2949
rect 49034 2937 49040 2949
rect 49840 2937 49846 2949
rect 49034 2909 49846 2937
rect 49034 2897 49040 2909
rect 49840 2897 49846 2909
rect 49898 2897 49904 2949
rect 50818 2937 50846 2974
rect 51472 2971 51478 3023
rect 51530 3011 51536 3023
rect 52723 3014 52781 3020
rect 52723 3011 52735 3014
rect 51530 2983 52735 3011
rect 51530 2971 51536 2983
rect 52723 2980 52735 2983
rect 52769 2980 52781 3014
rect 53491 3014 53549 3020
rect 53491 3011 53503 3014
rect 52723 2974 52781 2980
rect 52834 2983 53503 3011
rect 50050 2909 50846 2937
rect 50050 2875 50078 2909
rect 51376 2897 51382 2949
rect 51434 2937 51440 2949
rect 51856 2937 51862 2949
rect 51434 2909 51862 2937
rect 51434 2897 51440 2909
rect 51856 2897 51862 2909
rect 51914 2897 51920 2949
rect 52240 2897 52246 2949
rect 52298 2937 52304 2949
rect 52834 2937 52862 2983
rect 53491 2980 53503 2983
rect 53537 2980 53549 3014
rect 53491 2974 53549 2980
rect 53776 2971 53782 3023
rect 53834 3011 53840 3023
rect 55411 3014 55469 3020
rect 55411 3011 55423 3014
rect 53834 2983 55423 3011
rect 53834 2971 53840 2983
rect 55411 2980 55423 2983
rect 55457 2980 55469 3014
rect 55411 2974 55469 2980
rect 56179 3014 56237 3020
rect 56179 2980 56191 3014
rect 56225 2980 56237 3014
rect 56179 2974 56237 2980
rect 52298 2909 52862 2937
rect 52298 2897 52304 2909
rect 52912 2897 52918 2949
rect 52970 2937 52976 2949
rect 53680 2937 53686 2949
rect 52970 2909 53686 2937
rect 52970 2897 52976 2909
rect 53680 2897 53686 2909
rect 53738 2897 53744 2949
rect 54832 2897 54838 2949
rect 54890 2937 54896 2949
rect 56194 2937 56222 2974
rect 54890 2909 56222 2937
rect 54890 2897 54896 2909
rect 46387 2866 46445 2872
rect 46387 2863 46399 2866
rect 41218 2835 46399 2863
rect 46387 2832 46399 2835
rect 46433 2832 46445 2866
rect 46387 2826 46445 2832
rect 50032 2823 50038 2875
rect 50090 2823 50096 2875
rect 51763 2866 51821 2872
rect 51763 2832 51775 2866
rect 51809 2863 51821 2866
rect 52816 2863 52822 2875
rect 51809 2835 52822 2863
rect 51809 2832 51821 2835
rect 51763 2826 51821 2832
rect 52816 2823 52822 2835
rect 52874 2823 52880 2875
rect 53107 2866 53165 2872
rect 53107 2832 53119 2866
rect 53153 2832 53165 2866
rect 53107 2826 53165 2832
rect 43699 2792 43757 2798
rect 43699 2789 43711 2792
rect 34594 2761 43711 2789
rect 43699 2758 43711 2761
rect 43745 2758 43757 2792
rect 43699 2752 43757 2758
rect 46096 2749 46102 2801
rect 46154 2789 46160 2801
rect 46672 2789 46678 2801
rect 46154 2761 46678 2789
rect 46154 2749 46160 2761
rect 46672 2749 46678 2761
rect 46730 2749 46736 2801
rect 49075 2792 49133 2798
rect 49075 2758 49087 2792
rect 49121 2789 49133 2792
rect 53122 2789 53150 2826
rect 49121 2761 53150 2789
rect 49121 2758 49133 2761
rect 49075 2752 49133 2758
rect 1152 2690 58848 2712
rect 1152 2638 4294 2690
rect 4346 2638 4358 2690
rect 4410 2638 4422 2690
rect 4474 2638 4486 2690
rect 4538 2638 35014 2690
rect 35066 2638 35078 2690
rect 35130 2638 35142 2690
rect 35194 2638 35206 2690
rect 35258 2638 58848 2690
rect 1152 2616 58848 2638
rect 3952 2527 3958 2579
rect 4010 2567 4016 2579
rect 4240 2567 4246 2579
rect 4010 2539 4246 2567
rect 4010 2527 4016 2539
rect 4240 2527 4246 2539
rect 4298 2527 4304 2579
rect 4336 2527 4342 2579
rect 4394 2567 4400 2579
rect 4816 2567 4822 2579
rect 4394 2539 4822 2567
rect 4394 2527 4400 2539
rect 4816 2527 4822 2539
rect 4874 2527 4880 2579
rect 8752 2527 8758 2579
rect 8810 2567 8816 2579
rect 29776 2567 29782 2579
rect 8810 2539 29782 2567
rect 8810 2527 8816 2539
rect 29776 2527 29782 2539
rect 29834 2527 29840 2579
rect 35632 2527 35638 2579
rect 35690 2567 35696 2579
rect 36880 2567 36886 2579
rect 35690 2539 36886 2567
rect 35690 2527 35696 2539
rect 36880 2527 36886 2539
rect 36938 2527 36944 2579
rect 43216 2527 43222 2579
rect 43274 2567 43280 2579
rect 43984 2567 43990 2579
rect 43274 2539 43990 2567
rect 43274 2527 43280 2539
rect 43984 2527 43990 2539
rect 44042 2527 44048 2579
rect 20176 2453 20182 2505
rect 20234 2493 20240 2505
rect 20848 2493 20854 2505
rect 20234 2465 20854 2493
rect 20234 2453 20240 2465
rect 20848 2453 20854 2465
rect 20906 2453 20912 2505
rect 33808 2453 33814 2505
rect 33866 2493 33872 2505
rect 40816 2493 40822 2505
rect 33866 2465 40822 2493
rect 33866 2453 33872 2465
rect 40816 2453 40822 2465
rect 40874 2453 40880 2505
rect 33808 2305 33814 2357
rect 33866 2345 33872 2357
rect 34672 2345 34678 2357
rect 33866 2317 34678 2345
rect 33866 2305 33872 2317
rect 34672 2305 34678 2317
rect 34730 2305 34736 2357
rect 16240 2157 16246 2209
rect 16298 2197 16304 2209
rect 16432 2197 16438 2209
rect 16298 2169 16438 2197
rect 16298 2157 16304 2169
rect 16432 2157 16438 2169
rect 16490 2157 16496 2209
rect 4720 2009 4726 2061
rect 4778 2049 4784 2061
rect 5296 2049 5302 2061
rect 4778 2021 5302 2049
rect 4778 2009 4784 2021
rect 5296 2009 5302 2021
rect 5354 2009 5360 2061
rect 16528 1935 16534 1987
rect 16586 1975 16592 1987
rect 16720 1975 16726 1987
rect 16586 1947 16726 1975
rect 16586 1935 16592 1947
rect 16720 1935 16726 1947
rect 16778 1935 16784 1987
rect 4528 1861 4534 1913
rect 4586 1901 4592 1913
rect 4816 1901 4822 1913
rect 4586 1873 4822 1901
rect 4586 1861 4592 1873
rect 4816 1861 4822 1873
rect 4874 1861 4880 1913
rect 30352 1713 30358 1765
rect 30410 1753 30416 1765
rect 30640 1753 30646 1765
rect 30410 1725 30646 1753
rect 30410 1713 30416 1725
rect 30640 1713 30646 1725
rect 30698 1713 30704 1765
rect 50704 1713 50710 1765
rect 50762 1753 50768 1765
rect 50896 1753 50902 1765
rect 50762 1725 50902 1753
rect 50762 1713 50768 1725
rect 50896 1713 50902 1725
rect 50954 1713 50960 1765
rect 35344 1639 35350 1691
rect 35402 1639 35408 1691
rect 36304 1639 36310 1691
rect 36362 1639 36368 1691
rect 50512 1639 50518 1691
rect 50570 1679 50576 1691
rect 51088 1679 51094 1691
rect 50570 1651 51094 1679
rect 50570 1639 50576 1651
rect 51088 1639 51094 1651
rect 51146 1639 51152 1691
rect 35362 1395 35390 1639
rect 36322 1395 36350 1639
rect 50896 1565 50902 1617
rect 50954 1605 50960 1617
rect 51568 1605 51574 1617
rect 50954 1577 51574 1605
rect 50954 1565 50960 1577
rect 51568 1565 51574 1577
rect 51626 1565 51632 1617
rect 41008 1417 41014 1469
rect 41066 1457 41072 1469
rect 41296 1457 41302 1469
rect 41066 1429 41302 1457
rect 41066 1417 41072 1429
rect 41296 1417 41302 1429
rect 41354 1417 41360 1469
rect 35344 1343 35350 1395
rect 35402 1343 35408 1395
rect 36304 1343 36310 1395
rect 36362 1343 36368 1395
rect 33232 1269 33238 1321
rect 33290 1309 33296 1321
rect 33712 1309 33718 1321
rect 33290 1281 33718 1309
rect 33290 1269 33296 1281
rect 33712 1269 33718 1281
rect 33770 1269 33776 1321
rect 36112 1269 36118 1321
rect 36170 1309 36176 1321
rect 37264 1309 37270 1321
rect 36170 1281 37270 1309
rect 36170 1269 36176 1281
rect 37264 1269 37270 1281
rect 37322 1269 37328 1321
rect 34864 1195 34870 1247
rect 34922 1235 34928 1247
rect 35920 1235 35926 1247
rect 34922 1207 35926 1235
rect 34922 1195 34928 1207
rect 35920 1195 35926 1207
rect 35978 1195 35984 1247
<< via1 >>
rect 4294 57250 4346 57302
rect 4358 57250 4410 57302
rect 4422 57250 4474 57302
rect 4486 57250 4538 57302
rect 35014 57250 35066 57302
rect 35078 57250 35130 57302
rect 35142 57250 35194 57302
rect 35206 57250 35258 57302
rect 1750 56991 1802 57043
rect 214 56917 266 56969
rect 3286 56991 3338 57043
rect 4918 56917 4970 56969
rect 9622 56991 9674 57043
rect 11254 56991 11306 57043
rect 6454 56917 6506 56969
rect 8086 56960 8138 56969
rect 8086 56926 8095 56960
rect 8095 56926 8129 56960
rect 8129 56926 8138 56960
rect 8086 56917 8138 56926
rect 16438 56991 16490 57043
rect 18070 56991 18122 57043
rect 29110 56991 29162 57043
rect 12790 56917 12842 56969
rect 14422 56917 14474 56969
rect 15958 56917 16010 56969
rect 17494 56917 17546 56969
rect 19126 56917 19178 56969
rect 20662 56960 20714 56969
rect 20662 56926 20671 56960
rect 20671 56926 20705 56960
rect 20705 56926 20714 56960
rect 20662 56917 20714 56926
rect 22294 56917 22346 56969
rect 23830 56917 23882 56969
rect 25462 56917 25514 56969
rect 26998 56960 27050 56969
rect 26998 56926 27007 56960
rect 27007 56926 27041 56960
rect 27041 56926 27050 56960
rect 26998 56917 27050 56926
rect 28630 56917 28682 56969
rect 30166 56917 30218 56969
rect 31702 56917 31754 56969
rect 33334 56917 33386 56969
rect 34870 56917 34922 56969
rect 36502 56917 36554 56969
rect 41206 56917 41258 56969
rect 47542 56960 47594 56969
rect 47542 56926 47551 56960
rect 47551 56926 47585 56960
rect 47585 56926 47594 56960
rect 47542 56917 47594 56926
rect 52246 56917 52298 56969
rect 1750 56886 1802 56895
rect 1750 56852 1759 56886
rect 1759 56852 1793 56886
rect 1793 56852 1802 56886
rect 1750 56843 1802 56852
rect 2614 56886 2666 56895
rect 2614 56852 2623 56886
rect 2623 56852 2657 56886
rect 2657 56852 2666 56886
rect 2614 56843 2666 56852
rect 8278 56843 8330 56895
rect 11254 56886 11306 56895
rect 11254 56852 11263 56886
rect 11263 56852 11297 56886
rect 11297 56852 11306 56886
rect 11254 56843 11306 56852
rect 12214 56843 12266 56895
rect 14038 56886 14090 56895
rect 14038 56852 14047 56886
rect 14047 56852 14081 56886
rect 14081 56852 14090 56886
rect 14038 56843 14090 56852
rect 16150 56886 16202 56895
rect 16150 56852 16159 56886
rect 16159 56852 16193 56886
rect 16193 56852 16202 56886
rect 16150 56843 16202 56852
rect 6454 56769 6506 56821
rect 12406 56769 12458 56821
rect 21622 56886 21674 56895
rect 21622 56852 21631 56886
rect 21631 56852 21665 56886
rect 21665 56852 21674 56886
rect 21622 56843 21674 56852
rect 23350 56886 23402 56895
rect 23350 56852 23359 56886
rect 23359 56852 23393 56886
rect 23393 56852 23402 56886
rect 23350 56843 23402 56852
rect 26326 56843 26378 56895
rect 28822 56886 28874 56895
rect 28822 56852 28831 56886
rect 28831 56852 28865 56886
rect 28865 56852 28874 56886
rect 28822 56843 28874 56852
rect 31894 56886 31946 56895
rect 31894 56852 31903 56886
rect 31903 56852 31937 56886
rect 31937 56852 31946 56886
rect 31894 56843 31946 56852
rect 32758 56886 32810 56895
rect 32758 56852 32767 56886
rect 32767 56852 32801 56886
rect 32801 56852 32810 56886
rect 32758 56843 32810 56852
rect 34102 56886 34154 56895
rect 34102 56852 34111 56886
rect 34111 56852 34145 56886
rect 34145 56852 34154 56886
rect 34102 56843 34154 56852
rect 38038 56843 38090 56895
rect 39670 56843 39722 56895
rect 34870 56769 34922 56821
rect 42838 56843 42890 56895
rect 44374 56843 44426 56895
rect 45910 56843 45962 56895
rect 49078 56843 49130 56895
rect 50710 56843 50762 56895
rect 53878 56843 53930 56895
rect 55414 56843 55466 56895
rect 58582 56843 58634 56895
rect 9814 56738 9866 56747
rect 9814 56704 9823 56738
rect 9823 56704 9857 56738
rect 9857 56704 9866 56738
rect 9814 56695 9866 56704
rect 37942 56738 37994 56747
rect 37942 56704 37951 56738
rect 37951 56704 37985 56738
rect 37985 56704 37994 56738
rect 37942 56695 37994 56704
rect 39766 56738 39818 56747
rect 39766 56704 39775 56738
rect 39775 56704 39809 56738
rect 39809 56704 39818 56738
rect 39766 56695 39818 56704
rect 40438 56738 40490 56747
rect 40438 56704 40447 56738
rect 40447 56704 40481 56738
rect 40481 56704 40490 56738
rect 40438 56695 40490 56704
rect 40822 56738 40874 56747
rect 40822 56704 40831 56738
rect 40831 56704 40865 56738
rect 40865 56704 40874 56738
rect 40822 56695 40874 56704
rect 42934 56738 42986 56747
rect 42934 56704 42943 56738
rect 42943 56704 42977 56738
rect 42977 56704 42986 56738
rect 42934 56695 42986 56704
rect 44758 56738 44810 56747
rect 44758 56704 44767 56738
rect 44767 56704 44801 56738
rect 44801 56704 44810 56738
rect 44758 56695 44810 56704
rect 46102 56695 46154 56747
rect 48694 56738 48746 56747
rect 48694 56704 48703 56738
rect 48703 56704 48737 56738
rect 48737 56704 48746 56738
rect 48694 56695 48746 56704
rect 50806 56738 50858 56747
rect 50806 56704 50815 56738
rect 50815 56704 50849 56738
rect 50849 56704 50858 56738
rect 50806 56695 50858 56704
rect 53878 56695 53930 56747
rect 55510 56738 55562 56747
rect 55510 56704 55519 56738
rect 55519 56704 55553 56738
rect 55553 56704 55562 56738
rect 55510 56695 55562 56704
rect 56758 56738 56810 56747
rect 56758 56704 56767 56738
rect 56767 56704 56801 56738
rect 56801 56704 56810 56738
rect 56758 56695 56810 56704
rect 19654 56584 19706 56636
rect 19718 56584 19770 56636
rect 19782 56584 19834 56636
rect 19846 56584 19898 56636
rect 50374 56584 50426 56636
rect 50438 56584 50490 56636
rect 50502 56584 50554 56636
rect 50566 56584 50618 56636
rect 694 56473 746 56525
rect 2230 56473 2282 56525
rect 2806 56473 2858 56525
rect 3862 56473 3914 56525
rect 5398 56473 5450 56525
rect 5974 56473 6026 56525
rect 7030 56473 7082 56525
rect 8566 56473 8618 56525
rect 10198 56473 10250 56525
rect 10678 56473 10730 56525
rect 11734 56473 11786 56525
rect 12310 56473 12362 56525
rect 13366 56473 13418 56525
rect 14902 56473 14954 56525
rect 17014 56473 17066 56525
rect 18742 56516 18794 56525
rect 18742 56482 18751 56516
rect 18751 56482 18785 56516
rect 18785 56482 18794 56516
rect 18742 56473 18794 56482
rect 19990 56473 20042 56525
rect 21238 56473 21290 56525
rect 21718 56473 21770 56525
rect 22774 56473 22826 56525
rect 24406 56473 24458 56525
rect 25942 56473 25994 56525
rect 26518 56473 26570 56525
rect 27574 56473 27626 56525
rect 28054 56473 28106 56525
rect 29686 56516 29738 56525
rect 29686 56482 29695 56516
rect 29695 56482 29729 56516
rect 29729 56482 29738 56516
rect 29686 56473 29738 56482
rect 30646 56473 30698 56525
rect 32278 56473 32330 56525
rect 32854 56473 32906 56525
rect 33814 56473 33866 56525
rect 34390 56473 34442 56525
rect 35446 56473 35498 56525
rect 36022 56399 36074 56451
rect 37558 56473 37610 56525
rect 38614 56473 38666 56525
rect 40150 56473 40202 56525
rect 41782 56473 41834 56525
rect 42262 56473 42314 56525
rect 43318 56473 43370 56525
rect 43894 56473 43946 56525
rect 44950 56473 45002 56525
rect 46486 56473 46538 56525
rect 48022 56473 48074 56525
rect 48598 56473 48650 56525
rect 49654 56473 49706 56525
rect 50134 56473 50186 56525
rect 52822 56473 52874 56525
rect 53302 56473 53354 56525
rect 54358 56473 54410 56525
rect 54934 56473 54986 56525
rect 55990 56516 56042 56525
rect 55990 56482 55999 56516
rect 55999 56482 56033 56516
rect 56033 56482 56042 56516
rect 55990 56473 56042 56482
rect 39574 56399 39626 56451
rect 56758 56399 56810 56451
rect 42358 56325 42410 56377
rect 47062 56325 47114 56377
rect 12502 56251 12554 56303
rect 13750 56251 13802 56303
rect 43894 56251 43946 56303
rect 46870 56251 46922 56303
rect 1846 56177 1898 56229
rect 2710 56177 2762 56229
rect 2998 56220 3050 56229
rect 2998 56186 3007 56220
rect 3007 56186 3041 56220
rect 3041 56186 3050 56220
rect 2998 56177 3050 56186
rect 5014 56177 5066 56229
rect 5206 56220 5258 56229
rect 5206 56186 5215 56220
rect 5215 56186 5249 56220
rect 5249 56186 5258 56220
rect 5206 56177 5258 56186
rect 6358 56220 6410 56229
rect 6358 56186 6367 56220
rect 6367 56186 6401 56220
rect 6401 56186 6410 56220
rect 6358 56177 6410 56186
rect 8566 56220 8618 56229
rect 8566 56186 8575 56220
rect 8575 56186 8609 56220
rect 8609 56186 8618 56220
rect 8566 56177 8618 56186
rect 10390 56220 10442 56229
rect 10390 56186 10399 56220
rect 10399 56186 10433 56220
rect 10433 56186 10442 56220
rect 10390 56177 10442 56186
rect 10774 56220 10826 56229
rect 10774 56186 10783 56220
rect 10783 56186 10817 56220
rect 10817 56186 10826 56220
rect 10774 56177 10826 56186
rect 11926 56220 11978 56229
rect 11926 56186 11935 56220
rect 11935 56186 11969 56220
rect 11969 56186 11978 56220
rect 11926 56177 11978 56186
rect 12694 56220 12746 56229
rect 12694 56186 12703 56220
rect 12703 56186 12737 56220
rect 12737 56186 12746 56220
rect 12694 56177 12746 56186
rect 13558 56220 13610 56229
rect 13558 56186 13567 56220
rect 13567 56186 13601 56220
rect 13601 56186 13610 56220
rect 13558 56177 13610 56186
rect 15190 56177 15242 56229
rect 16822 56220 16874 56229
rect 15382 56103 15434 56155
rect 16822 56186 16831 56220
rect 16831 56186 16865 56220
rect 16865 56186 16874 56220
rect 16822 56177 16874 56186
rect 18646 56220 18698 56229
rect 18646 56186 18655 56220
rect 18655 56186 18689 56220
rect 18689 56186 18698 56220
rect 18646 56177 18698 56186
rect 20854 56177 20906 56229
rect 21430 56220 21482 56229
rect 21430 56186 21439 56220
rect 21439 56186 21473 56220
rect 21473 56186 21482 56220
rect 21430 56177 21482 56186
rect 22102 56220 22154 56229
rect 22102 56186 22111 56220
rect 22111 56186 22145 56220
rect 22145 56186 22154 56220
rect 22102 56177 22154 56186
rect 22966 56220 23018 56229
rect 22966 56186 22975 56220
rect 22975 56186 23009 56220
rect 23009 56186 23018 56220
rect 24406 56220 24458 56229
rect 22966 56177 23018 56186
rect 24406 56186 24415 56220
rect 24415 56186 24449 56220
rect 24449 56186 24458 56220
rect 24406 56177 24458 56186
rect 26134 56220 26186 56229
rect 26134 56186 26143 56220
rect 26143 56186 26177 56220
rect 26177 56186 26186 56220
rect 26134 56177 26186 56186
rect 26902 56220 26954 56229
rect 26902 56186 26911 56220
rect 26911 56186 26945 56220
rect 26945 56186 26954 56220
rect 26902 56177 26954 56186
rect 27766 56220 27818 56229
rect 27766 56186 27775 56220
rect 27775 56186 27809 56220
rect 27809 56186 27818 56220
rect 27766 56177 27818 56186
rect 28150 56220 28202 56229
rect 28150 56186 28159 56220
rect 28159 56186 28193 56220
rect 28193 56186 28202 56220
rect 28150 56177 28202 56186
rect 29590 56220 29642 56229
rect 29590 56186 29599 56220
rect 29599 56186 29633 56220
rect 29633 56186 29642 56220
rect 29590 56177 29642 56186
rect 30934 56220 30986 56229
rect 30934 56186 30943 56220
rect 30943 56186 30977 56220
rect 30977 56186 30986 56220
rect 30934 56177 30986 56186
rect 31318 56220 31370 56229
rect 31318 56186 31327 56220
rect 31327 56186 31361 56220
rect 31361 56186 31370 56220
rect 31318 56177 31370 56186
rect 32470 56220 32522 56229
rect 31222 56103 31274 56155
rect 32470 56186 32479 56220
rect 32479 56186 32513 56220
rect 32513 56186 32522 56220
rect 32470 56177 32522 56186
rect 34006 56220 34058 56229
rect 34006 56186 34015 56220
rect 34015 56186 34049 56220
rect 34049 56186 34058 56220
rect 34006 56177 34058 56186
rect 34774 56220 34826 56229
rect 34774 56186 34783 56220
rect 34783 56186 34817 56220
rect 34817 56186 34826 56220
rect 34774 56177 34826 56186
rect 35350 56177 35402 56229
rect 36886 56220 36938 56229
rect 36886 56186 36895 56220
rect 36895 56186 36929 56220
rect 36929 56186 36938 56220
rect 36886 56177 36938 56186
rect 37462 56220 37514 56229
rect 37462 56186 37471 56220
rect 37471 56186 37505 56220
rect 37505 56186 37514 56220
rect 37462 56177 37514 56186
rect 38422 56220 38474 56229
rect 38422 56186 38431 56220
rect 38431 56186 38465 56220
rect 38465 56186 38474 56220
rect 38422 56177 38474 56186
rect 39862 56220 39914 56229
rect 39862 56186 39871 56220
rect 39871 56186 39905 56220
rect 39905 56186 39914 56220
rect 39862 56177 39914 56186
rect 42070 56177 42122 56229
rect 42646 56220 42698 56229
rect 42646 56186 42655 56220
rect 42655 56186 42689 56220
rect 42689 56186 42698 56220
rect 42646 56177 42698 56186
rect 43510 56220 43562 56229
rect 43510 56186 43519 56220
rect 43519 56186 43553 56220
rect 43553 56186 43562 56220
rect 43510 56177 43562 56186
rect 44182 56220 44234 56229
rect 44182 56186 44191 56220
rect 44191 56186 44225 56220
rect 44225 56186 44234 56220
rect 44182 56177 44234 56186
rect 46678 56220 46730 56229
rect 46678 56186 46687 56220
rect 46687 56186 46721 56220
rect 46721 56186 46730 56220
rect 46678 56177 46730 56186
rect 48214 56220 48266 56229
rect 48214 56186 48223 56220
rect 48223 56186 48257 56220
rect 48257 56186 48266 56220
rect 48214 56177 48266 56186
rect 48598 56220 48650 56229
rect 48598 56186 48607 56220
rect 48607 56186 48641 56220
rect 48641 56186 48650 56220
rect 48598 56177 48650 56186
rect 50230 56220 50282 56229
rect 50230 56186 50239 56220
rect 50239 56186 50273 56220
rect 50273 56186 50282 56220
rect 50230 56177 50282 56186
rect 51286 56177 51338 56229
rect 57046 56251 57098 56303
rect 52918 56220 52970 56229
rect 51190 56103 51242 56155
rect 52918 56186 52927 56220
rect 52927 56186 52961 56220
rect 52961 56186 52970 56220
rect 52918 56177 52970 56186
rect 53974 56220 54026 56229
rect 53974 56186 53983 56220
rect 53983 56186 54017 56220
rect 54017 56186 54026 56220
rect 53974 56177 54026 56186
rect 54550 56220 54602 56229
rect 54550 56186 54559 56220
rect 54559 56186 54593 56220
rect 54593 56186 54602 56220
rect 54550 56177 54602 56186
rect 54934 56220 54986 56229
rect 54934 56186 54943 56220
rect 54943 56186 54977 56220
rect 54977 56186 54986 56220
rect 54934 56177 54986 56186
rect 36982 56029 37034 56081
rect 40822 56029 40874 56081
rect 4294 55918 4346 55970
rect 4358 55918 4410 55970
rect 4422 55918 4474 55970
rect 4486 55918 4538 55970
rect 35014 55918 35066 55970
rect 35078 55918 35130 55970
rect 35142 55918 35194 55970
rect 35206 55918 35258 55970
rect 1174 55659 1226 55711
rect 4630 55659 4682 55711
rect 7510 55659 7562 55711
rect 9142 55659 9194 55711
rect 13846 55659 13898 55711
rect 20182 55659 20234 55711
rect 23446 55702 23498 55711
rect 23446 55668 23455 55702
rect 23455 55668 23489 55702
rect 23489 55668 23498 55702
rect 23446 55659 23498 55668
rect 24886 55659 24938 55711
rect 20566 55585 20618 55637
rect 4630 55511 4682 55563
rect 14134 55511 14186 55563
rect 26134 55585 26186 55637
rect 39094 55659 39146 55711
rect 40726 55659 40778 55711
rect 45430 55659 45482 55711
rect 46966 55659 47018 55711
rect 51766 55659 51818 55711
rect 56470 55659 56522 55711
rect 57526 55659 57578 55711
rect 45334 55585 45386 55637
rect 24310 55511 24362 55563
rect 24982 55554 25034 55563
rect 24982 55520 24991 55554
rect 24991 55520 25025 55554
rect 25025 55520 25034 55554
rect 24982 55511 25034 55520
rect 39190 55554 39242 55563
rect 39190 55520 39199 55554
rect 39199 55520 39233 55554
rect 39233 55520 39242 55554
rect 39190 55511 39242 55520
rect 40822 55511 40874 55563
rect 51958 55554 52010 55563
rect 1942 55406 1994 55415
rect 1942 55372 1951 55406
rect 1951 55372 1985 55406
rect 1985 55372 1994 55406
rect 1942 55363 1994 55372
rect 7318 55406 7370 55415
rect 7318 55372 7327 55406
rect 7327 55372 7361 55406
rect 7361 55372 7370 55406
rect 7318 55363 7370 55372
rect 8950 55406 9002 55415
rect 8950 55372 8959 55406
rect 8959 55372 8993 55406
rect 8993 55372 9002 55406
rect 8950 55363 9002 55372
rect 17398 55406 17450 55415
rect 17398 55372 17407 55406
rect 17407 55372 17441 55406
rect 17441 55372 17450 55406
rect 17398 55363 17450 55372
rect 20086 55406 20138 55415
rect 20086 55372 20095 55406
rect 20095 55372 20129 55406
rect 20129 55372 20138 55406
rect 20086 55363 20138 55372
rect 20758 55406 20810 55415
rect 20758 55372 20767 55406
rect 20767 55372 20801 55406
rect 20801 55372 20810 55406
rect 20758 55363 20810 55372
rect 51958 55520 51967 55554
rect 51967 55520 52001 55554
rect 52001 55520 52010 55554
rect 51958 55511 52010 55520
rect 45814 55406 45866 55415
rect 45814 55372 45823 55406
rect 45823 55372 45857 55406
rect 45857 55372 45866 55406
rect 45814 55363 45866 55372
rect 55606 55406 55658 55415
rect 55606 55372 55615 55406
rect 55615 55372 55649 55406
rect 55649 55372 55658 55406
rect 55606 55363 55658 55372
rect 56278 55406 56330 55415
rect 56278 55372 56287 55406
rect 56287 55372 56321 55406
rect 56321 55372 56330 55406
rect 57334 55406 57386 55415
rect 56278 55363 56330 55372
rect 57334 55372 57343 55406
rect 57343 55372 57377 55406
rect 57377 55372 57386 55406
rect 57334 55363 57386 55372
rect 19654 55252 19706 55304
rect 19718 55252 19770 55304
rect 19782 55252 19834 55304
rect 19846 55252 19898 55304
rect 50374 55252 50426 55304
rect 50438 55252 50490 55304
rect 50502 55252 50554 55304
rect 50566 55252 50618 55304
rect 59158 55141 59210 55193
rect 15094 55067 15146 55119
rect 55606 55067 55658 55119
rect 42358 55036 42410 55045
rect 42358 55002 42367 55036
rect 42367 55002 42401 55036
rect 42401 55002 42410 55036
rect 42358 54993 42410 55002
rect 57814 54888 57866 54897
rect 57814 54854 57823 54888
rect 57823 54854 57857 54888
rect 57857 54854 57866 54888
rect 57814 54845 57866 54854
rect 5014 54771 5066 54823
rect 15286 54697 15338 54749
rect 20470 54740 20522 54749
rect 20470 54706 20479 54740
rect 20479 54706 20513 54740
rect 20513 54706 20522 54740
rect 20470 54697 20522 54706
rect 22390 54740 22442 54749
rect 22390 54706 22399 54740
rect 22399 54706 22433 54740
rect 22433 54706 22442 54740
rect 22390 54697 22442 54706
rect 4294 54586 4346 54638
rect 4358 54586 4410 54638
rect 4422 54586 4474 54638
rect 4486 54586 4538 54638
rect 35014 54586 35066 54638
rect 35078 54586 35130 54638
rect 35142 54586 35194 54638
rect 35206 54586 35258 54638
rect 58102 54327 58154 54379
rect 58102 54074 58154 54083
rect 58102 54040 58111 54074
rect 58111 54040 58145 54074
rect 58145 54040 58154 54074
rect 58102 54031 58154 54040
rect 19654 53920 19706 53972
rect 19718 53920 19770 53972
rect 19782 53920 19834 53972
rect 19846 53920 19898 53972
rect 50374 53920 50426 53972
rect 50438 53920 50490 53972
rect 50502 53920 50554 53972
rect 50566 53920 50618 53972
rect 59638 53809 59690 53861
rect 57718 53365 57770 53417
rect 4294 53254 4346 53306
rect 4358 53254 4410 53306
rect 4422 53254 4474 53306
rect 4486 53254 4538 53306
rect 35014 53254 35066 53306
rect 35078 53254 35130 53306
rect 35142 53254 35194 53306
rect 35206 53254 35258 53306
rect 35350 52995 35402 53047
rect 14998 52847 15050 52899
rect 26902 52847 26954 52899
rect 19654 52588 19706 52640
rect 19718 52588 19770 52640
rect 19782 52588 19834 52640
rect 19846 52588 19898 52640
rect 50374 52588 50426 52640
rect 50438 52588 50490 52640
rect 50502 52588 50554 52640
rect 50566 52588 50618 52640
rect 4294 51922 4346 51974
rect 4358 51922 4410 51974
rect 4422 51922 4474 51974
rect 4486 51922 4538 51974
rect 35014 51922 35066 51974
rect 35078 51922 35130 51974
rect 35142 51922 35194 51974
rect 35206 51922 35258 51974
rect 19414 51515 19466 51567
rect 54550 51367 54602 51419
rect 19654 51256 19706 51308
rect 19718 51256 19770 51308
rect 19782 51256 19834 51308
rect 19846 51256 19898 51308
rect 50374 51256 50426 51308
rect 50438 51256 50490 51308
rect 50502 51256 50554 51308
rect 50566 51256 50618 51308
rect 12502 51188 12554 51197
rect 12502 51154 12511 51188
rect 12511 51154 12545 51188
rect 12545 51154 12554 51188
rect 12502 51145 12554 51154
rect 11926 50849 11978 50901
rect 55030 50701 55082 50753
rect 56854 50701 56906 50753
rect 4294 50590 4346 50642
rect 4358 50590 4410 50642
rect 4422 50590 4474 50642
rect 4486 50590 4538 50642
rect 35014 50590 35066 50642
rect 35078 50590 35130 50642
rect 35142 50590 35194 50642
rect 35206 50590 35258 50642
rect 54934 50405 54986 50457
rect 40918 50035 40970 50087
rect 19654 49924 19706 49976
rect 19718 49924 19770 49976
rect 19782 49924 19834 49976
rect 19846 49924 19898 49976
rect 50374 49924 50426 49976
rect 50438 49924 50490 49976
rect 50502 49924 50554 49976
rect 50566 49924 50618 49976
rect 32470 49517 32522 49569
rect 44854 49412 44906 49421
rect 44854 49378 44863 49412
rect 44863 49378 44897 49412
rect 44897 49378 44906 49412
rect 44854 49369 44906 49378
rect 48118 49412 48170 49421
rect 48118 49378 48127 49412
rect 48127 49378 48161 49412
rect 48161 49378 48170 49412
rect 48118 49369 48170 49378
rect 4294 49258 4346 49310
rect 4358 49258 4410 49310
rect 4422 49258 4474 49310
rect 4486 49258 4538 49310
rect 35014 49258 35066 49310
rect 35078 49258 35130 49310
rect 35142 49258 35194 49310
rect 35206 49258 35258 49310
rect 7222 49042 7274 49051
rect 7222 49008 7231 49042
rect 7231 49008 7265 49042
rect 7265 49008 7274 49042
rect 7222 48999 7274 49008
rect 29686 48851 29738 48903
rect 3574 48703 3626 48755
rect 43510 48703 43562 48755
rect 19654 48592 19706 48644
rect 19718 48592 19770 48644
rect 19782 48592 19834 48644
rect 19846 48592 19898 48644
rect 50374 48592 50426 48644
rect 50438 48592 50490 48644
rect 50502 48592 50554 48644
rect 50566 48592 50618 48644
rect 4726 48037 4778 48089
rect 48886 48037 48938 48089
rect 4294 47926 4346 47978
rect 4358 47926 4410 47978
rect 4422 47926 4474 47978
rect 4486 47926 4538 47978
rect 35014 47926 35066 47978
rect 35078 47926 35130 47978
rect 35142 47926 35194 47978
rect 35206 47926 35258 47978
rect 39670 47593 39722 47645
rect 48214 47519 48266 47571
rect 19654 47260 19706 47312
rect 19718 47260 19770 47312
rect 19782 47260 19834 47312
rect 19846 47260 19898 47312
rect 50374 47260 50426 47312
rect 50438 47260 50490 47312
rect 50502 47260 50554 47312
rect 50566 47260 50618 47312
rect 43894 46853 43946 46905
rect 16630 46779 16682 46831
rect 4822 46748 4874 46757
rect 4822 46714 4831 46748
rect 4831 46714 4865 46748
rect 4865 46714 4874 46748
rect 4822 46705 4874 46714
rect 19990 46705 20042 46757
rect 45430 46748 45482 46757
rect 45430 46714 45439 46748
rect 45439 46714 45473 46748
rect 45473 46714 45482 46748
rect 45430 46705 45482 46714
rect 4294 46594 4346 46646
rect 4358 46594 4410 46646
rect 4422 46594 4474 46646
rect 4486 46594 4538 46646
rect 35014 46594 35066 46646
rect 35078 46594 35130 46646
rect 35142 46594 35194 46646
rect 35206 46594 35258 46646
rect 4822 46483 4874 46535
rect 57142 46483 57194 46535
rect 27958 46156 28010 46165
rect 27958 46122 27967 46156
rect 27967 46122 28001 46156
rect 28001 46122 28010 46156
rect 27958 46113 28010 46122
rect 46966 46039 47018 46091
rect 19654 45928 19706 45980
rect 19718 45928 19770 45980
rect 19782 45928 19834 45980
rect 19846 45928 19898 45980
rect 50374 45928 50426 45980
rect 50438 45928 50490 45980
rect 50502 45928 50554 45980
rect 50566 45928 50618 45980
rect 20470 45373 20522 45425
rect 31606 45373 31658 45425
rect 4294 45262 4346 45314
rect 4358 45262 4410 45314
rect 4422 45262 4474 45314
rect 4486 45262 4538 45314
rect 35014 45262 35066 45314
rect 35078 45262 35130 45314
rect 35142 45262 35194 45314
rect 35206 45262 35258 45314
rect 12118 44855 12170 44907
rect 19654 44596 19706 44648
rect 19718 44596 19770 44648
rect 19782 44596 19834 44648
rect 19846 44596 19898 44648
rect 50374 44596 50426 44648
rect 50438 44596 50490 44648
rect 50502 44596 50554 44648
rect 50566 44596 50618 44648
rect 17974 44041 18026 44093
rect 47734 44084 47786 44093
rect 47734 44050 47743 44084
rect 47743 44050 47777 44084
rect 47777 44050 47786 44084
rect 47734 44041 47786 44050
rect 4294 43930 4346 43982
rect 4358 43930 4410 43982
rect 4422 43930 4474 43982
rect 4486 43930 4538 43982
rect 35014 43930 35066 43982
rect 35078 43930 35130 43982
rect 35142 43930 35194 43982
rect 35206 43930 35258 43982
rect 25654 43819 25706 43871
rect 47734 43819 47786 43871
rect 54070 43597 54122 43649
rect 13654 43523 13706 43575
rect 22294 43375 22346 43427
rect 52246 43523 52298 43575
rect 19654 43264 19706 43316
rect 19718 43264 19770 43316
rect 19782 43264 19834 43316
rect 19846 43264 19898 43316
rect 50374 43264 50426 43316
rect 50438 43264 50490 43316
rect 50502 43264 50554 43316
rect 50566 43264 50618 43316
rect 11446 42783 11498 42835
rect 11350 42709 11402 42761
rect 25942 42752 25994 42761
rect 25942 42718 25951 42752
rect 25951 42718 25985 42752
rect 25985 42718 25994 42752
rect 25942 42709 25994 42718
rect 4294 42598 4346 42650
rect 4358 42598 4410 42650
rect 4422 42598 4474 42650
rect 4486 42598 4538 42650
rect 35014 42598 35066 42650
rect 35078 42598 35130 42650
rect 35142 42598 35194 42650
rect 35206 42598 35258 42650
rect 11350 42487 11402 42539
rect 26134 42487 26186 42539
rect 14134 42265 14186 42317
rect 16534 42234 16586 42243
rect 16534 42200 16543 42234
rect 16543 42200 16577 42234
rect 16577 42200 16586 42234
rect 16534 42191 16586 42200
rect 19654 41932 19706 41984
rect 19718 41932 19770 41984
rect 19782 41932 19834 41984
rect 19846 41932 19898 41984
rect 50374 41932 50426 41984
rect 50438 41932 50490 41984
rect 50502 41932 50554 41984
rect 50566 41932 50618 41984
rect 22966 41747 23018 41799
rect 25174 41377 25226 41429
rect 4294 41266 4346 41318
rect 4358 41266 4410 41318
rect 4422 41266 4474 41318
rect 4486 41266 4538 41318
rect 35014 41266 35066 41318
rect 35078 41266 35130 41318
rect 35142 41266 35194 41318
rect 35206 41266 35258 41318
rect 28918 40859 28970 40911
rect 33910 40754 33962 40763
rect 33910 40720 33919 40754
rect 33919 40720 33953 40754
rect 33953 40720 33962 40754
rect 48310 40859 48362 40911
rect 33910 40711 33962 40720
rect 19654 40600 19706 40652
rect 19718 40600 19770 40652
rect 19782 40600 19834 40652
rect 19846 40600 19898 40652
rect 50374 40600 50426 40652
rect 50438 40600 50490 40652
rect 50502 40600 50554 40652
rect 50566 40600 50618 40652
rect 46870 40489 46922 40541
rect 25078 40045 25130 40097
rect 57238 40045 57290 40097
rect 4294 39934 4346 39986
rect 4358 39934 4410 39986
rect 4422 39934 4474 39986
rect 4486 39934 4538 39986
rect 35014 39934 35066 39986
rect 35078 39934 35130 39986
rect 35142 39934 35194 39986
rect 35206 39934 35258 39986
rect 23734 39823 23786 39875
rect 57238 39823 57290 39875
rect 57910 39379 57962 39431
rect 19654 39268 19706 39320
rect 19718 39268 19770 39320
rect 19782 39268 19834 39320
rect 19846 39268 19898 39320
rect 50374 39268 50426 39320
rect 50438 39268 50490 39320
rect 50502 39268 50554 39320
rect 50566 39268 50618 39320
rect 32758 39157 32810 39209
rect 1846 38861 1898 38913
rect 10678 38756 10730 38765
rect 10678 38722 10687 38756
rect 10687 38722 10721 38756
rect 10721 38722 10730 38756
rect 10678 38713 10730 38722
rect 30550 38713 30602 38765
rect 31510 38713 31562 38765
rect 57622 38756 57674 38765
rect 57622 38722 57631 38756
rect 57631 38722 57665 38756
rect 57665 38722 57674 38756
rect 57622 38713 57674 38722
rect 4294 38602 4346 38654
rect 4358 38602 4410 38654
rect 4422 38602 4474 38654
rect 4486 38602 4538 38654
rect 35014 38602 35066 38654
rect 35078 38602 35130 38654
rect 35142 38602 35194 38654
rect 35206 38602 35258 38654
rect 12694 38195 12746 38247
rect 13846 38121 13898 38173
rect 32662 38047 32714 38099
rect 19654 37936 19706 37988
rect 19718 37936 19770 37988
rect 19782 37936 19834 37988
rect 19846 37936 19898 37988
rect 50374 37936 50426 37988
rect 50438 37936 50490 37988
rect 50502 37936 50554 37988
rect 50566 37936 50618 37988
rect 5014 37424 5066 37433
rect 5014 37390 5023 37424
rect 5023 37390 5057 37424
rect 5057 37390 5066 37424
rect 5014 37381 5066 37390
rect 6070 37424 6122 37433
rect 6070 37390 6079 37424
rect 6079 37390 6113 37424
rect 6113 37390 6122 37424
rect 6070 37381 6122 37390
rect 30934 37381 30986 37433
rect 4294 37270 4346 37322
rect 4358 37270 4410 37322
rect 4422 37270 4474 37322
rect 4486 37270 4538 37322
rect 35014 37270 35066 37322
rect 35078 37270 35130 37322
rect 35142 37270 35194 37322
rect 35206 37270 35258 37322
rect 5014 37159 5066 37211
rect 52918 37159 52970 37211
rect 14902 36906 14954 36915
rect 14902 36872 14911 36906
rect 14911 36872 14945 36906
rect 14945 36872 14954 36906
rect 14902 36863 14954 36872
rect 18454 36715 18506 36767
rect 19654 36604 19706 36656
rect 19718 36604 19770 36656
rect 19782 36604 19834 36656
rect 19846 36604 19898 36656
rect 50374 36604 50426 36656
rect 50438 36604 50490 36656
rect 50502 36604 50554 36656
rect 50566 36604 50618 36656
rect 14902 36493 14954 36545
rect 32374 36493 32426 36545
rect 19510 36197 19562 36249
rect 2902 36049 2954 36101
rect 12502 36049 12554 36101
rect 18646 36123 18698 36175
rect 17878 36049 17930 36101
rect 44374 36092 44426 36101
rect 44374 36058 44383 36092
rect 44383 36058 44417 36092
rect 44417 36058 44426 36092
rect 44374 36049 44426 36058
rect 4294 35938 4346 35990
rect 4358 35938 4410 35990
rect 4422 35938 4474 35990
rect 4486 35938 4538 35990
rect 35014 35938 35066 35990
rect 35078 35938 35130 35990
rect 35142 35938 35194 35990
rect 35206 35938 35258 35990
rect 3286 35531 3338 35583
rect 20662 35574 20714 35583
rect 20662 35540 20671 35574
rect 20671 35540 20705 35574
rect 20705 35540 20714 35574
rect 20662 35531 20714 35540
rect 21718 35531 21770 35583
rect 32566 35531 32618 35583
rect 56662 35383 56714 35435
rect 19654 35272 19706 35324
rect 19718 35272 19770 35324
rect 19782 35272 19834 35324
rect 19846 35272 19898 35324
rect 50374 35272 50426 35324
rect 50438 35272 50490 35324
rect 50502 35272 50554 35324
rect 50566 35272 50618 35324
rect 40822 34791 40874 34843
rect 26806 34717 26858 34769
rect 31414 34760 31466 34769
rect 31414 34726 31423 34760
rect 31423 34726 31457 34760
rect 31457 34726 31466 34760
rect 31414 34717 31466 34726
rect 53206 34760 53258 34769
rect 53206 34726 53215 34760
rect 53215 34726 53249 34760
rect 53249 34726 53258 34760
rect 53206 34717 53258 34726
rect 57046 34760 57098 34769
rect 57046 34726 57055 34760
rect 57055 34726 57089 34760
rect 57089 34726 57098 34760
rect 57046 34717 57098 34726
rect 4294 34606 4346 34658
rect 4358 34606 4410 34658
rect 4422 34606 4474 34658
rect 4486 34606 4538 34658
rect 35014 34606 35066 34658
rect 35078 34606 35130 34658
rect 35142 34606 35194 34658
rect 35206 34606 35258 34658
rect 24406 34273 24458 34325
rect 53398 34125 53450 34177
rect 19654 33940 19706 33992
rect 19718 33940 19770 33992
rect 19782 33940 19834 33992
rect 19846 33940 19898 33992
rect 50374 33940 50426 33992
rect 50438 33940 50490 33992
rect 50502 33940 50554 33992
rect 50566 33940 50618 33992
rect 21718 33829 21770 33881
rect 51478 33829 51530 33881
rect 56278 33459 56330 33511
rect 10582 33385 10634 33437
rect 38134 33385 38186 33437
rect 4294 33274 4346 33326
rect 4358 33274 4410 33326
rect 4422 33274 4474 33326
rect 4486 33274 4538 33326
rect 35014 33274 35066 33326
rect 35078 33274 35130 33326
rect 35142 33274 35194 33326
rect 35206 33274 35258 33326
rect 10390 32719 10442 32771
rect 19654 32608 19706 32660
rect 19718 32608 19770 32660
rect 19782 32608 19834 32660
rect 19846 32608 19898 32660
rect 50374 32608 50426 32660
rect 50438 32608 50490 32660
rect 50502 32608 50554 32660
rect 50566 32608 50618 32660
rect 51958 32127 52010 32179
rect 24502 32053 24554 32105
rect 27382 32096 27434 32105
rect 27382 32062 27391 32096
rect 27391 32062 27425 32096
rect 27425 32062 27434 32096
rect 27382 32053 27434 32062
rect 53302 32053 53354 32105
rect 4294 31942 4346 31994
rect 4358 31942 4410 31994
rect 4422 31942 4474 31994
rect 4486 31942 4538 31994
rect 35014 31942 35066 31994
rect 35078 31942 35130 31994
rect 35142 31942 35194 31994
rect 35206 31942 35258 31994
rect 27382 31831 27434 31883
rect 50134 31831 50186 31883
rect 24502 31757 24554 31809
rect 35446 31757 35498 31809
rect 35350 31683 35402 31735
rect 6454 31609 6506 31661
rect 8086 31609 8138 31661
rect 19654 31276 19706 31328
rect 19718 31276 19770 31328
rect 19782 31276 19834 31328
rect 19846 31276 19898 31328
rect 50374 31276 50426 31328
rect 50438 31276 50490 31328
rect 50502 31276 50554 31328
rect 50566 31276 50618 31328
rect 34006 30869 34058 30921
rect 12598 30721 12650 30773
rect 19030 30764 19082 30773
rect 19030 30730 19039 30764
rect 19039 30730 19073 30764
rect 19073 30730 19082 30764
rect 19030 30721 19082 30730
rect 24022 30721 24074 30773
rect 51862 30721 51914 30773
rect 55318 30764 55370 30773
rect 55318 30730 55327 30764
rect 55327 30730 55361 30764
rect 55361 30730 55370 30764
rect 55318 30721 55370 30730
rect 4294 30610 4346 30662
rect 4358 30610 4410 30662
rect 4422 30610 4474 30662
rect 4486 30610 4538 30662
rect 35014 30610 35066 30662
rect 35078 30610 35130 30662
rect 35142 30610 35194 30662
rect 35206 30610 35258 30662
rect 29494 30499 29546 30551
rect 55318 30499 55370 30551
rect 19030 30425 19082 30477
rect 38230 30425 38282 30477
rect 52150 30351 52202 30403
rect 51574 30277 51626 30329
rect 19654 29944 19706 29996
rect 19718 29944 19770 29996
rect 19782 29944 19834 29996
rect 19846 29944 19898 29996
rect 50374 29944 50426 29996
rect 50438 29944 50490 29996
rect 50502 29944 50554 29996
rect 50566 29944 50618 29996
rect 6262 29432 6314 29441
rect 6262 29398 6271 29432
rect 6271 29398 6305 29432
rect 6305 29398 6314 29432
rect 6262 29389 6314 29398
rect 37078 29432 37130 29441
rect 37078 29398 37087 29432
rect 37087 29398 37121 29432
rect 37121 29398 37130 29432
rect 37078 29389 37130 29398
rect 49078 29389 49130 29441
rect 4294 29278 4346 29330
rect 4358 29278 4410 29330
rect 4422 29278 4474 29330
rect 4486 29278 4538 29330
rect 35014 29278 35066 29330
rect 35078 29278 35130 29330
rect 35142 29278 35194 29330
rect 35206 29278 35258 29330
rect 37078 29167 37130 29219
rect 49366 29167 49418 29219
rect 13942 28871 13994 28923
rect 44086 28871 44138 28923
rect 19654 28612 19706 28664
rect 19718 28612 19770 28664
rect 19782 28612 19834 28664
rect 19846 28612 19898 28664
rect 50374 28612 50426 28664
rect 50438 28612 50490 28664
rect 50502 28612 50554 28664
rect 50566 28612 50618 28664
rect 2998 28057 3050 28109
rect 45622 28057 45674 28109
rect 4294 27946 4346 27998
rect 4358 27946 4410 27998
rect 4422 27946 4474 27998
rect 4486 27946 4538 27998
rect 35014 27946 35066 27998
rect 35078 27946 35130 27998
rect 35142 27946 35194 27998
rect 35206 27946 35258 27998
rect 24310 27878 24362 27887
rect 24310 27844 24319 27878
rect 24319 27844 24353 27878
rect 24353 27844 24362 27878
rect 24310 27835 24362 27844
rect 35542 27613 35594 27665
rect 52534 27539 52586 27591
rect 13558 27465 13610 27517
rect 42742 27465 42794 27517
rect 19654 27280 19706 27332
rect 19718 27280 19770 27332
rect 19782 27280 19834 27332
rect 19846 27280 19898 27332
rect 50374 27280 50426 27332
rect 50438 27280 50490 27332
rect 50502 27280 50554 27332
rect 50566 27280 50618 27332
rect 6358 26947 6410 26999
rect 16822 26873 16874 26925
rect 42166 26873 42218 26925
rect 6838 26799 6890 26851
rect 56662 26799 56714 26851
rect 14902 26725 14954 26777
rect 16054 26725 16106 26777
rect 4294 26614 4346 26666
rect 4358 26614 4410 26666
rect 4422 26614 4474 26666
rect 4486 26614 4538 26666
rect 35014 26614 35066 26666
rect 35078 26614 35130 26666
rect 35142 26614 35194 26666
rect 35206 26614 35258 26666
rect 19414 26059 19466 26111
rect 23830 26059 23882 26111
rect 19654 25948 19706 26000
rect 19718 25948 19770 26000
rect 19782 25948 19834 26000
rect 19846 25948 19898 26000
rect 50374 25948 50426 26000
rect 50438 25948 50490 26000
rect 50502 25948 50554 26000
rect 50566 25948 50618 26000
rect 56950 25393 57002 25445
rect 4294 25282 4346 25334
rect 4358 25282 4410 25334
rect 4422 25282 4474 25334
rect 4486 25282 4538 25334
rect 35014 25282 35066 25334
rect 35078 25282 35130 25334
rect 35142 25282 35194 25334
rect 35206 25282 35258 25334
rect 16630 25171 16682 25223
rect 23638 25171 23690 25223
rect 42070 25171 42122 25223
rect 34774 24949 34826 25001
rect 25462 24918 25514 24927
rect 25462 24884 25471 24918
rect 25471 24884 25505 24918
rect 25505 24884 25514 24918
rect 25462 24875 25514 24884
rect 50710 24875 50762 24927
rect 32470 24801 32522 24853
rect 19654 24616 19706 24668
rect 19718 24616 19770 24668
rect 19782 24616 19834 24668
rect 19846 24616 19898 24668
rect 50374 24616 50426 24668
rect 50438 24616 50490 24668
rect 50502 24616 50554 24668
rect 50566 24616 50618 24668
rect 3574 24283 3626 24335
rect 23254 24283 23306 24335
rect 15286 24209 15338 24261
rect 39094 24209 39146 24261
rect 7126 24135 7178 24187
rect 31414 24135 31466 24187
rect 21430 24061 21482 24113
rect 4294 23950 4346 24002
rect 4358 23950 4410 24002
rect 4422 23950 4474 24002
rect 4486 23950 4538 24002
rect 35014 23950 35066 24002
rect 35078 23950 35130 24002
rect 35142 23950 35194 24002
rect 35206 23950 35258 24002
rect 17398 23839 17450 23891
rect 41878 23839 41930 23891
rect 15958 23765 16010 23817
rect 45430 23765 45482 23817
rect 3670 23691 3722 23743
rect 53206 23691 53258 23743
rect 19654 23284 19706 23336
rect 19718 23284 19770 23336
rect 19782 23284 19834 23336
rect 19846 23284 19898 23336
rect 50374 23284 50426 23336
rect 50438 23284 50490 23336
rect 50502 23284 50554 23336
rect 50566 23284 50618 23336
rect 8566 22877 8618 22929
rect 39574 22877 39626 22929
rect 1942 22803 1994 22855
rect 13558 22772 13610 22781
rect 13558 22738 13567 22772
rect 13567 22738 13601 22772
rect 13601 22738 13610 22772
rect 13558 22729 13610 22738
rect 17782 22772 17834 22781
rect 17782 22738 17791 22772
rect 17791 22738 17825 22772
rect 17825 22738 17834 22772
rect 17782 22729 17834 22738
rect 26902 22772 26954 22781
rect 26902 22738 26911 22772
rect 26911 22738 26945 22772
rect 26945 22738 26954 22772
rect 26902 22729 26954 22738
rect 30934 22772 30986 22781
rect 30934 22738 30943 22772
rect 30943 22738 30977 22772
rect 30977 22738 30986 22772
rect 30934 22729 30986 22738
rect 51094 22803 51146 22855
rect 4294 22618 4346 22670
rect 4358 22618 4410 22670
rect 4422 22618 4474 22670
rect 4486 22618 4538 22670
rect 35014 22618 35066 22670
rect 35078 22618 35130 22670
rect 35142 22618 35194 22670
rect 35206 22618 35258 22670
rect 8854 22507 8906 22559
rect 13558 22507 13610 22559
rect 32758 22507 32810 22559
rect 8566 22433 8618 22485
rect 36886 22433 36938 22485
rect 16534 22359 16586 22411
rect 40246 22359 40298 22411
rect 19510 22285 19562 22337
rect 20950 22285 21002 22337
rect 35638 22137 35690 22189
rect 8758 22063 8810 22115
rect 19654 21952 19706 22004
rect 19718 21952 19770 22004
rect 19782 21952 19834 22004
rect 19846 21952 19898 22004
rect 50374 21952 50426 22004
rect 50438 21952 50490 22004
rect 50502 21952 50554 22004
rect 50566 21952 50618 22004
rect 3574 21841 3626 21893
rect 26902 21841 26954 21893
rect 8758 21545 8810 21597
rect 58102 21545 58154 21597
rect 8374 21471 8426 21523
rect 55510 21471 55562 21523
rect 7990 21397 8042 21449
rect 53878 21397 53930 21449
rect 4294 21286 4346 21338
rect 4358 21286 4410 21338
rect 4422 21286 4474 21338
rect 4486 21286 4538 21338
rect 35014 21286 35066 21338
rect 35078 21286 35130 21338
rect 35142 21286 35194 21338
rect 35206 21286 35258 21338
rect 8758 21101 8810 21153
rect 8374 21027 8426 21079
rect 7942 20953 7994 21005
rect 21622 20879 21674 20931
rect 44662 20731 44714 20783
rect 19654 20620 19706 20672
rect 19718 20620 19770 20672
rect 19782 20620 19834 20672
rect 19846 20620 19898 20672
rect 50374 20620 50426 20672
rect 50438 20620 50490 20672
rect 50502 20620 50554 20672
rect 50566 20620 50618 20672
rect 20854 20509 20906 20561
rect 10870 20287 10922 20339
rect 17974 20287 18026 20339
rect 21526 20065 21578 20117
rect 43894 20065 43946 20117
rect 49654 20108 49706 20117
rect 49654 20074 49663 20108
rect 49663 20074 49697 20108
rect 49697 20074 49706 20108
rect 49654 20065 49706 20074
rect 4294 19954 4346 20006
rect 4358 19954 4410 20006
rect 4422 19954 4474 20006
rect 4486 19954 4538 20006
rect 35014 19954 35066 20006
rect 35078 19954 35130 20006
rect 35142 19954 35194 20006
rect 35206 19954 35258 20006
rect 8278 19769 8330 19821
rect 53974 19843 54026 19895
rect 38230 19769 38282 19821
rect 45046 19769 45098 19821
rect 17782 19695 17834 19747
rect 43990 19695 44042 19747
rect 45814 19621 45866 19673
rect 10966 19547 11018 19599
rect 7942 19473 7994 19525
rect 20854 19399 20906 19451
rect 19654 19288 19706 19340
rect 19718 19288 19770 19340
rect 19782 19288 19834 19340
rect 19846 19288 19898 19340
rect 50374 19288 50426 19340
rect 50438 19288 50490 19340
rect 50502 19288 50554 19340
rect 50566 19288 50618 19340
rect 7990 19177 8042 19229
rect 48694 19177 48746 19229
rect 8278 19029 8330 19081
rect 50806 19029 50858 19081
rect 8662 18955 8714 19007
rect 13462 18955 13514 19007
rect 25942 18807 25994 18859
rect 27862 18807 27914 18859
rect 34678 18733 34730 18785
rect 54646 18733 54698 18785
rect 4294 18622 4346 18674
rect 4358 18622 4410 18674
rect 4422 18622 4474 18674
rect 4486 18622 4538 18674
rect 35014 18622 35066 18674
rect 35078 18622 35130 18674
rect 35142 18622 35194 18674
rect 35206 18622 35258 18674
rect 8182 18437 8234 18489
rect 48598 18437 48650 18489
rect 17302 18215 17354 18267
rect 30838 18258 30890 18267
rect 30838 18224 30847 18258
rect 30847 18224 30881 18258
rect 30881 18224 30890 18258
rect 30838 18215 30890 18224
rect 42838 18258 42890 18267
rect 42838 18224 42847 18258
rect 42847 18224 42881 18258
rect 42881 18224 42890 18258
rect 42838 18215 42890 18224
rect 7942 18141 7994 18193
rect 8374 18141 8426 18193
rect 12022 18141 12074 18193
rect 8182 18067 8234 18119
rect 45814 18110 45866 18119
rect 45814 18076 45823 18110
rect 45823 18076 45857 18110
rect 45857 18076 45866 18110
rect 45814 18067 45866 18076
rect 19654 17956 19706 18008
rect 19718 17956 19770 18008
rect 19782 17956 19834 18008
rect 19846 17956 19898 18008
rect 50374 17956 50426 18008
rect 50438 17956 50490 18008
rect 50502 17956 50554 18008
rect 50566 17956 50618 18008
rect 12022 17771 12074 17823
rect 42934 17771 42986 17823
rect 8374 17697 8426 17749
rect 44758 17697 44810 17749
rect 7990 17623 8042 17675
rect 46102 17623 46154 17675
rect 5206 17549 5258 17601
rect 8566 17475 8618 17527
rect 45814 17475 45866 17527
rect 12406 17401 12458 17453
rect 4294 17290 4346 17342
rect 4358 17290 4410 17342
rect 4422 17290 4474 17342
rect 4486 17290 4538 17342
rect 35014 17290 35066 17342
rect 35078 17290 35130 17342
rect 35142 17290 35194 17342
rect 35206 17290 35258 17342
rect 42646 17105 42698 17157
rect 21526 17031 21578 17083
rect 48598 17031 48650 17083
rect 11062 16957 11114 17009
rect 21526 16883 21578 16935
rect 12022 16809 12074 16861
rect 8182 16735 8234 16787
rect 19654 16624 19706 16676
rect 19718 16624 19770 16676
rect 19782 16624 19834 16676
rect 19846 16624 19898 16676
rect 50374 16624 50426 16676
rect 50438 16624 50490 16676
rect 50502 16624 50554 16676
rect 50566 16624 50618 16676
rect 10006 16513 10058 16565
rect 42838 16513 42890 16565
rect 12022 16439 12074 16491
rect 37942 16439 37994 16491
rect 8182 16365 8234 16417
rect 39766 16365 39818 16417
rect 57334 16143 57386 16195
rect 8278 16069 8330 16121
rect 13942 16069 13994 16121
rect 49558 16112 49610 16121
rect 49558 16078 49567 16112
rect 49567 16078 49601 16112
rect 49601 16078 49610 16112
rect 49558 16069 49610 16078
rect 4294 15958 4346 16010
rect 4358 15958 4410 16010
rect 4422 15958 4474 16010
rect 4486 15958 4538 16010
rect 35014 15958 35066 16010
rect 35078 15958 35130 16010
rect 35142 15958 35194 16010
rect 35206 15958 35258 16010
rect 16630 15847 16682 15899
rect 20086 15847 20138 15899
rect 27766 15847 27818 15899
rect 35734 15847 35786 15899
rect 49558 15847 49610 15899
rect 37462 15773 37514 15825
rect 8374 15551 8426 15603
rect 34102 15477 34154 15529
rect 8758 15403 8810 15455
rect 12982 15403 13034 15455
rect 34870 15403 34922 15455
rect 19654 15292 19706 15344
rect 19718 15292 19770 15344
rect 19782 15292 19834 15344
rect 19846 15292 19898 15344
rect 50374 15292 50426 15344
rect 50438 15292 50490 15344
rect 50502 15292 50554 15344
rect 50566 15292 50618 15344
rect 8758 15181 8810 15233
rect 12982 15181 13034 15233
rect 39862 15181 39914 15233
rect 8374 15107 8426 15159
rect 31894 15107 31946 15159
rect 7318 14811 7370 14863
rect 36598 14811 36650 14863
rect 4054 14737 4106 14789
rect 20470 14780 20522 14789
rect 20470 14746 20479 14780
rect 20479 14746 20513 14780
rect 20513 14746 20522 14780
rect 20470 14737 20522 14746
rect 21238 14737 21290 14789
rect 54454 14737 54506 14789
rect 4294 14626 4346 14678
rect 4358 14626 4410 14678
rect 4422 14626 4474 14678
rect 4486 14626 4538 14678
rect 35014 14626 35066 14678
rect 35078 14626 35130 14678
rect 35142 14626 35194 14678
rect 35206 14626 35258 14678
rect 36598 14558 36650 14567
rect 8182 14441 8234 14493
rect 36598 14524 36607 14558
rect 36607 14524 36641 14558
rect 36641 14524 36650 14558
rect 36598 14515 36650 14524
rect 31318 14441 31370 14493
rect 7606 14410 7658 14419
rect 7606 14376 7615 14410
rect 7615 14376 7649 14410
rect 7649 14376 7658 14410
rect 7606 14367 7658 14376
rect 8182 14145 8234 14197
rect 30838 14145 30890 14197
rect 42838 14145 42890 14197
rect 34390 14071 34442 14123
rect 46678 14071 46730 14123
rect 19654 13960 19706 14012
rect 19718 13960 19770 14012
rect 19782 13960 19834 14012
rect 19846 13960 19898 14012
rect 50374 13960 50426 14012
rect 50438 13960 50490 14012
rect 50502 13960 50554 14012
rect 50566 13960 50618 14012
rect 27574 13849 27626 13901
rect 40918 13849 40970 13901
rect 8182 13775 8234 13827
rect 28822 13775 28874 13827
rect 37750 13775 37802 13827
rect 51862 13775 51914 13827
rect 33814 13701 33866 13753
rect 56950 13701 57002 13753
rect 26038 13627 26090 13679
rect 57046 13627 57098 13679
rect 9910 13405 9962 13457
rect 11446 13448 11498 13457
rect 11446 13414 11455 13448
rect 11455 13414 11489 13448
rect 11489 13414 11498 13448
rect 11446 13405 11498 13414
rect 29590 13479 29642 13531
rect 57718 13405 57770 13457
rect 4294 13294 4346 13346
rect 4358 13294 4410 13346
rect 4422 13294 4474 13346
rect 4486 13294 4538 13346
rect 35014 13294 35066 13346
rect 35078 13294 35130 13346
rect 35142 13294 35194 13346
rect 35206 13294 35258 13346
rect 9910 13183 9962 13235
rect 43702 13183 43754 13235
rect 28150 13109 28202 13161
rect 29014 13109 29066 13161
rect 32662 13109 32714 13161
rect 8566 13035 8618 13087
rect 13750 13035 13802 13087
rect 12886 12961 12938 13013
rect 30166 12961 30218 13013
rect 26326 12813 26378 12865
rect 19654 12628 19706 12680
rect 19718 12628 19770 12680
rect 19782 12628 19834 12680
rect 19846 12628 19898 12680
rect 50374 12628 50426 12680
rect 50438 12628 50490 12680
rect 50502 12628 50554 12680
rect 50566 12628 50618 12680
rect 20278 12517 20330 12569
rect 20854 12517 20906 12569
rect 57238 12517 57290 12569
rect 20662 12369 20714 12421
rect 20854 12369 20906 12421
rect 51094 12369 51146 12421
rect 52822 12369 52874 12421
rect 2326 12295 2378 12347
rect 44182 12295 44234 12347
rect 7798 12147 7850 12199
rect 24982 12147 25034 12199
rect 57526 12147 57578 12199
rect 20374 12116 20426 12125
rect 20374 12082 20383 12116
rect 20383 12082 20417 12116
rect 20417 12082 20426 12116
rect 20374 12073 20426 12082
rect 31030 12116 31082 12125
rect 31030 12082 31039 12116
rect 31039 12082 31073 12116
rect 31073 12082 31082 12116
rect 31030 12073 31082 12082
rect 41782 12073 41834 12125
rect 44758 12073 44810 12125
rect 45334 12073 45386 12125
rect 4294 11962 4346 12014
rect 4358 11962 4410 12014
rect 4422 11962 4474 12014
rect 4486 11962 4538 12014
rect 35014 11962 35066 12014
rect 35078 11962 35130 12014
rect 35142 11962 35194 12014
rect 35206 11962 35258 12014
rect 2326 11894 2378 11903
rect 2326 11860 2335 11894
rect 2335 11860 2369 11894
rect 2369 11860 2378 11894
rect 2326 11851 2378 11860
rect 2710 11851 2762 11903
rect 7798 11777 7850 11829
rect 20374 11777 20426 11829
rect 50806 11777 50858 11829
rect 2518 11629 2570 11681
rect 3574 11629 3626 11681
rect 2998 11598 3050 11607
rect 2998 11564 3007 11598
rect 3007 11564 3041 11598
rect 3041 11564 3050 11598
rect 2998 11555 3050 11564
rect 24502 11703 24554 11755
rect 31030 11703 31082 11755
rect 27958 11629 28010 11681
rect 44758 11703 44810 11755
rect 44854 11703 44906 11755
rect 23350 11555 23402 11607
rect 31510 11555 31562 11607
rect 36502 11555 36554 11607
rect 52630 11629 52682 11681
rect 20854 11481 20906 11533
rect 24118 11481 24170 11533
rect 59734 11555 59786 11607
rect 56278 11407 56330 11459
rect 19654 11296 19706 11348
rect 19718 11296 19770 11348
rect 19782 11296 19834 11348
rect 19846 11296 19898 11348
rect 50374 11296 50426 11348
rect 50438 11296 50490 11348
rect 50502 11296 50554 11348
rect 50566 11296 50618 11348
rect 54646 11037 54698 11089
rect 17014 10963 17066 11015
rect 30166 10963 30218 11015
rect 57910 11037 57962 11089
rect 21526 10889 21578 10941
rect 34582 10889 34634 10941
rect 2998 10815 3050 10867
rect 41206 10815 41258 10867
rect 48790 10815 48842 10867
rect 56758 10889 56810 10941
rect 56854 10815 56906 10867
rect 40438 10741 40490 10793
rect 44758 10784 44810 10793
rect 44758 10750 44767 10784
rect 44767 10750 44801 10784
rect 44801 10750 44810 10784
rect 44758 10741 44810 10750
rect 51862 10741 51914 10793
rect 4294 10630 4346 10682
rect 4358 10630 4410 10682
rect 4422 10630 4474 10682
rect 4486 10630 4538 10682
rect 35014 10630 35066 10682
rect 35078 10630 35130 10682
rect 35142 10630 35194 10682
rect 35206 10630 35258 10682
rect 11446 10445 11498 10497
rect 12310 10371 12362 10423
rect 55030 10414 55082 10423
rect 55030 10380 55039 10414
rect 55039 10380 55073 10414
rect 55073 10380 55082 10414
rect 55030 10371 55082 10380
rect 58582 10519 58634 10571
rect 22390 10297 22442 10349
rect 17590 10223 17642 10275
rect 48694 10223 48746 10275
rect 56470 10149 56522 10201
rect 22102 10075 22154 10127
rect 35542 10075 35594 10127
rect 36118 10075 36170 10127
rect 55702 10075 55754 10127
rect 56086 10075 56138 10127
rect 19654 9964 19706 10016
rect 19718 9964 19770 10016
rect 19782 9964 19834 10016
rect 19846 9964 19898 10016
rect 50374 9964 50426 10016
rect 50438 9964 50490 10016
rect 50502 9964 50554 10016
rect 50566 9964 50618 10016
rect 22966 9853 23018 9905
rect 24022 9853 24074 9905
rect 32374 9853 32426 9905
rect 33142 9853 33194 9905
rect 35638 9853 35690 9905
rect 36214 9853 36266 9905
rect 54070 9853 54122 9905
rect 6070 9779 6122 9831
rect 15862 9779 15914 9831
rect 21910 9779 21962 9831
rect 25174 9779 25226 9831
rect 32758 9779 32810 9831
rect 34006 9779 34058 9831
rect 35446 9779 35498 9831
rect 36982 9779 37034 9831
rect 6262 9705 6314 9757
rect 14710 9705 14762 9757
rect 19222 9705 19274 9757
rect 23734 9705 23786 9757
rect 34294 9705 34346 9757
rect 35734 9705 35786 9757
rect 36790 9705 36842 9757
rect 54454 9748 54506 9757
rect 5686 9631 5738 9683
rect 13846 9631 13898 9683
rect 13942 9631 13994 9683
rect 24502 9631 24554 9683
rect 10678 9557 10730 9609
rect 24310 9557 24362 9609
rect 30358 9557 30410 9609
rect 38422 9557 38474 9609
rect 54454 9714 54463 9748
rect 54463 9714 54497 9748
rect 54497 9714 54506 9748
rect 54454 9705 54506 9714
rect 57814 9779 57866 9831
rect 49654 9631 49706 9683
rect 17686 9483 17738 9535
rect 32566 9483 32618 9535
rect 50230 9483 50282 9535
rect 8278 9409 8330 9461
rect 16150 9409 16202 9461
rect 16246 9409 16298 9461
rect 20278 9409 20330 9461
rect 50998 9409 51050 9461
rect 53782 9452 53834 9461
rect 53782 9418 53791 9452
rect 53791 9418 53825 9452
rect 53825 9418 53834 9452
rect 53782 9409 53834 9418
rect 54262 9557 54314 9609
rect 54934 9483 54986 9535
rect 55318 9557 55370 9609
rect 57622 9674 57674 9683
rect 57622 9640 57631 9674
rect 57631 9640 57665 9674
rect 57665 9640 57674 9674
rect 57622 9631 57674 9640
rect 4294 9298 4346 9350
rect 4358 9298 4410 9350
rect 4422 9298 4474 9350
rect 4486 9298 4538 9350
rect 35014 9298 35066 9350
rect 35078 9298 35130 9350
rect 35142 9298 35194 9350
rect 35206 9298 35258 9350
rect 12502 9113 12554 9165
rect 7942 8891 7994 8943
rect 21526 9187 21578 9239
rect 53782 9187 53834 9239
rect 30934 9113 30986 9165
rect 23926 9039 23978 9091
rect 29686 9039 29738 9091
rect 30358 9082 30410 9091
rect 30358 9048 30367 9082
rect 30367 9048 30401 9082
rect 30401 9048 30410 9082
rect 30358 9039 30410 9048
rect 36790 9082 36842 9091
rect 36790 9048 36799 9082
rect 36799 9048 36833 9082
rect 36833 9048 36842 9082
rect 36790 9039 36842 9048
rect 48694 9113 48746 9165
rect 15190 8965 15242 9017
rect 55894 8965 55946 9017
rect 57238 9008 57290 9017
rect 43030 8891 43082 8943
rect 53206 8891 53258 8943
rect 57238 8974 57247 9008
rect 57247 8974 57281 9008
rect 57281 8974 57290 9008
rect 57238 8965 57290 8974
rect 12598 8817 12650 8869
rect 10198 8743 10250 8795
rect 14902 8743 14954 8795
rect 35062 8817 35114 8869
rect 57334 8891 57386 8943
rect 18838 8743 18890 8795
rect 44950 8743 45002 8795
rect 53878 8743 53930 8795
rect 54646 8743 54698 8795
rect 19654 8632 19706 8684
rect 19718 8632 19770 8684
rect 19782 8632 19834 8684
rect 19846 8632 19898 8684
rect 50374 8632 50426 8684
rect 50438 8632 50490 8684
rect 50502 8632 50554 8684
rect 50566 8632 50618 8684
rect 3670 8521 3722 8573
rect 5590 8521 5642 8573
rect 12790 8521 12842 8573
rect 3286 8416 3338 8425
rect 3286 8382 3295 8416
rect 3295 8382 3329 8416
rect 3329 8382 3338 8416
rect 3286 8373 3338 8382
rect 7222 8299 7274 8351
rect 9430 8299 9482 8351
rect 42166 8521 42218 8573
rect 48598 8564 48650 8573
rect 48598 8530 48607 8564
rect 48607 8530 48641 8564
rect 48641 8530 48650 8564
rect 48598 8521 48650 8530
rect 58966 8521 59018 8573
rect 10582 8416 10634 8425
rect 10582 8382 10591 8416
rect 10591 8382 10625 8416
rect 10625 8382 10634 8416
rect 10582 8373 10634 8382
rect 11350 8416 11402 8425
rect 11350 8382 11359 8416
rect 11359 8382 11393 8416
rect 11393 8382 11402 8416
rect 11350 8373 11402 8382
rect 12118 8416 12170 8425
rect 12118 8382 12127 8416
rect 12127 8382 12161 8416
rect 12161 8382 12170 8416
rect 12118 8373 12170 8382
rect 12886 8416 12938 8425
rect 12886 8382 12895 8416
rect 12895 8382 12929 8416
rect 12929 8382 12938 8416
rect 12886 8373 12938 8382
rect 13654 8416 13706 8425
rect 13654 8382 13663 8416
rect 13663 8382 13697 8416
rect 13697 8382 13706 8416
rect 13654 8373 13706 8382
rect 33910 8373 33962 8425
rect 34390 8416 34442 8425
rect 34390 8382 34399 8416
rect 34399 8382 34433 8416
rect 34433 8382 34442 8416
rect 34390 8373 34442 8382
rect 35062 8416 35114 8425
rect 35062 8382 35071 8416
rect 35071 8382 35105 8416
rect 35105 8382 35114 8416
rect 35062 8373 35114 8382
rect 44374 8447 44426 8499
rect 42166 8416 42218 8425
rect 42166 8382 42175 8416
rect 42175 8382 42209 8416
rect 42209 8382 42218 8416
rect 42166 8373 42218 8382
rect 16246 8342 16298 8351
rect 16246 8308 16255 8342
rect 16255 8308 16289 8342
rect 16289 8308 16298 8342
rect 16246 8299 16298 8308
rect 17014 8342 17066 8351
rect 17014 8308 17023 8342
rect 17023 8308 17057 8342
rect 17057 8308 17066 8342
rect 17014 8299 17066 8308
rect 17110 8299 17162 8351
rect 50710 8447 50762 8499
rect 48886 8373 48938 8425
rect 52534 8416 52586 8425
rect 52534 8382 52543 8416
rect 52543 8382 52577 8416
rect 52577 8382 52586 8416
rect 52534 8373 52586 8382
rect 53302 8416 53354 8425
rect 53302 8382 53311 8416
rect 53311 8382 53345 8416
rect 53345 8382 53354 8416
rect 53302 8373 53354 8382
rect 48790 8299 48842 8351
rect 52918 8299 52970 8351
rect 59830 8373 59882 8425
rect 1654 8268 1706 8277
rect 1654 8234 1663 8268
rect 1663 8234 1697 8268
rect 1697 8234 1706 8268
rect 1654 8225 1706 8234
rect 2134 8225 2186 8277
rect 2710 8225 2762 8277
rect 2998 8225 3050 8277
rect 7702 8225 7754 8277
rect 4822 8151 4874 8203
rect 9622 8225 9674 8277
rect 9718 8268 9770 8277
rect 9718 8234 9743 8268
rect 9743 8234 9770 8268
rect 9718 8225 9770 8234
rect 9910 8225 9962 8277
rect 9814 8151 9866 8203
rect 10294 8225 10346 8277
rect 10582 8225 10634 8277
rect 11350 8225 11402 8277
rect 12118 8225 12170 8277
rect 16150 8268 16202 8277
rect 16150 8234 16159 8268
rect 16159 8234 16193 8268
rect 16193 8234 16202 8268
rect 16150 8225 16202 8234
rect 16342 8225 16394 8277
rect 48022 8225 48074 8277
rect 48598 8225 48650 8277
rect 48694 8151 48746 8203
rect 49462 8225 49514 8277
rect 53110 8225 53162 8277
rect 53494 8225 53546 8277
rect 56950 8299 57002 8351
rect 58390 8225 58442 8277
rect 51190 8151 51242 8203
rect 56662 8151 56714 8203
rect 6166 8120 6218 8129
rect 6166 8086 6175 8120
rect 6175 8086 6209 8120
rect 6209 8086 6218 8120
rect 6166 8077 6218 8086
rect 7606 8077 7658 8129
rect 7798 8077 7850 8129
rect 8566 8077 8618 8129
rect 9622 8077 9674 8129
rect 17782 8120 17834 8129
rect 17782 8086 17791 8120
rect 17791 8086 17825 8120
rect 17825 8086 17834 8120
rect 17782 8077 17834 8086
rect 22102 8120 22154 8129
rect 22102 8086 22111 8120
rect 22111 8086 22145 8120
rect 22145 8086 22154 8120
rect 22102 8077 22154 8086
rect 28054 8077 28106 8129
rect 52534 8077 52586 8129
rect 57718 8077 57770 8129
rect 4294 7966 4346 8018
rect 4358 7966 4410 8018
rect 4422 7966 4474 8018
rect 4486 7966 4538 8018
rect 35014 7966 35066 8018
rect 35078 7966 35130 8018
rect 35142 7966 35194 8018
rect 35206 7966 35258 8018
rect 2902 7898 2954 7907
rect 2902 7864 2911 7898
rect 2911 7864 2945 7898
rect 2945 7864 2954 7898
rect 2902 7855 2954 7864
rect 2518 7750 2570 7759
rect 2518 7716 2527 7750
rect 2527 7716 2561 7750
rect 2561 7716 2570 7750
rect 2518 7707 2570 7716
rect 8566 7855 8618 7907
rect 7798 7781 7850 7833
rect 11254 7781 11306 7833
rect 22102 7855 22154 7907
rect 17110 7781 17162 7833
rect 24310 7824 24362 7833
rect 24310 7790 24319 7824
rect 24319 7790 24353 7824
rect 24353 7790 24362 7824
rect 25078 7824 25130 7833
rect 24310 7781 24362 7790
rect 4054 7750 4106 7759
rect 4054 7716 4063 7750
rect 4063 7716 4097 7750
rect 4097 7716 4106 7750
rect 4054 7707 4106 7716
rect 4918 7707 4970 7759
rect 5590 7750 5642 7759
rect 5590 7716 5599 7750
rect 5599 7716 5633 7750
rect 5633 7716 5642 7750
rect 5590 7707 5642 7716
rect 7942 7707 7994 7759
rect 10198 7750 10250 7759
rect 1462 7633 1514 7685
rect 10198 7716 10207 7750
rect 10207 7716 10241 7750
rect 10241 7716 10250 7750
rect 10198 7707 10250 7716
rect 10966 7750 11018 7759
rect 10966 7716 10975 7750
rect 10975 7716 11009 7750
rect 11009 7716 11018 7750
rect 10966 7707 11018 7716
rect 12406 7750 12458 7759
rect 12406 7716 12415 7750
rect 12415 7716 12449 7750
rect 12449 7716 12458 7750
rect 12406 7707 12458 7716
rect 12502 7707 12554 7759
rect 15958 7707 16010 7759
rect 20950 7750 21002 7759
rect 20950 7716 20959 7750
rect 20959 7716 20993 7750
rect 20993 7716 21002 7750
rect 20950 7707 21002 7716
rect 23926 7750 23978 7759
rect 23926 7716 23935 7750
rect 23935 7716 23969 7750
rect 23969 7716 23978 7750
rect 23926 7707 23978 7716
rect 25078 7790 25087 7824
rect 25087 7790 25121 7824
rect 25121 7790 25130 7824
rect 28918 7855 28970 7907
rect 36502 7898 36554 7907
rect 36502 7864 36511 7898
rect 36511 7864 36545 7898
rect 36545 7864 36554 7898
rect 36502 7855 36554 7864
rect 39094 7855 39146 7907
rect 40246 7855 40298 7907
rect 25078 7781 25130 7790
rect 24790 7707 24842 7759
rect 37462 7781 37514 7833
rect 44758 7855 44810 7907
rect 26134 7750 26186 7759
rect 26134 7716 26143 7750
rect 26143 7716 26177 7750
rect 26177 7716 26186 7750
rect 26134 7707 26186 7716
rect 28918 7707 28970 7759
rect 30166 7750 30218 7759
rect 30166 7716 30175 7750
rect 30175 7716 30209 7750
rect 30209 7716 30218 7750
rect 30166 7707 30218 7716
rect 33814 7750 33866 7759
rect 33814 7716 33823 7750
rect 33823 7716 33857 7750
rect 33857 7716 33866 7750
rect 33814 7707 33866 7716
rect 34582 7750 34634 7759
rect 34582 7716 34591 7750
rect 34591 7716 34625 7750
rect 34625 7716 34634 7750
rect 34582 7707 34634 7716
rect 35350 7750 35402 7759
rect 35350 7716 35359 7750
rect 35359 7716 35393 7750
rect 35393 7716 35402 7750
rect 35350 7707 35402 7716
rect 36118 7750 36170 7759
rect 36118 7716 36127 7750
rect 36127 7716 36161 7750
rect 36161 7716 36170 7750
rect 36118 7707 36170 7716
rect 36502 7707 36554 7759
rect 9430 7676 9482 7685
rect 9430 7642 9439 7676
rect 9439 7642 9473 7676
rect 9473 7642 9482 7676
rect 9430 7633 9482 7642
rect 7030 7559 7082 7611
rect 8230 7559 8282 7611
rect 14230 7559 14282 7611
rect 9142 7485 9194 7537
rect 11734 7485 11786 7537
rect 15958 7559 16010 7611
rect 2422 7454 2474 7463
rect 2422 7420 2431 7454
rect 2431 7420 2465 7454
rect 2465 7420 2474 7454
rect 2422 7411 2474 7420
rect 3286 7411 3338 7463
rect 3382 7411 3434 7463
rect 4054 7411 4106 7463
rect 5302 7411 5354 7463
rect 8758 7411 8810 7463
rect 9910 7411 9962 7463
rect 10966 7411 11018 7463
rect 23158 7485 23210 7537
rect 25462 7559 25514 7611
rect 38806 7707 38858 7759
rect 40246 7707 40298 7759
rect 41782 7707 41834 7759
rect 42742 7707 42794 7759
rect 43990 7707 44042 7759
rect 45046 7707 45098 7759
rect 45622 7750 45674 7759
rect 45622 7716 45631 7750
rect 45631 7716 45665 7750
rect 45665 7716 45674 7750
rect 45622 7707 45674 7716
rect 45814 7707 45866 7759
rect 51190 7855 51242 7907
rect 51478 7898 51530 7907
rect 51478 7864 51487 7898
rect 51487 7864 51521 7898
rect 51521 7864 51530 7898
rect 51478 7855 51530 7864
rect 46486 7707 46538 7759
rect 39094 7633 39146 7685
rect 30166 7485 30218 7537
rect 30646 7559 30698 7611
rect 32374 7602 32426 7611
rect 32374 7568 32383 7602
rect 32383 7568 32417 7602
rect 32417 7568 32426 7602
rect 32374 7559 32426 7568
rect 43894 7633 43946 7685
rect 51670 7781 51722 7833
rect 49366 7750 49418 7759
rect 49366 7716 49375 7750
rect 49375 7716 49409 7750
rect 49409 7716 49418 7750
rect 49366 7707 49418 7716
rect 50998 7707 51050 7759
rect 52630 7750 52682 7759
rect 52630 7716 52639 7750
rect 52639 7716 52673 7750
rect 52673 7716 52682 7750
rect 52630 7707 52682 7716
rect 53398 7750 53450 7759
rect 53398 7716 53407 7750
rect 53407 7716 53441 7750
rect 53441 7716 53450 7750
rect 53398 7707 53450 7716
rect 40150 7559 40202 7611
rect 52534 7633 52586 7685
rect 58774 7707 58826 7759
rect 55798 7676 55850 7685
rect 55798 7642 55807 7676
rect 55807 7642 55841 7676
rect 55841 7642 55850 7676
rect 55798 7633 55850 7642
rect 56182 7633 56234 7685
rect 56662 7633 56714 7685
rect 47926 7602 47978 7611
rect 47926 7568 47935 7602
rect 47935 7568 47969 7602
rect 47969 7568 47978 7602
rect 47926 7559 47978 7568
rect 57142 7559 57194 7611
rect 48118 7485 48170 7537
rect 49174 7485 49226 7537
rect 15670 7411 15722 7463
rect 20758 7411 20810 7463
rect 23734 7411 23786 7463
rect 24694 7454 24746 7463
rect 24694 7420 24703 7454
rect 24703 7420 24737 7454
rect 24737 7420 24746 7454
rect 24694 7411 24746 7420
rect 25942 7411 25994 7463
rect 26710 7411 26762 7463
rect 28150 7411 28202 7463
rect 29206 7411 29258 7463
rect 29590 7411 29642 7463
rect 31030 7411 31082 7463
rect 33622 7411 33674 7463
rect 34390 7411 34442 7463
rect 34774 7411 34826 7463
rect 35830 7411 35882 7463
rect 36598 7411 36650 7463
rect 38038 7411 38090 7463
rect 39478 7411 39530 7463
rect 41782 7454 41834 7463
rect 41782 7420 41791 7454
rect 41791 7420 41825 7454
rect 41825 7420 41834 7454
rect 41782 7411 41834 7420
rect 42454 7411 42506 7463
rect 43894 7411 43946 7463
rect 44758 7454 44810 7463
rect 44758 7420 44767 7454
rect 44767 7420 44801 7454
rect 44801 7420 44810 7454
rect 44758 7411 44810 7420
rect 45046 7411 45098 7463
rect 47254 7411 47306 7463
rect 48406 7411 48458 7463
rect 59350 7485 59402 7537
rect 51670 7411 51722 7463
rect 52342 7411 52394 7463
rect 52726 7411 52778 7463
rect 19654 7300 19706 7352
rect 19718 7300 19770 7352
rect 19782 7300 19834 7352
rect 19846 7300 19898 7352
rect 50374 7300 50426 7352
rect 50438 7300 50490 7352
rect 50502 7300 50554 7352
rect 50566 7300 50618 7352
rect 1846 7189 1898 7241
rect 7798 7189 7850 7241
rect 32374 7189 32426 7241
rect 47926 7189 47978 7241
rect 6838 7084 6890 7093
rect 6838 7050 6847 7084
rect 6847 7050 6881 7084
rect 6881 7050 6890 7084
rect 6838 7041 6890 7050
rect 7606 7084 7658 7093
rect 7606 7050 7615 7084
rect 7615 7050 7649 7084
rect 7649 7050 7658 7084
rect 7606 7041 7658 7050
rect 8374 7084 8426 7093
rect 8374 7050 8383 7084
rect 8383 7050 8417 7084
rect 8417 7050 8426 7084
rect 8374 7041 8426 7050
rect 10006 7041 10058 7093
rect 10870 7041 10922 7093
rect 13462 7041 13514 7093
rect 14998 7084 15050 7093
rect 14998 7050 15007 7084
rect 15007 7050 15041 7084
rect 15041 7050 15050 7084
rect 14998 7041 15050 7050
rect 16054 7041 16106 7093
rect 16630 7084 16682 7093
rect 16630 7050 16639 7084
rect 16639 7050 16673 7084
rect 16673 7050 16682 7084
rect 16630 7041 16682 7050
rect 17302 7084 17354 7093
rect 17302 7050 17311 7084
rect 17311 7050 17345 7084
rect 17345 7050 17354 7084
rect 17302 7041 17354 7050
rect 1654 7010 1706 7019
rect 1654 6976 1663 7010
rect 1663 6976 1697 7010
rect 1697 6976 1706 7010
rect 1654 6967 1706 6976
rect 2518 7010 2570 7019
rect 2518 6976 2527 7010
rect 2527 6976 2561 7010
rect 2561 6976 2570 7010
rect 2518 6967 2570 6976
rect 3670 6967 3722 7019
rect 11254 7010 11306 7019
rect 5782 6893 5834 6945
rect 5878 6893 5930 6945
rect 6550 6893 6602 6945
rect 6934 6893 6986 6945
rect 7318 6819 7370 6871
rect 5206 6745 5258 6797
rect 8182 6745 8234 6797
rect 9814 6893 9866 6945
rect 11254 6976 11263 7010
rect 11263 6976 11297 7010
rect 11297 6976 11306 7010
rect 11254 6967 11306 6976
rect 12694 7010 12746 7019
rect 12694 6976 12703 7010
rect 12703 6976 12737 7010
rect 12737 6976 12746 7010
rect 12694 6967 12746 6976
rect 15958 6967 16010 7019
rect 17878 7115 17930 7167
rect 19990 7158 20042 7167
rect 19990 7124 19999 7158
rect 19999 7124 20033 7158
rect 20033 7124 20042 7158
rect 22294 7158 22346 7167
rect 19990 7115 20042 7124
rect 18838 7084 18890 7093
rect 18838 7050 18847 7084
rect 18847 7050 18881 7084
rect 18881 7050 18890 7084
rect 18838 7041 18890 7050
rect 22294 7124 22303 7158
rect 22303 7124 22337 7158
rect 22337 7124 22346 7158
rect 22294 7115 22346 7124
rect 21238 7041 21290 7093
rect 21910 7084 21962 7093
rect 21910 7050 21919 7084
rect 21919 7050 21953 7084
rect 21953 7050 21962 7084
rect 21910 7041 21962 7050
rect 23254 7115 23306 7167
rect 23830 7158 23882 7167
rect 23830 7124 23839 7158
rect 23839 7124 23873 7158
rect 23873 7124 23882 7158
rect 26038 7158 26090 7167
rect 23830 7115 23882 7124
rect 26038 7124 26047 7158
rect 26047 7124 26081 7158
rect 26081 7124 26090 7158
rect 26806 7158 26858 7167
rect 26038 7115 26090 7124
rect 25654 7084 25706 7093
rect 25654 7050 25663 7084
rect 25663 7050 25697 7084
rect 25697 7050 25706 7084
rect 25654 7041 25706 7050
rect 26806 7124 26815 7158
rect 26815 7124 26849 7158
rect 26849 7124 26858 7158
rect 27574 7158 27626 7167
rect 26806 7115 26858 7124
rect 27574 7124 27583 7158
rect 27583 7124 27617 7158
rect 27617 7124 27626 7158
rect 30550 7158 30602 7167
rect 27574 7115 27626 7124
rect 30550 7124 30559 7158
rect 30559 7124 30593 7158
rect 30593 7124 30602 7158
rect 38134 7158 38186 7167
rect 30550 7115 30602 7124
rect 28054 7041 28106 7093
rect 29494 7084 29546 7093
rect 20662 6967 20714 7019
rect 23158 6967 23210 7019
rect 29494 7050 29503 7084
rect 29503 7050 29537 7084
rect 29537 7050 29546 7084
rect 29494 7041 29546 7050
rect 38134 7124 38143 7158
rect 38143 7124 38177 7158
rect 38177 7124 38186 7158
rect 38134 7115 38186 7124
rect 31606 7084 31658 7093
rect 31606 7050 31615 7084
rect 31615 7050 31649 7084
rect 31649 7050 31658 7084
rect 31606 7041 31658 7050
rect 32470 7084 32522 7093
rect 32470 7050 32479 7084
rect 32479 7050 32513 7084
rect 32513 7050 32522 7084
rect 32470 7041 32522 7050
rect 34006 7084 34058 7093
rect 34006 7050 34015 7084
rect 34015 7050 34049 7084
rect 34049 7050 34058 7084
rect 34006 7041 34058 7050
rect 36214 7084 36266 7093
rect 36214 7050 36223 7084
rect 36223 7050 36257 7084
rect 36257 7050 36266 7084
rect 36214 7041 36266 7050
rect 36982 7084 37034 7093
rect 36982 7050 36991 7084
rect 36991 7050 37025 7084
rect 37025 7050 37034 7084
rect 36982 7041 37034 7050
rect 37750 7084 37802 7093
rect 37750 7050 37759 7084
rect 37759 7050 37793 7084
rect 37793 7050 37802 7084
rect 37750 7041 37802 7050
rect 38518 7115 38570 7167
rect 39670 7158 39722 7167
rect 39670 7124 39679 7158
rect 39679 7124 39713 7158
rect 39713 7124 39722 7158
rect 41878 7158 41930 7167
rect 39670 7115 39722 7124
rect 41878 7124 41887 7158
rect 41887 7124 41921 7158
rect 41921 7124 41930 7158
rect 41878 7115 41930 7124
rect 42262 7158 42314 7167
rect 42262 7124 42289 7158
rect 42289 7124 42314 7158
rect 42262 7115 42314 7124
rect 37462 6967 37514 7019
rect 38998 6967 39050 7019
rect 43510 7115 43562 7167
rect 44950 7158 45002 7167
rect 44950 7124 44959 7158
rect 44959 7124 44993 7158
rect 44993 7124 45002 7158
rect 44950 7115 45002 7124
rect 43030 7084 43082 7093
rect 43030 7050 43039 7084
rect 43039 7050 43073 7084
rect 43073 7050 43082 7084
rect 43030 7041 43082 7050
rect 43414 7041 43466 7093
rect 43798 7041 43850 7093
rect 52246 7115 52298 7167
rect 48310 7084 48362 7093
rect 48310 7050 48319 7084
rect 48319 7050 48353 7084
rect 48353 7050 48362 7084
rect 48310 7041 48362 7050
rect 49078 7084 49130 7093
rect 49078 7050 49087 7084
rect 49087 7050 49121 7084
rect 49121 7050 49130 7084
rect 49078 7041 49130 7050
rect 50134 7041 50186 7093
rect 52150 7041 52202 7093
rect 52822 7084 52874 7093
rect 52822 7050 52831 7084
rect 52831 7050 52865 7084
rect 52865 7050 52874 7084
rect 52822 7041 52874 7050
rect 13462 6893 13514 6945
rect 14614 6893 14666 6945
rect 15382 6893 15434 6945
rect 17110 6893 17162 6945
rect 17878 6893 17930 6945
rect 18550 6893 18602 6945
rect 20374 6936 20426 6945
rect 20374 6902 20383 6936
rect 20383 6902 20417 6936
rect 20417 6902 20426 6936
rect 20374 6893 20426 6902
rect 20662 6819 20714 6871
rect 21142 6893 21194 6945
rect 21910 6893 21962 6945
rect 23350 6893 23402 6945
rect 24214 6936 24266 6945
rect 24214 6902 24223 6936
rect 24223 6902 24257 6936
rect 24257 6902 24266 6936
rect 24214 6893 24266 6902
rect 24502 6893 24554 6945
rect 25174 6819 25226 6871
rect 26902 6893 26954 6945
rect 26998 6819 27050 6871
rect 29398 6936 29450 6945
rect 27766 6819 27818 6871
rect 29398 6902 29407 6936
rect 29407 6902 29441 6936
rect 29441 6902 29450 6936
rect 29398 6893 29450 6902
rect 29974 6893 30026 6945
rect 31798 6893 31850 6945
rect 32374 6936 32426 6945
rect 32374 6902 32383 6936
rect 32383 6902 32417 6936
rect 32417 6902 32426 6936
rect 32374 6893 32426 6902
rect 32182 6819 32234 6871
rect 32950 6745 33002 6797
rect 34582 6893 34634 6945
rect 35734 6893 35786 6945
rect 35926 6893 35978 6945
rect 36406 6893 36458 6945
rect 36982 6893 37034 6945
rect 38518 6936 38570 6945
rect 38518 6902 38527 6936
rect 38527 6902 38561 6936
rect 38561 6902 38570 6936
rect 38518 6893 38570 6902
rect 37654 6745 37706 6797
rect 39862 6819 39914 6871
rect 41878 6893 41930 6945
rect 54742 7010 54794 7019
rect 41110 6745 41162 6797
rect 43798 6936 43850 6945
rect 43798 6902 43807 6936
rect 43807 6902 43841 6936
rect 43841 6902 43850 6936
rect 43798 6893 43850 6902
rect 43606 6819 43658 6871
rect 43414 6788 43466 6797
rect 43414 6754 43423 6788
rect 43423 6754 43457 6788
rect 43457 6754 43466 6788
rect 43414 6745 43466 6754
rect 44278 6745 44330 6797
rect 45430 6893 45482 6945
rect 46774 6893 46826 6945
rect 46870 6819 46922 6871
rect 48310 6893 48362 6945
rect 50134 6893 50186 6945
rect 51382 6893 51434 6945
rect 52438 6893 52490 6945
rect 54742 6976 54751 7010
rect 54751 6976 54785 7010
rect 54785 6976 54794 7010
rect 54742 6967 54794 6976
rect 55414 6967 55466 7019
rect 58486 6967 58538 7019
rect 56374 6893 56426 6945
rect 4294 6634 4346 6686
rect 4358 6634 4410 6686
rect 4422 6634 4474 6686
rect 4486 6634 4538 6686
rect 35014 6634 35066 6686
rect 35078 6634 35130 6686
rect 35142 6634 35194 6686
rect 35206 6634 35258 6686
rect 15094 6566 15146 6575
rect 15094 6532 15103 6566
rect 15103 6532 15137 6566
rect 15137 6532 15146 6566
rect 15862 6566 15914 6575
rect 15094 6523 15146 6532
rect 8950 6449 9002 6501
rect 5686 6418 5738 6427
rect 5686 6384 5695 6418
rect 5695 6384 5729 6418
rect 5729 6384 5738 6418
rect 5686 6375 5738 6384
rect 7126 6418 7178 6427
rect 7126 6384 7135 6418
rect 7135 6384 7169 6418
rect 7169 6384 7178 6418
rect 7126 6375 7178 6384
rect 13942 6418 13994 6427
rect 13942 6384 13951 6418
rect 13951 6384 13985 6418
rect 13985 6384 13994 6418
rect 13942 6375 13994 6384
rect 14710 6418 14762 6427
rect 14710 6384 14719 6418
rect 14719 6384 14753 6418
rect 14753 6384 14762 6418
rect 14710 6375 14762 6384
rect 15862 6532 15871 6566
rect 15871 6532 15905 6566
rect 15905 6532 15914 6566
rect 15862 6523 15914 6532
rect 20566 6523 20618 6575
rect 24118 6566 24170 6575
rect 17686 6418 17738 6427
rect 1558 6344 1610 6353
rect 1558 6310 1567 6344
rect 1567 6310 1601 6344
rect 1601 6310 1610 6344
rect 1558 6301 1610 6310
rect 2038 6301 2090 6353
rect 3190 6344 3242 6353
rect 3190 6310 3199 6344
rect 3199 6310 3233 6344
rect 3233 6310 3242 6344
rect 3190 6301 3242 6310
rect 3862 6301 3914 6353
rect 4630 6301 4682 6353
rect 9430 6344 9482 6353
rect 9430 6310 9439 6344
rect 9439 6310 9473 6344
rect 9473 6310 9482 6344
rect 9430 6301 9482 6310
rect 10102 6301 10154 6353
rect 10870 6301 10922 6353
rect 11638 6301 11690 6353
rect 12310 6301 12362 6353
rect 14902 6301 14954 6353
rect 17686 6384 17695 6418
rect 17695 6384 17729 6418
rect 17729 6384 17738 6418
rect 17686 6375 17738 6384
rect 18454 6418 18506 6427
rect 18454 6384 18463 6418
rect 18463 6384 18497 6418
rect 18497 6384 18506 6418
rect 18454 6375 18506 6384
rect 19222 6418 19274 6427
rect 19222 6384 19231 6418
rect 19231 6384 19265 6418
rect 19265 6384 19274 6418
rect 19222 6375 19274 6384
rect 20470 6375 20522 6427
rect 24118 6532 24127 6566
rect 24127 6532 24161 6566
rect 24161 6532 24170 6566
rect 27862 6566 27914 6575
rect 24118 6523 24170 6532
rect 21526 6418 21578 6427
rect 19318 6301 19370 6353
rect 21526 6384 21535 6418
rect 21535 6384 21569 6418
rect 21569 6384 21578 6418
rect 21526 6375 21578 6384
rect 22966 6418 23018 6427
rect 22966 6384 22975 6418
rect 22975 6384 23009 6418
rect 23009 6384 23018 6418
rect 22966 6375 23018 6384
rect 23638 6418 23690 6427
rect 23638 6384 23647 6418
rect 23647 6384 23681 6418
rect 23681 6384 23690 6418
rect 23638 6375 23690 6384
rect 27862 6532 27871 6566
rect 27871 6532 27905 6566
rect 27905 6532 27914 6566
rect 33142 6566 33194 6575
rect 27862 6523 27914 6532
rect 33142 6532 33151 6566
rect 33151 6532 33185 6566
rect 33185 6532 33194 6566
rect 34678 6566 34730 6575
rect 33142 6523 33194 6532
rect 29014 6418 29066 6427
rect 29014 6384 29023 6418
rect 29023 6384 29057 6418
rect 29057 6384 29066 6418
rect 29014 6375 29066 6384
rect 34678 6532 34687 6566
rect 34687 6532 34721 6566
rect 34721 6532 34730 6566
rect 34678 6523 34730 6532
rect 34294 6418 34346 6427
rect 34294 6384 34303 6418
rect 34303 6384 34337 6418
rect 34337 6384 34346 6418
rect 34294 6375 34346 6384
rect 35734 6523 35786 6575
rect 41302 6523 41354 6575
rect 42262 6523 42314 6575
rect 57046 6449 57098 6501
rect 25654 6344 25706 6353
rect 25654 6310 25663 6344
rect 25663 6310 25697 6344
rect 25697 6310 25706 6344
rect 25654 6301 25706 6310
rect 26806 6344 26858 6353
rect 26806 6310 26815 6344
rect 26815 6310 26849 6344
rect 26849 6310 26858 6344
rect 26806 6301 26858 6310
rect 29686 6344 29738 6353
rect 29686 6310 29695 6344
rect 29695 6310 29729 6344
rect 29729 6310 29738 6344
rect 29686 6301 29738 6310
rect 31222 6344 31274 6353
rect 31222 6310 31231 6344
rect 31231 6310 31265 6344
rect 31265 6310 31274 6344
rect 31222 6301 31274 6310
rect 33814 6301 33866 6353
rect 35446 6375 35498 6427
rect 41206 6418 41258 6427
rect 41206 6384 41215 6418
rect 41215 6384 41249 6418
rect 41249 6384 41258 6418
rect 41206 6375 41258 6384
rect 42838 6418 42890 6427
rect 42838 6384 42847 6418
rect 42847 6384 42881 6418
rect 42881 6384 42890 6418
rect 42838 6375 42890 6384
rect 44086 6418 44138 6427
rect 44086 6384 44095 6418
rect 44095 6384 44129 6418
rect 44129 6384 44138 6418
rect 44086 6375 44138 6384
rect 44662 6375 44714 6427
rect 50806 6418 50858 6427
rect 50806 6384 50815 6418
rect 50815 6384 50849 6418
rect 50849 6384 50858 6418
rect 50806 6375 50858 6384
rect 51574 6418 51626 6427
rect 51574 6384 51583 6418
rect 51583 6384 51617 6418
rect 51617 6384 51626 6418
rect 51574 6375 51626 6384
rect 36310 6344 36362 6353
rect 36310 6310 36319 6344
rect 36319 6310 36353 6344
rect 36353 6310 36362 6344
rect 36310 6301 36362 6310
rect 38902 6344 38954 6353
rect 38902 6310 38911 6344
rect 38911 6310 38945 6344
rect 38945 6310 38954 6344
rect 38902 6301 38954 6310
rect 40342 6344 40394 6353
rect 40342 6310 40351 6344
rect 40351 6310 40385 6344
rect 40385 6310 40394 6344
rect 40342 6301 40394 6310
rect 41878 6344 41930 6353
rect 41878 6310 41887 6344
rect 41887 6310 41921 6344
rect 41921 6310 41930 6344
rect 41878 6301 41930 6310
rect 45526 6344 45578 6353
rect 45526 6310 45535 6344
rect 45535 6310 45569 6344
rect 45569 6310 45578 6344
rect 45526 6301 45578 6310
rect 46966 6344 47018 6353
rect 46966 6310 46975 6344
rect 46975 6310 47009 6344
rect 47009 6310 47018 6344
rect 46966 6301 47018 6310
rect 47734 6344 47786 6353
rect 47734 6310 47743 6344
rect 47743 6310 47777 6344
rect 47777 6310 47786 6344
rect 47734 6301 47786 6310
rect 48790 6301 48842 6353
rect 49558 6301 49610 6353
rect 53974 6301 54026 6353
rect 55222 6344 55274 6353
rect 55222 6310 55231 6344
rect 55231 6310 55265 6344
rect 55265 6310 55274 6344
rect 55222 6301 55274 6310
rect 30646 6270 30698 6279
rect 30646 6236 30655 6270
rect 30655 6236 30689 6270
rect 30689 6236 30698 6270
rect 30646 6227 30698 6236
rect 8086 6153 8138 6205
rect 8374 6153 8426 6205
rect 14134 6153 14186 6205
rect 5494 6079 5546 6131
rect 6262 6079 6314 6131
rect 13078 6079 13130 6131
rect 13942 6079 13994 6131
rect 16822 6153 16874 6205
rect 18262 6153 18314 6205
rect 18358 6122 18410 6131
rect 18358 6088 18367 6122
rect 18367 6088 18401 6122
rect 18401 6088 18410 6122
rect 18358 6079 18410 6088
rect 18934 6153 18986 6205
rect 36886 6227 36938 6279
rect 40630 6227 40682 6279
rect 21430 6122 21482 6131
rect 21430 6088 21439 6122
rect 21439 6088 21473 6122
rect 21473 6088 21482 6122
rect 21430 6079 21482 6088
rect 21526 6079 21578 6131
rect 23638 6079 23690 6131
rect 23926 6079 23978 6131
rect 26326 6079 26378 6131
rect 40822 6153 40874 6205
rect 28438 6079 28490 6131
rect 29782 6079 29834 6131
rect 30742 6079 30794 6131
rect 33526 6122 33578 6131
rect 33526 6088 33535 6122
rect 33535 6088 33569 6122
rect 33569 6088 33578 6122
rect 33526 6079 33578 6088
rect 33718 6079 33770 6131
rect 36886 6122 36938 6131
rect 36886 6088 36895 6122
rect 36895 6088 36929 6122
rect 36929 6088 36938 6122
rect 36886 6079 36938 6088
rect 39958 6079 40010 6131
rect 55126 6227 55178 6279
rect 42646 6153 42698 6205
rect 51574 6153 51626 6205
rect 44086 6079 44138 6131
rect 49750 6079 49802 6131
rect 51094 6079 51146 6131
rect 55030 6153 55082 6205
rect 58102 6301 58154 6353
rect 58870 6227 58922 6279
rect 19654 5968 19706 6020
rect 19718 5968 19770 6020
rect 19782 5968 19834 6020
rect 19846 5968 19898 6020
rect 50374 5968 50426 6020
rect 50438 5968 50490 6020
rect 50502 5968 50554 6020
rect 50566 5968 50618 6020
rect 5782 5857 5834 5909
rect 17590 5857 17642 5909
rect 2614 5783 2666 5835
rect 8374 5783 8426 5835
rect 8854 5783 8906 5835
rect 9814 5783 9866 5835
rect 5014 5709 5066 5761
rect 7030 5709 7082 5761
rect 1078 5635 1130 5687
rect 2902 5678 2954 5687
rect 2902 5644 2911 5678
rect 2911 5644 2945 5678
rect 2945 5644 2954 5678
rect 2902 5635 2954 5644
rect 4918 5635 4970 5687
rect 5110 5678 5162 5687
rect 5110 5644 5119 5678
rect 5119 5644 5153 5678
rect 5153 5644 5162 5678
rect 5110 5635 5162 5644
rect 6838 5678 6890 5687
rect 6838 5644 6847 5678
rect 6847 5644 6881 5678
rect 6881 5644 6890 5678
rect 6838 5635 6890 5644
rect 7222 5635 7274 5687
rect 5782 5487 5834 5539
rect 7606 5487 7658 5539
rect 8758 5635 8810 5687
rect 43414 5709 43466 5761
rect 10198 5635 10250 5687
rect 10486 5635 10538 5687
rect 12598 5678 12650 5687
rect 12598 5644 12607 5678
rect 12607 5644 12641 5678
rect 12641 5644 12650 5678
rect 12598 5635 12650 5644
rect 13366 5678 13418 5687
rect 13366 5644 13375 5678
rect 13375 5644 13409 5678
rect 13409 5644 13418 5678
rect 13366 5635 13418 5644
rect 14998 5678 15050 5687
rect 14998 5644 15007 5678
rect 15007 5644 15041 5678
rect 15041 5644 15050 5678
rect 14998 5635 15050 5644
rect 15862 5678 15914 5687
rect 15862 5644 15871 5678
rect 15871 5644 15905 5678
rect 15905 5644 15914 5678
rect 15862 5635 15914 5644
rect 16246 5635 16298 5687
rect 17302 5678 17354 5687
rect 17302 5644 17311 5678
rect 17311 5644 17345 5678
rect 17345 5644 17354 5678
rect 18742 5678 18794 5687
rect 17302 5635 17354 5644
rect 18742 5644 18751 5678
rect 18751 5644 18785 5678
rect 18785 5644 18794 5678
rect 18742 5635 18794 5644
rect 20182 5678 20234 5687
rect 20182 5644 20191 5678
rect 20191 5644 20225 5678
rect 20225 5644 20234 5678
rect 20182 5635 20234 5644
rect 20566 5635 20618 5687
rect 21814 5635 21866 5687
rect 23062 5635 23114 5687
rect 23446 5635 23498 5687
rect 24598 5635 24650 5687
rect 26230 5678 26282 5687
rect 26230 5644 26239 5678
rect 26239 5644 26273 5678
rect 26273 5644 26282 5678
rect 26230 5635 26282 5644
rect 27382 5635 27434 5687
rect 27862 5635 27914 5687
rect 28822 5635 28874 5687
rect 30262 5635 30314 5687
rect 30838 5635 30890 5687
rect 31702 5635 31754 5687
rect 33142 5678 33194 5687
rect 33142 5644 33151 5678
rect 33151 5644 33185 5678
rect 33185 5644 33194 5678
rect 33142 5635 33194 5644
rect 33238 5635 33290 5687
rect 34678 5678 34730 5687
rect 34678 5644 34687 5678
rect 34687 5644 34721 5678
rect 34721 5644 34730 5678
rect 34678 5635 34730 5644
rect 36022 5678 36074 5687
rect 36022 5644 36031 5678
rect 36031 5644 36065 5678
rect 36065 5644 36074 5678
rect 36022 5635 36074 5644
rect 36214 5635 36266 5687
rect 37558 5678 37610 5687
rect 37558 5644 37567 5678
rect 37567 5644 37601 5678
rect 37601 5644 37610 5678
rect 37558 5635 37610 5644
rect 39094 5678 39146 5687
rect 36886 5561 36938 5613
rect 37462 5561 37514 5613
rect 39094 5644 39103 5678
rect 39103 5644 39137 5678
rect 39137 5644 39146 5678
rect 39094 5635 39146 5644
rect 39286 5635 39338 5687
rect 40726 5635 40778 5687
rect 42070 5678 42122 5687
rect 42070 5644 42079 5678
rect 42079 5644 42113 5678
rect 42113 5644 42122 5678
rect 42070 5635 42122 5644
rect 42262 5635 42314 5687
rect 43222 5635 43274 5687
rect 43702 5635 43754 5687
rect 44662 5635 44714 5687
rect 46102 5635 46154 5687
rect 46678 5635 46730 5687
rect 47542 5635 47594 5687
rect 48982 5678 49034 5687
rect 48982 5644 48991 5678
rect 48991 5644 49025 5678
rect 49025 5644 49034 5678
rect 48982 5635 49034 5644
rect 49654 5678 49706 5687
rect 49654 5644 49663 5678
rect 49663 5644 49697 5678
rect 49697 5644 49706 5678
rect 49654 5635 49706 5644
rect 50710 5635 50762 5687
rect 52150 5678 52202 5687
rect 52150 5644 52159 5678
rect 52159 5644 52193 5678
rect 52193 5644 52202 5678
rect 52150 5635 52202 5644
rect 52534 5635 52586 5687
rect 53686 5678 53738 5687
rect 53686 5644 53695 5678
rect 53695 5644 53729 5678
rect 53729 5644 53738 5678
rect 53686 5635 53738 5644
rect 57430 5678 57482 5687
rect 53590 5561 53642 5613
rect 57430 5644 57439 5678
rect 57439 5644 57473 5678
rect 57473 5644 57482 5678
rect 57430 5635 57482 5644
rect 59638 5561 59690 5613
rect 21718 5487 21770 5539
rect 26038 5487 26090 5539
rect 6166 5413 6218 5465
rect 17782 5413 17834 5465
rect 38998 5487 39050 5539
rect 30646 5413 30698 5465
rect 4294 5302 4346 5354
rect 4358 5302 4410 5354
rect 4422 5302 4474 5354
rect 4486 5302 4538 5354
rect 35014 5302 35066 5354
rect 35078 5302 35130 5354
rect 35142 5302 35194 5354
rect 35206 5302 35258 5354
rect 4726 5191 4778 5243
rect 57142 5191 57194 5243
rect 310 4969 362 5021
rect 1846 4969 1898 5021
rect 3094 5012 3146 5021
rect 3094 4978 3103 5012
rect 3103 4978 3137 5012
rect 3137 4978 3146 5012
rect 3094 4969 3146 4978
rect 4150 5012 4202 5021
rect 4150 4978 4159 5012
rect 4159 4978 4193 5012
rect 4193 4978 4202 5012
rect 4150 4969 4202 4978
rect 5398 5012 5450 5021
rect 5398 4978 5407 5012
rect 5407 4978 5441 5012
rect 5441 4978 5450 5012
rect 5398 4969 5450 4978
rect 6070 4969 6122 5021
rect 9238 5012 9290 5021
rect 9238 4978 9247 5012
rect 9247 4978 9281 5012
rect 9281 4978 9290 5012
rect 9238 4969 9290 4978
rect 10006 5012 10058 5021
rect 10006 4978 10015 5012
rect 10015 4978 10049 5012
rect 10049 4978 10058 5012
rect 10006 4969 10058 4978
rect 10678 4969 10730 5021
rect 11830 4969 11882 5021
rect 12982 5012 13034 5021
rect 12982 4978 12991 5012
rect 12991 4978 13025 5012
rect 13025 4978 13034 5012
rect 12982 4969 13034 4978
rect 13942 5012 13994 5021
rect 13942 4978 13951 5012
rect 13951 4978 13985 5012
rect 13985 4978 13994 5012
rect 13942 4969 13994 4978
rect 14422 4969 14474 5021
rect 14806 4969 14858 5021
rect 16534 4969 16586 5021
rect 17494 5012 17546 5021
rect 17494 4978 17503 5012
rect 17503 4978 17537 5012
rect 17537 4978 17546 5012
rect 17494 4969 17546 4978
rect 17974 4969 18026 5021
rect 19030 5012 19082 5021
rect 19030 4978 19039 5012
rect 19039 4978 19073 5012
rect 19073 4978 19082 5012
rect 19030 4969 19082 4978
rect 19126 4969 19178 5021
rect 20662 5012 20714 5021
rect 20662 4978 20671 5012
rect 20671 4978 20705 5012
rect 20705 4978 20714 5012
rect 20662 4969 20714 4978
rect 20854 4969 20906 5021
rect 22774 5012 22826 5021
rect 22774 4978 22783 5012
rect 22783 4978 22817 5012
rect 22817 4978 22826 5012
rect 22774 4969 22826 4978
rect 23542 5012 23594 5021
rect 23542 4978 23551 5012
rect 23551 4978 23585 5012
rect 23585 4978 23594 5012
rect 23542 4969 23594 4978
rect 25078 5012 25130 5021
rect 7942 4895 7994 4947
rect 23158 4895 23210 4947
rect 25078 4978 25087 5012
rect 25087 4978 25121 5012
rect 25121 4978 25130 5012
rect 25078 4969 25130 4978
rect 26614 5012 26666 5021
rect 24886 4895 24938 4947
rect 26614 4978 26623 5012
rect 26623 4978 26657 5012
rect 26657 4978 26666 5012
rect 26614 4969 26666 4978
rect 28054 5012 28106 5021
rect 28054 4978 28063 5012
rect 28063 4978 28097 5012
rect 28097 4978 28106 5012
rect 28054 4969 28106 4978
rect 28918 5012 28970 5021
rect 28918 4978 28927 5012
rect 28927 4978 28961 5012
rect 28961 4978 28970 5012
rect 28918 4969 28970 4978
rect 29302 4969 29354 5021
rect 30358 5012 30410 5021
rect 30358 4978 30367 5012
rect 30367 4978 30401 5012
rect 30401 4978 30410 5012
rect 30358 4969 30410 4978
rect 31126 5012 31178 5021
rect 31126 4978 31135 5012
rect 31135 4978 31169 5012
rect 31169 4978 31178 5012
rect 31126 4969 31178 4978
rect 31894 5012 31946 5021
rect 31894 4978 31903 5012
rect 31903 4978 31937 5012
rect 31937 4978 31946 5012
rect 31894 4969 31946 4978
rect 33334 5012 33386 5021
rect 33334 4978 33343 5012
rect 33343 4978 33377 5012
rect 33377 4978 33386 5012
rect 33334 4969 33386 4978
rect 34102 5012 34154 5021
rect 34102 4978 34111 5012
rect 34111 4978 34145 5012
rect 34145 4978 34154 5012
rect 34102 4969 34154 4978
rect 34870 5012 34922 5021
rect 34870 4978 34879 5012
rect 34879 4978 34913 5012
rect 34913 4978 34922 5012
rect 34870 4969 34922 4978
rect 35350 4969 35402 5021
rect 36118 4969 36170 5021
rect 36886 4969 36938 5021
rect 38614 5012 38666 5021
rect 38614 4978 38623 5012
rect 38623 4978 38657 5012
rect 38657 4978 38666 5012
rect 38614 4969 38666 4978
rect 39382 5012 39434 5021
rect 39382 4978 39391 5012
rect 39391 4978 39425 5012
rect 39425 4978 39434 5012
rect 39382 4969 39434 4978
rect 39574 4969 39626 5021
rect 40918 5012 40970 5021
rect 40918 4978 40927 5012
rect 40927 4978 40961 5012
rect 40961 4978 40970 5012
rect 40918 4969 40970 4978
rect 41686 5012 41738 5021
rect 41686 4978 41695 5012
rect 41695 4978 41729 5012
rect 41729 4978 41738 5012
rect 41686 4969 41738 4978
rect 42166 4969 42218 5021
rect 43318 4969 43370 5021
rect 44854 4969 44906 5021
rect 45430 5012 45482 5021
rect 45430 4978 45439 5012
rect 45439 4978 45473 5012
rect 45473 4978 45482 5012
rect 45430 4969 45482 4978
rect 46198 5012 46250 5021
rect 46198 4978 46207 5012
rect 46207 4978 46241 5012
rect 46241 4978 46250 5012
rect 46198 4969 46250 4978
rect 46294 4969 46346 5021
rect 47638 4969 47690 5021
rect 49366 5012 49418 5021
rect 49366 4978 49375 5012
rect 49375 4978 49409 5012
rect 49409 4978 49418 5012
rect 49366 4969 49418 4978
rect 50422 5012 50474 5021
rect 50422 4978 50431 5012
rect 50431 4978 50465 5012
rect 50465 4978 50474 5012
rect 50422 4969 50474 4978
rect 50902 4969 50954 5021
rect 51862 5012 51914 5021
rect 51862 4978 51871 5012
rect 51871 4978 51905 5012
rect 51905 4978 51914 5012
rect 51862 4969 51914 4978
rect 52246 4969 52298 5021
rect 53302 4969 53354 5021
rect 57046 5012 57098 5021
rect 8374 4821 8426 4873
rect 57046 4978 57055 5012
rect 57055 4978 57089 5012
rect 57089 4978 57098 5012
rect 57046 4969 57098 4978
rect 57814 4895 57866 4947
rect 59254 4821 59306 4873
rect 19654 4636 19706 4688
rect 19718 4636 19770 4688
rect 19782 4636 19834 4688
rect 19846 4636 19898 4688
rect 50374 4636 50426 4688
rect 50438 4636 50490 4688
rect 50502 4636 50554 4688
rect 50566 4636 50618 4688
rect 790 4377 842 4429
rect 1174 4303 1226 4355
rect 14038 4377 14090 4429
rect 1366 4229 1418 4281
rect 3766 4229 3818 4281
rect 4726 4303 4778 4355
rect 5014 4229 5066 4281
rect 7414 4346 7466 4355
rect 5686 4229 5738 4281
rect 7414 4312 7423 4346
rect 7423 4312 7457 4346
rect 7457 4312 7466 4346
rect 7414 4303 7466 4312
rect 9622 4346 9674 4355
rect 3478 4155 3530 4207
rect 4918 4155 4970 4207
rect 6454 4155 6506 4207
rect 9622 4312 9631 4346
rect 9631 4312 9665 4346
rect 9665 4312 9674 4346
rect 9622 4303 9674 4312
rect 10390 4346 10442 4355
rect 10390 4312 10399 4346
rect 10399 4312 10433 4346
rect 10433 4312 10442 4346
rect 10390 4303 10442 4312
rect 10774 4303 10826 4355
rect 13558 4346 13610 4355
rect 9814 4229 9866 4281
rect 10198 4229 10250 4281
rect 11158 4155 11210 4207
rect 3958 4081 4010 4133
rect 5110 4081 5162 4133
rect 9046 4081 9098 4133
rect 10678 4081 10730 4133
rect 11446 4081 11498 4133
rect 13558 4312 13567 4346
rect 13567 4312 13601 4346
rect 13601 4312 13610 4346
rect 13558 4303 13610 4312
rect 15478 4346 15530 4355
rect 15478 4312 15487 4346
rect 15487 4312 15521 4346
rect 15521 4312 15530 4346
rect 15478 4303 15530 4312
rect 15958 4303 16010 4355
rect 16438 4303 16490 4355
rect 16918 4229 16970 4281
rect 20278 4346 20330 4355
rect 17590 4229 17642 4281
rect 20278 4312 20287 4346
rect 20287 4312 20321 4346
rect 20321 4312 20330 4346
rect 20278 4303 20330 4312
rect 21046 4346 21098 4355
rect 21046 4312 21055 4346
rect 21055 4312 21089 4346
rect 21089 4312 21098 4346
rect 21046 4303 21098 4312
rect 21814 4346 21866 4355
rect 21814 4312 21823 4346
rect 21823 4312 21857 4346
rect 21857 4312 21866 4346
rect 21814 4303 21866 4312
rect 23254 4346 23306 4355
rect 23254 4312 23263 4346
rect 23263 4312 23297 4346
rect 23297 4312 23306 4346
rect 23254 4303 23306 4312
rect 25462 4346 25514 4355
rect 22006 4229 22058 4281
rect 25462 4312 25471 4346
rect 25471 4312 25505 4346
rect 25505 4312 25514 4346
rect 25462 4303 25514 4312
rect 26134 4303 26186 4355
rect 26518 4303 26570 4355
rect 28342 4346 28394 4355
rect 28342 4312 28351 4346
rect 28351 4312 28385 4346
rect 28385 4312 28394 4346
rect 28342 4303 28394 4312
rect 29110 4346 29162 4355
rect 29110 4312 29119 4346
rect 29119 4312 29153 4346
rect 29153 4312 29162 4346
rect 29110 4303 29162 4312
rect 30934 4346 30986 4355
rect 30934 4312 30943 4346
rect 30943 4312 30977 4346
rect 30977 4312 30986 4346
rect 30934 4303 30986 4312
rect 31702 4346 31754 4355
rect 31702 4312 31711 4346
rect 31711 4312 31745 4346
rect 31745 4312 31754 4346
rect 31702 4303 31754 4312
rect 32758 4346 32810 4355
rect 32758 4312 32767 4346
rect 32767 4312 32801 4346
rect 32801 4312 32810 4346
rect 32758 4303 32810 4312
rect 33910 4346 33962 4355
rect 33910 4312 33919 4346
rect 33919 4312 33953 4346
rect 33953 4312 33962 4346
rect 33910 4303 33962 4312
rect 34582 4303 34634 4355
rect 34198 4229 34250 4281
rect 36790 4346 36842 4355
rect 36790 4312 36799 4346
rect 36799 4312 36833 4346
rect 36833 4312 36842 4346
rect 36790 4303 36842 4312
rect 37174 4229 37226 4281
rect 38998 4346 39050 4355
rect 38998 4312 39007 4346
rect 39007 4312 39041 4346
rect 39041 4312 39050 4346
rect 38998 4303 39050 4312
rect 39766 4346 39818 4355
rect 39766 4312 39775 4346
rect 39775 4312 39809 4346
rect 39809 4312 39818 4346
rect 39766 4303 39818 4312
rect 41974 4346 42026 4355
rect 41974 4312 41983 4346
rect 41983 4312 42017 4346
rect 42017 4312 42026 4346
rect 41974 4303 42026 4312
rect 42358 4303 42410 4355
rect 43414 4303 43466 4355
rect 44950 4346 45002 4355
rect 44950 4312 44959 4346
rect 44959 4312 44993 4346
rect 44993 4312 45002 4346
rect 44950 4303 45002 4312
rect 46774 4346 46826 4355
rect 46774 4312 46783 4346
rect 46783 4312 46817 4346
rect 46817 4312 46826 4346
rect 46774 4303 46826 4312
rect 47446 4229 47498 4281
rect 47830 4303 47882 4355
rect 49846 4346 49898 4355
rect 48598 4229 48650 4281
rect 49846 4312 49855 4346
rect 49855 4312 49889 4346
rect 49889 4312 49898 4346
rect 49846 4303 49898 4312
rect 52630 4346 52682 4355
rect 49942 4229 49994 4281
rect 50998 4229 51050 4281
rect 52630 4312 52639 4346
rect 52639 4312 52673 4346
rect 52673 4312 52682 4346
rect 52630 4303 52682 4312
rect 53014 4229 53066 4281
rect 54070 4303 54122 4355
rect 55606 4346 55658 4355
rect 55606 4312 55615 4346
rect 55615 4312 55649 4346
rect 55649 4312 55658 4346
rect 55606 4303 55658 4312
rect 56662 4303 56714 4355
rect 55126 4272 55178 4281
rect 55126 4238 55135 4272
rect 55135 4238 55169 4272
rect 55169 4238 55178 4272
rect 55126 4229 55178 4238
rect 56374 4229 56426 4281
rect 59446 4229 59498 4281
rect 43510 4155 43562 4207
rect 55894 4081 55946 4133
rect 57910 4081 57962 4133
rect 4294 3970 4346 4022
rect 4358 3970 4410 4022
rect 4422 3970 4474 4022
rect 4486 3970 4538 4022
rect 35014 3970 35066 4022
rect 35078 3970 35130 4022
rect 35142 3970 35194 4022
rect 35206 3970 35258 4022
rect 1942 3859 1994 3911
rect 3286 3859 3338 3911
rect 7894 3859 7946 3911
rect 9238 3859 9290 3911
rect 21238 3859 21290 3911
rect 22774 3859 22826 3911
rect 29782 3859 29834 3911
rect 31990 3859 32042 3911
rect 33526 3859 33578 3911
rect 35542 3859 35594 3911
rect 39190 3859 39242 3911
rect 57334 3859 57386 3911
rect 59158 3859 59210 3911
rect 502 3785 554 3837
rect 1654 3785 1706 3837
rect 2326 3785 2378 3837
rect 3094 3785 3146 3837
rect 8278 3785 8330 3837
rect 10006 3785 10058 3837
rect 16726 3785 16778 3837
rect 17302 3785 17354 3837
rect 19414 3785 19466 3837
rect 20662 3785 20714 3837
rect 22294 3785 22346 3837
rect 23638 3785 23690 3837
rect 26422 3785 26474 3837
rect 28054 3785 28106 3837
rect 28822 3785 28874 3837
rect 29014 3785 29066 3837
rect 30358 3785 30410 3837
rect 33430 3785 33482 3837
rect 34870 3785 34922 3837
rect 37846 3785 37898 3837
rect 39382 3785 39434 3837
rect 40054 3785 40106 3837
rect 41686 3785 41738 3837
rect 49270 3785 49322 3837
rect 50710 3785 50762 3837
rect 51286 3785 51338 3837
rect 54358 3785 54410 3837
rect 55222 3785 55274 3837
rect 57142 3785 57194 3837
rect 118 3637 170 3689
rect 1654 3637 1706 3689
rect 2710 3637 2762 3689
rect 982 3563 1034 3615
rect 2422 3563 2474 3615
rect 5206 3711 5258 3763
rect 24118 3711 24170 3763
rect 24694 3711 24746 3763
rect 28726 3711 28778 3763
rect 5590 3680 5642 3689
rect 598 3415 650 3467
rect 1462 3415 1514 3467
rect 2422 3415 2474 3467
rect 3094 3489 3146 3541
rect 3382 3415 3434 3467
rect 5590 3646 5599 3680
rect 5599 3646 5633 3680
rect 5633 3646 5642 3680
rect 5590 3637 5642 3646
rect 6358 3637 6410 3689
rect 7030 3637 7082 3689
rect 7798 3637 7850 3689
rect 8566 3637 8618 3689
rect 9334 3637 9386 3689
rect 10006 3489 10058 3541
rect 13174 3637 13226 3689
rect 13654 3680 13706 3689
rect 13654 3646 13663 3680
rect 13663 3646 13697 3680
rect 13697 3646 13706 3680
rect 13654 3637 13706 3646
rect 14038 3637 14090 3689
rect 14806 3637 14858 3689
rect 15286 3637 15338 3689
rect 17398 3637 17450 3689
rect 18070 3637 18122 3689
rect 18454 3637 18506 3689
rect 19222 3637 19274 3689
rect 19990 3637 20042 3689
rect 20662 3637 20714 3689
rect 22102 3637 22154 3689
rect 22870 3637 22922 3689
rect 23638 3637 23690 3689
rect 24406 3637 24458 3689
rect 24694 3563 24746 3615
rect 25558 3563 25610 3615
rect 25942 3563 25994 3615
rect 17302 3489 17354 3541
rect 17494 3489 17546 3541
rect 22582 3489 22634 3541
rect 23350 3489 23402 3541
rect 25846 3489 25898 3541
rect 27286 3637 27338 3689
rect 42838 3711 42890 3763
rect 43798 3711 43850 3763
rect 44566 3711 44618 3763
rect 28054 3489 28106 3541
rect 29494 3563 29546 3615
rect 30454 3637 30506 3689
rect 31318 3637 31370 3689
rect 32470 3637 32522 3689
rect 33526 3637 33578 3689
rect 34294 3637 34346 3689
rect 34966 3637 35018 3689
rect 35734 3637 35786 3689
rect 36502 3637 36554 3689
rect 37942 3637 37994 3689
rect 38710 3637 38762 3689
rect 30742 3563 30794 3615
rect 31798 3563 31850 3615
rect 31414 3489 31466 3541
rect 32374 3489 32426 3541
rect 37366 3489 37418 3541
rect 38518 3489 38570 3541
rect 39382 3489 39434 3541
rect 40150 3489 40202 3541
rect 41014 3637 41066 3689
rect 41590 3489 41642 3541
rect 42742 3637 42794 3689
rect 43798 3563 43850 3615
rect 45238 3563 45290 3615
rect 46006 3489 46058 3541
rect 47158 3637 47210 3689
rect 48214 3637 48266 3689
rect 47542 3489 47594 3541
rect 48310 3489 48362 3541
rect 55894 3711 55946 3763
rect 50710 3637 50762 3689
rect 50806 3637 50858 3689
rect 51286 3637 51338 3689
rect 52054 3637 52106 3689
rect 53398 3637 53450 3689
rect 57334 3711 57386 3763
rect 54454 3489 54506 3541
rect 55222 3415 55274 3467
rect 56278 3563 56330 3615
rect 56374 3489 56426 3541
rect 57142 3489 57194 3541
rect 19654 3304 19706 3356
rect 19718 3304 19770 3356
rect 19782 3304 19834 3356
rect 19846 3304 19898 3356
rect 50374 3304 50426 3356
rect 50438 3304 50490 3356
rect 50502 3304 50554 3356
rect 50566 3304 50618 3356
rect 1462 3193 1514 3245
rect 2134 3193 2186 3245
rect 12022 3193 12074 3245
rect 13366 3193 13418 3245
rect 17494 3193 17546 3245
rect 18358 3193 18410 3245
rect 19702 3193 19754 3245
rect 20374 3193 20426 3245
rect 23350 3193 23402 3245
rect 24214 3193 24266 3245
rect 25942 3193 25994 3245
rect 26902 3193 26954 3245
rect 27382 3193 27434 3245
rect 28438 3193 28490 3245
rect 28534 3193 28586 3245
rect 29398 3193 29450 3245
rect 30454 3193 30506 3245
rect 31894 3193 31946 3245
rect 32662 3193 32714 3245
rect 34102 3193 34154 3245
rect 38518 3193 38570 3245
rect 39574 3193 39626 3245
rect 41206 3193 41258 3245
rect 41686 3193 41738 3245
rect 44086 3193 44138 3245
rect 45430 3193 45482 3245
rect 48502 3193 48554 3245
rect 49654 3193 49706 3245
rect 52054 3193 52106 3245
rect 52438 3193 52490 3245
rect 56854 3193 56906 3245
rect 58294 3193 58346 3245
rect 214 3119 266 3171
rect 1750 3119 1802 3171
rect 12214 3119 12266 3171
rect 12982 3119 13034 3171
rect 20086 3119 20138 3171
rect 21430 3119 21482 3171
rect 22966 3119 23018 3171
rect 23926 3119 23978 3171
rect 24982 3119 25034 3171
rect 26614 3119 26666 3171
rect 28246 3119 28298 3171
rect 29302 3119 29354 3171
rect 29782 3119 29834 3171
rect 30550 3119 30602 3171
rect 31798 3119 31850 3171
rect 31990 3119 32042 3171
rect 32566 3119 32618 3171
rect 33718 3119 33770 3171
rect 35542 3119 35594 3171
rect 8950 3045 9002 3097
rect 18358 3045 18410 3097
rect 19030 3045 19082 3097
rect 19798 3045 19850 3097
rect 20182 3045 20234 3097
rect 22390 3045 22442 3097
rect 23542 3045 23594 3097
rect 23830 3045 23882 3097
rect 25078 3045 25130 3097
rect 25366 3045 25418 3097
rect 26230 3045 26282 3097
rect 27478 3045 27530 3097
rect 28918 3045 28970 3097
rect 29398 3045 29450 3097
rect 31126 3045 31178 3097
rect 31894 3045 31946 3097
rect 33334 3045 33386 3097
rect 34006 3045 34058 3097
rect 34486 3045 34538 3097
rect 37078 3119 37130 3171
rect 38614 3119 38666 3171
rect 39670 3119 39722 3171
rect 40918 3119 40970 3171
rect 41110 3119 41162 3171
rect 42166 3119 42218 3171
rect 44854 3119 44906 3171
rect 45142 3119 45194 3171
rect 46294 3119 46346 3171
rect 48118 3119 48170 3171
rect 48982 3119 49034 3171
rect 57334 3119 57386 3171
rect 58006 3119 58058 3171
rect 35926 3045 35978 3097
rect 36118 3045 36170 3097
rect 36694 3045 36746 3097
rect 37558 3045 37610 3097
rect 38326 3045 38378 3097
rect 22 2971 74 3023
rect 694 2897 746 2949
rect 2134 2897 2186 2949
rect 4918 3014 4970 3023
rect 4918 2980 4927 3014
rect 4927 2980 4961 3014
rect 4961 2980 4970 3014
rect 4918 2971 4970 2980
rect 5206 2971 5258 3023
rect 5974 2971 6026 3023
rect 6742 2897 6794 2949
rect 8182 2971 8234 3023
rect 12982 3014 13034 3023
rect 8950 2897 9002 2949
rect 12982 2980 12991 3014
rect 12991 2980 13025 3014
rect 13025 2980 13034 3014
rect 12982 2971 13034 2980
rect 13366 2971 13418 3023
rect 14518 2971 14570 3023
rect 16630 3014 16682 3023
rect 16630 2980 16639 3014
rect 16639 2980 16673 3014
rect 16673 2980 16682 3014
rect 16630 2971 16682 2980
rect 17014 2971 17066 3023
rect 15382 2897 15434 2949
rect 16534 2897 16586 2949
rect 17686 2897 17738 2949
rect 18838 2971 18890 3023
rect 19606 2897 19658 2949
rect 21430 2971 21482 3023
rect 20950 2897 21002 2949
rect 21718 2897 21770 2949
rect 22486 2897 22538 2949
rect 24022 2971 24074 3023
rect 24214 2897 24266 2949
rect 24886 2897 24938 2949
rect 25078 2897 25130 2949
rect 26902 2971 26954 3023
rect 27670 2897 27722 2949
rect 29878 2971 29930 3023
rect 30550 2897 30602 2949
rect 32086 2971 32138 3023
rect 32278 2897 32330 2949
rect 33142 2897 33194 2949
rect 33334 2897 33386 2949
rect 35350 2971 35402 3023
rect 37270 2971 37322 3023
rect 40822 3045 40874 3097
rect 41206 3045 41258 3097
rect 40534 2971 40586 3023
rect 42166 2971 42218 3023
rect 42646 2971 42698 3023
rect 43222 3045 43274 3097
rect 44758 3045 44810 3097
rect 46198 3045 46250 3097
rect 46390 3045 46442 3097
rect 43030 2971 43082 3023
rect 35446 2897 35498 2949
rect 36022 2897 36074 2949
rect 37558 2897 37610 2949
rect 38134 2897 38186 2949
rect 39094 2897 39146 2949
rect 39190 2897 39242 2949
rect 39958 2897 40010 2949
rect 2614 2823 2666 2875
rect 5110 2749 5162 2801
rect 5782 2749 5834 2801
rect 8758 2792 8810 2801
rect 8758 2758 8767 2792
rect 8767 2758 8801 2792
rect 8801 2758 8810 2792
rect 8758 2749 8810 2758
rect 14230 2823 14282 2875
rect 33814 2749 33866 2801
rect 40822 2823 40874 2875
rect 41494 2897 41546 2949
rect 42070 2897 42122 2949
rect 42550 2897 42602 2949
rect 43318 2897 43370 2949
rect 44182 2897 44234 2949
rect 45622 2971 45674 3023
rect 51766 3045 51818 3097
rect 52246 3045 52298 3097
rect 53206 3045 53258 3097
rect 49654 2971 49706 3023
rect 46294 2897 46346 2949
rect 47638 2897 47690 2949
rect 48982 2897 49034 2949
rect 49846 2897 49898 2949
rect 51478 2971 51530 3023
rect 51382 2897 51434 2949
rect 51862 2897 51914 2949
rect 52246 2897 52298 2949
rect 53782 2971 53834 3023
rect 52918 2897 52970 2949
rect 53686 2897 53738 2949
rect 54838 2897 54890 2949
rect 50038 2823 50090 2875
rect 52822 2823 52874 2875
rect 46102 2749 46154 2801
rect 46678 2749 46730 2801
rect 4294 2638 4346 2690
rect 4358 2638 4410 2690
rect 4422 2638 4474 2690
rect 4486 2638 4538 2690
rect 35014 2638 35066 2690
rect 35078 2638 35130 2690
rect 35142 2638 35194 2690
rect 35206 2638 35258 2690
rect 3958 2527 4010 2579
rect 4246 2527 4298 2579
rect 4342 2527 4394 2579
rect 4822 2527 4874 2579
rect 8758 2527 8810 2579
rect 29782 2527 29834 2579
rect 35638 2527 35690 2579
rect 36886 2527 36938 2579
rect 43222 2527 43274 2579
rect 43990 2527 44042 2579
rect 20182 2453 20234 2505
rect 20854 2453 20906 2505
rect 33814 2453 33866 2505
rect 40822 2453 40874 2505
rect 33814 2305 33866 2357
rect 34678 2305 34730 2357
rect 16246 2157 16298 2209
rect 16438 2157 16490 2209
rect 4726 2009 4778 2061
rect 5302 2009 5354 2061
rect 16534 1935 16586 1987
rect 16726 1935 16778 1987
rect 4534 1861 4586 1913
rect 4822 1861 4874 1913
rect 30358 1713 30410 1765
rect 30646 1713 30698 1765
rect 50710 1713 50762 1765
rect 50902 1713 50954 1765
rect 35350 1639 35402 1691
rect 36310 1639 36362 1691
rect 50518 1639 50570 1691
rect 51094 1639 51146 1691
rect 50902 1565 50954 1617
rect 51574 1565 51626 1617
rect 41014 1417 41066 1469
rect 41302 1417 41354 1469
rect 35350 1343 35402 1395
rect 36310 1343 36362 1395
rect 33238 1269 33290 1321
rect 33718 1269 33770 1321
rect 36118 1269 36170 1321
rect 37270 1269 37322 1321
rect 34870 1195 34922 1247
rect 35926 1195 35978 1247
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 226 56975 254 59200
rect 214 56969 266 56975
rect 214 56911 266 56917
rect 706 56531 734 59200
rect 694 56525 746 56531
rect 694 56467 746 56473
rect 1186 55717 1214 59200
rect 1762 57049 1790 59200
rect 1750 57043 1802 57049
rect 1750 56985 1802 56991
rect 1750 56895 1802 56901
rect 1750 56837 1802 56843
rect 1174 55711 1226 55717
rect 1174 55653 1226 55659
rect 1762 17294 1790 56837
rect 2242 56531 2270 59200
rect 2614 56895 2666 56901
rect 2614 56837 2666 56843
rect 2230 56525 2282 56531
rect 2230 56467 2282 56473
rect 1846 56229 1898 56235
rect 1846 56171 1898 56177
rect 1858 38919 1886 56171
rect 1942 55415 1994 55421
rect 1942 55357 1994 55363
rect 1846 38913 1898 38919
rect 1846 38855 1898 38861
rect 1954 22861 1982 55357
rect 1942 22855 1994 22861
rect 1942 22797 1994 22803
rect 1762 17266 1886 17294
rect 1654 8277 1706 8283
rect 1654 8219 1706 8225
rect 1462 7685 1514 7691
rect 1462 7627 1514 7633
rect 1078 5687 1130 5693
rect 1078 5629 1130 5635
rect 310 5021 362 5027
rect 310 4963 362 4969
rect 118 3689 170 3695
rect 118 3631 170 3637
rect 22 3023 74 3029
rect 22 2965 74 2971
rect 34 800 62 2965
rect 130 800 158 3631
rect 214 3171 266 3177
rect 214 3113 266 3119
rect 226 800 254 3113
rect 322 800 350 4963
rect 790 4429 842 4435
rect 790 4371 842 4377
rect 502 3837 554 3843
rect 502 3779 554 3785
rect 514 800 542 3779
rect 598 3467 650 3473
rect 598 3409 650 3415
rect 610 800 638 3409
rect 694 2949 746 2955
rect 694 2891 746 2897
rect 706 800 734 2891
rect 802 800 830 4371
rect 982 3615 1034 3621
rect 982 3557 1034 3563
rect 994 800 1022 3557
rect 1090 800 1118 5629
rect 1174 4355 1226 4361
rect 1174 4297 1226 4303
rect 1186 800 1214 4297
rect 1366 4281 1418 4287
rect 1366 4223 1418 4229
rect 1378 800 1406 4223
rect 1474 3473 1502 7627
rect 1666 7214 1694 8219
rect 1858 7247 1886 17266
rect 2326 12347 2378 12353
rect 2326 12289 2378 12295
rect 2338 11909 2366 12289
rect 2326 11903 2378 11909
rect 2326 11845 2378 11851
rect 2518 11681 2570 11687
rect 2518 11623 2570 11629
rect 2134 8277 2186 8283
rect 2134 8219 2186 8225
rect 1846 7241 1898 7247
rect 1666 7186 1790 7214
rect 1654 7019 1706 7025
rect 1654 6961 1706 6967
rect 1558 6353 1610 6359
rect 1558 6295 1610 6301
rect 1462 3467 1514 3473
rect 1462 3409 1514 3415
rect 1462 3245 1514 3251
rect 1462 3187 1514 3193
rect 1474 800 1502 3187
rect 1570 800 1598 6295
rect 1666 3843 1694 6961
rect 1654 3837 1706 3843
rect 1654 3779 1706 3785
rect 1654 3689 1706 3695
rect 1654 3631 1706 3637
rect 1666 800 1694 3631
rect 1762 3177 1790 7186
rect 1846 7183 1898 7189
rect 2038 6353 2090 6359
rect 2038 6295 2090 6301
rect 1846 5021 1898 5027
rect 1846 4963 1898 4969
rect 1750 3171 1802 3177
rect 1750 3113 1802 3119
rect 1858 800 1886 4963
rect 1942 3911 1994 3917
rect 1942 3853 1994 3859
rect 1954 800 1982 3853
rect 2050 800 2078 6295
rect 2146 3251 2174 8219
rect 2530 7765 2558 11623
rect 2518 7759 2570 7765
rect 2518 7701 2570 7707
rect 2422 7463 2474 7469
rect 2422 7405 2474 7411
rect 2326 3837 2378 3843
rect 2326 3779 2378 3785
rect 2134 3245 2186 3251
rect 2134 3187 2186 3193
rect 2134 2949 2186 2955
rect 2134 2891 2186 2897
rect 2146 800 2174 2891
rect 2338 800 2366 3779
rect 2434 3621 2462 7405
rect 2518 7019 2570 7025
rect 2518 6961 2570 6967
rect 2422 3615 2474 3621
rect 2422 3557 2474 3563
rect 2422 3467 2474 3473
rect 2422 3409 2474 3415
rect 2434 800 2462 3409
rect 2530 800 2558 6961
rect 2626 5841 2654 56837
rect 2818 56531 2846 59200
rect 3298 57049 3326 59200
rect 3286 57043 3338 57049
rect 3286 56985 3338 56991
rect 3874 56531 3902 59200
rect 4354 57614 4382 59200
rect 4354 57586 4670 57614
rect 4268 57304 4564 57324
rect 4324 57302 4348 57304
rect 4404 57302 4428 57304
rect 4484 57302 4508 57304
rect 4346 57250 4348 57302
rect 4410 57250 4422 57302
rect 4484 57250 4486 57302
rect 4324 57248 4348 57250
rect 4404 57248 4428 57250
rect 4484 57248 4508 57250
rect 4268 57228 4564 57248
rect 2806 56525 2858 56531
rect 2806 56467 2858 56473
rect 3862 56525 3914 56531
rect 3862 56467 3914 56473
rect 2710 56229 2762 56235
rect 2710 56171 2762 56177
rect 2998 56229 3050 56235
rect 2998 56171 3050 56177
rect 2722 11909 2750 56171
rect 2902 36101 2954 36107
rect 2902 36043 2954 36049
rect 2710 11903 2762 11909
rect 2710 11845 2762 11851
rect 2710 8277 2762 8283
rect 2710 8219 2762 8225
rect 2614 5835 2666 5841
rect 2614 5777 2666 5783
rect 2722 3788 2750 8219
rect 2914 7913 2942 36043
rect 3010 28115 3038 56171
rect 4268 55972 4564 55992
rect 4324 55970 4348 55972
rect 4404 55970 4428 55972
rect 4484 55970 4508 55972
rect 4346 55918 4348 55970
rect 4410 55918 4422 55970
rect 4484 55918 4486 55970
rect 4324 55916 4348 55918
rect 4404 55916 4428 55918
rect 4484 55916 4508 55918
rect 4268 55896 4564 55916
rect 4642 55717 4670 57586
rect 4930 56975 4958 59200
rect 4918 56969 4970 56975
rect 4918 56911 4970 56917
rect 5410 56531 5438 59200
rect 5986 56531 6014 59200
rect 6466 56975 6494 59200
rect 6454 56969 6506 56975
rect 6454 56911 6506 56917
rect 6454 56821 6506 56827
rect 6454 56763 6506 56769
rect 5398 56525 5450 56531
rect 5398 56467 5450 56473
rect 5974 56525 6026 56531
rect 5974 56467 6026 56473
rect 5014 56229 5066 56235
rect 5014 56171 5066 56177
rect 5206 56229 5258 56235
rect 5206 56171 5258 56177
rect 6358 56229 6410 56235
rect 6358 56171 6410 56177
rect 4630 55711 4682 55717
rect 4630 55653 4682 55659
rect 4630 55563 4682 55569
rect 4630 55505 4682 55511
rect 4268 54640 4564 54660
rect 4324 54638 4348 54640
rect 4404 54638 4428 54640
rect 4484 54638 4508 54640
rect 4346 54586 4348 54638
rect 4410 54586 4422 54638
rect 4484 54586 4486 54638
rect 4324 54584 4348 54586
rect 4404 54584 4428 54586
rect 4484 54584 4508 54586
rect 4268 54564 4564 54584
rect 4268 53308 4564 53328
rect 4324 53306 4348 53308
rect 4404 53306 4428 53308
rect 4484 53306 4508 53308
rect 4346 53254 4348 53306
rect 4410 53254 4422 53306
rect 4484 53254 4486 53306
rect 4324 53252 4348 53254
rect 4404 53252 4428 53254
rect 4484 53252 4508 53254
rect 4268 53232 4564 53252
rect 4268 51976 4564 51996
rect 4324 51974 4348 51976
rect 4404 51974 4428 51976
rect 4484 51974 4508 51976
rect 4346 51922 4348 51974
rect 4410 51922 4422 51974
rect 4484 51922 4486 51974
rect 4324 51920 4348 51922
rect 4404 51920 4428 51922
rect 4484 51920 4508 51922
rect 4268 51900 4564 51920
rect 4268 50644 4564 50664
rect 4324 50642 4348 50644
rect 4404 50642 4428 50644
rect 4484 50642 4508 50644
rect 4346 50590 4348 50642
rect 4410 50590 4422 50642
rect 4484 50590 4486 50642
rect 4324 50588 4348 50590
rect 4404 50588 4428 50590
rect 4484 50588 4508 50590
rect 4268 50568 4564 50588
rect 4268 49312 4564 49332
rect 4324 49310 4348 49312
rect 4404 49310 4428 49312
rect 4484 49310 4508 49312
rect 4346 49258 4348 49310
rect 4410 49258 4422 49310
rect 4484 49258 4486 49310
rect 4324 49256 4348 49258
rect 4404 49256 4428 49258
rect 4484 49256 4508 49258
rect 4268 49236 4564 49256
rect 3574 48755 3626 48761
rect 3574 48697 3626 48703
rect 3286 35583 3338 35589
rect 3286 35525 3338 35531
rect 2998 28109 3050 28115
rect 2998 28051 3050 28057
rect 2998 11607 3050 11613
rect 2998 11549 3050 11555
rect 3010 10873 3038 11549
rect 2998 10867 3050 10873
rect 2998 10809 3050 10815
rect 3298 8431 3326 35525
rect 3586 24341 3614 48697
rect 4268 47980 4564 48000
rect 4324 47978 4348 47980
rect 4404 47978 4428 47980
rect 4484 47978 4508 47980
rect 4346 47926 4348 47978
rect 4410 47926 4422 47978
rect 4484 47926 4486 47978
rect 4324 47924 4348 47926
rect 4404 47924 4428 47926
rect 4484 47924 4508 47926
rect 4268 47904 4564 47924
rect 4268 46648 4564 46668
rect 4324 46646 4348 46648
rect 4404 46646 4428 46648
rect 4484 46646 4508 46648
rect 4346 46594 4348 46646
rect 4410 46594 4422 46646
rect 4484 46594 4486 46646
rect 4324 46592 4348 46594
rect 4404 46592 4428 46594
rect 4484 46592 4508 46594
rect 4268 46572 4564 46592
rect 4268 45316 4564 45336
rect 4324 45314 4348 45316
rect 4404 45314 4428 45316
rect 4484 45314 4508 45316
rect 4346 45262 4348 45314
rect 4410 45262 4422 45314
rect 4484 45262 4486 45314
rect 4324 45260 4348 45262
rect 4404 45260 4428 45262
rect 4484 45260 4508 45262
rect 4268 45240 4564 45260
rect 4268 43984 4564 44004
rect 4324 43982 4348 43984
rect 4404 43982 4428 43984
rect 4484 43982 4508 43984
rect 4346 43930 4348 43982
rect 4410 43930 4422 43982
rect 4484 43930 4486 43982
rect 4324 43928 4348 43930
rect 4404 43928 4428 43930
rect 4484 43928 4508 43930
rect 4268 43908 4564 43928
rect 4268 42652 4564 42672
rect 4324 42650 4348 42652
rect 4404 42650 4428 42652
rect 4484 42650 4508 42652
rect 4346 42598 4348 42650
rect 4410 42598 4422 42650
rect 4484 42598 4486 42650
rect 4324 42596 4348 42598
rect 4404 42596 4428 42598
rect 4484 42596 4508 42598
rect 4268 42576 4564 42596
rect 4268 41320 4564 41340
rect 4324 41318 4348 41320
rect 4404 41318 4428 41320
rect 4484 41318 4508 41320
rect 4346 41266 4348 41318
rect 4410 41266 4422 41318
rect 4484 41266 4486 41318
rect 4324 41264 4348 41266
rect 4404 41264 4428 41266
rect 4484 41264 4508 41266
rect 4268 41244 4564 41264
rect 4268 39988 4564 40008
rect 4324 39986 4348 39988
rect 4404 39986 4428 39988
rect 4484 39986 4508 39988
rect 4346 39934 4348 39986
rect 4410 39934 4422 39986
rect 4484 39934 4486 39986
rect 4324 39932 4348 39934
rect 4404 39932 4428 39934
rect 4484 39932 4508 39934
rect 4268 39912 4564 39932
rect 4268 38656 4564 38676
rect 4324 38654 4348 38656
rect 4404 38654 4428 38656
rect 4484 38654 4508 38656
rect 4346 38602 4348 38654
rect 4410 38602 4422 38654
rect 4484 38602 4486 38654
rect 4324 38600 4348 38602
rect 4404 38600 4428 38602
rect 4484 38600 4508 38602
rect 4268 38580 4564 38600
rect 4268 37324 4564 37344
rect 4324 37322 4348 37324
rect 4404 37322 4428 37324
rect 4484 37322 4508 37324
rect 4346 37270 4348 37322
rect 4410 37270 4422 37322
rect 4484 37270 4486 37322
rect 4324 37268 4348 37270
rect 4404 37268 4428 37270
rect 4484 37268 4508 37270
rect 4268 37248 4564 37268
rect 4268 35992 4564 36012
rect 4324 35990 4348 35992
rect 4404 35990 4428 35992
rect 4484 35990 4508 35992
rect 4346 35938 4348 35990
rect 4410 35938 4422 35990
rect 4484 35938 4486 35990
rect 4324 35936 4348 35938
rect 4404 35936 4428 35938
rect 4484 35936 4508 35938
rect 4268 35916 4564 35936
rect 4268 34660 4564 34680
rect 4324 34658 4348 34660
rect 4404 34658 4428 34660
rect 4484 34658 4508 34660
rect 4346 34606 4348 34658
rect 4410 34606 4422 34658
rect 4484 34606 4486 34658
rect 4324 34604 4348 34606
rect 4404 34604 4428 34606
rect 4484 34604 4508 34606
rect 4268 34584 4564 34604
rect 4268 33328 4564 33348
rect 4324 33326 4348 33328
rect 4404 33326 4428 33328
rect 4484 33326 4508 33328
rect 4346 33274 4348 33326
rect 4410 33274 4422 33326
rect 4484 33274 4486 33326
rect 4324 33272 4348 33274
rect 4404 33272 4428 33274
rect 4484 33272 4508 33274
rect 4268 33252 4564 33272
rect 4268 31996 4564 32016
rect 4324 31994 4348 31996
rect 4404 31994 4428 31996
rect 4484 31994 4508 31996
rect 4346 31942 4348 31994
rect 4410 31942 4422 31994
rect 4484 31942 4486 31994
rect 4324 31940 4348 31942
rect 4404 31940 4428 31942
rect 4484 31940 4508 31942
rect 4268 31920 4564 31940
rect 4268 30664 4564 30684
rect 4324 30662 4348 30664
rect 4404 30662 4428 30664
rect 4484 30662 4508 30664
rect 4346 30610 4348 30662
rect 4410 30610 4422 30662
rect 4484 30610 4486 30662
rect 4324 30608 4348 30610
rect 4404 30608 4428 30610
rect 4484 30608 4508 30610
rect 4268 30588 4564 30608
rect 4268 29332 4564 29352
rect 4324 29330 4348 29332
rect 4404 29330 4428 29332
rect 4484 29330 4508 29332
rect 4346 29278 4348 29330
rect 4410 29278 4422 29330
rect 4484 29278 4486 29330
rect 4324 29276 4348 29278
rect 4404 29276 4428 29278
rect 4484 29276 4508 29278
rect 4268 29256 4564 29276
rect 4268 28000 4564 28020
rect 4324 27998 4348 28000
rect 4404 27998 4428 28000
rect 4484 27998 4508 28000
rect 4346 27946 4348 27998
rect 4410 27946 4422 27998
rect 4484 27946 4486 27998
rect 4324 27944 4348 27946
rect 4404 27944 4428 27946
rect 4484 27944 4508 27946
rect 4268 27924 4564 27944
rect 4268 26668 4564 26688
rect 4324 26666 4348 26668
rect 4404 26666 4428 26668
rect 4484 26666 4508 26668
rect 4346 26614 4348 26666
rect 4410 26614 4422 26666
rect 4484 26614 4486 26666
rect 4324 26612 4348 26614
rect 4404 26612 4428 26614
rect 4484 26612 4508 26614
rect 4268 26592 4564 26612
rect 4268 25336 4564 25356
rect 4324 25334 4348 25336
rect 4404 25334 4428 25336
rect 4484 25334 4508 25336
rect 4346 25282 4348 25334
rect 4410 25282 4422 25334
rect 4484 25282 4486 25334
rect 4324 25280 4348 25282
rect 4404 25280 4428 25282
rect 4484 25280 4508 25282
rect 4268 25260 4564 25280
rect 3574 24335 3626 24341
rect 3574 24277 3626 24283
rect 4268 24004 4564 24024
rect 4324 24002 4348 24004
rect 4404 24002 4428 24004
rect 4484 24002 4508 24004
rect 4346 23950 4348 24002
rect 4410 23950 4422 24002
rect 4484 23950 4486 24002
rect 4324 23948 4348 23950
rect 4404 23948 4428 23950
rect 4484 23948 4508 23950
rect 4268 23928 4564 23948
rect 3670 23743 3722 23749
rect 3670 23685 3722 23691
rect 3574 21893 3626 21899
rect 3574 21835 3626 21841
rect 3586 11687 3614 21835
rect 3574 11681 3626 11687
rect 3574 11623 3626 11629
rect 3682 8579 3710 23685
rect 4268 22672 4564 22692
rect 4324 22670 4348 22672
rect 4404 22670 4428 22672
rect 4484 22670 4508 22672
rect 4346 22618 4348 22670
rect 4410 22618 4422 22670
rect 4484 22618 4486 22670
rect 4324 22616 4348 22618
rect 4404 22616 4428 22618
rect 4484 22616 4508 22618
rect 4268 22596 4564 22616
rect 4268 21340 4564 21360
rect 4324 21338 4348 21340
rect 4404 21338 4428 21340
rect 4484 21338 4508 21340
rect 4346 21286 4348 21338
rect 4410 21286 4422 21338
rect 4484 21286 4486 21338
rect 4324 21284 4348 21286
rect 4404 21284 4428 21286
rect 4484 21284 4508 21286
rect 4268 21264 4564 21284
rect 4268 20008 4564 20028
rect 4324 20006 4348 20008
rect 4404 20006 4428 20008
rect 4484 20006 4508 20008
rect 4346 19954 4348 20006
rect 4410 19954 4422 20006
rect 4484 19954 4486 20006
rect 4324 19952 4348 19954
rect 4404 19952 4428 19954
rect 4484 19952 4508 19954
rect 4268 19932 4564 19952
rect 4268 18676 4564 18696
rect 4324 18674 4348 18676
rect 4404 18674 4428 18676
rect 4484 18674 4508 18676
rect 4346 18622 4348 18674
rect 4410 18622 4422 18674
rect 4484 18622 4486 18674
rect 4324 18620 4348 18622
rect 4404 18620 4428 18622
rect 4484 18620 4508 18622
rect 4268 18600 4564 18620
rect 4268 17344 4564 17364
rect 4324 17342 4348 17344
rect 4404 17342 4428 17344
rect 4484 17342 4508 17344
rect 4346 17290 4348 17342
rect 4410 17290 4422 17342
rect 4484 17290 4486 17342
rect 4324 17288 4348 17290
rect 4404 17288 4428 17290
rect 4484 17288 4508 17290
rect 4268 17268 4564 17288
rect 4268 16012 4564 16032
rect 4324 16010 4348 16012
rect 4404 16010 4428 16012
rect 4484 16010 4508 16012
rect 4346 15958 4348 16010
rect 4410 15958 4422 16010
rect 4484 15958 4486 16010
rect 4324 15956 4348 15958
rect 4404 15956 4428 15958
rect 4484 15956 4508 15958
rect 4268 15936 4564 15956
rect 4054 14789 4106 14795
rect 4054 14731 4106 14737
rect 3670 8573 3722 8579
rect 3670 8515 3722 8521
rect 3286 8425 3338 8431
rect 3286 8367 3338 8373
rect 2998 8277 3050 8283
rect 2998 8219 3050 8225
rect 2902 7907 2954 7913
rect 2902 7849 2954 7855
rect 2902 5687 2954 5693
rect 2902 5629 2954 5635
rect 2626 3760 2750 3788
rect 2626 2881 2654 3760
rect 2710 3689 2762 3695
rect 2710 3631 2762 3637
rect 2614 2875 2666 2881
rect 2614 2817 2666 2823
rect 2722 800 2750 3631
rect 2914 2900 2942 5629
rect 2818 2872 2942 2900
rect 2818 800 2846 2872
rect 3010 2752 3038 8219
rect 4066 7765 4094 14731
rect 4268 14680 4564 14700
rect 4324 14678 4348 14680
rect 4404 14678 4428 14680
rect 4484 14678 4508 14680
rect 4346 14626 4348 14678
rect 4410 14626 4422 14678
rect 4484 14626 4486 14678
rect 4324 14624 4348 14626
rect 4404 14624 4428 14626
rect 4484 14624 4508 14626
rect 4268 14604 4564 14624
rect 4268 13348 4564 13368
rect 4324 13346 4348 13348
rect 4404 13346 4428 13348
rect 4484 13346 4508 13348
rect 4346 13294 4348 13346
rect 4410 13294 4422 13346
rect 4484 13294 4486 13346
rect 4324 13292 4348 13294
rect 4404 13292 4428 13294
rect 4484 13292 4508 13294
rect 4268 13272 4564 13292
rect 4642 12974 4670 55505
rect 5026 54829 5054 56171
rect 5014 54823 5066 54829
rect 5014 54765 5066 54771
rect 4726 48089 4778 48095
rect 4726 48031 4778 48037
rect 4738 25934 4766 48031
rect 4822 46757 4874 46763
rect 4822 46699 4874 46705
rect 4834 46541 4862 46699
rect 4822 46535 4874 46541
rect 4822 46477 4874 46483
rect 5014 37433 5066 37439
rect 5014 37375 5066 37381
rect 5026 37217 5054 37375
rect 5014 37211 5066 37217
rect 5014 37153 5066 37159
rect 4738 25906 5054 25934
rect 4642 12946 4766 12974
rect 4268 12016 4564 12036
rect 4324 12014 4348 12016
rect 4404 12014 4428 12016
rect 4484 12014 4508 12016
rect 4346 11962 4348 12014
rect 4410 11962 4422 12014
rect 4484 11962 4486 12014
rect 4324 11960 4348 11962
rect 4404 11960 4428 11962
rect 4484 11960 4508 11962
rect 4268 11940 4564 11960
rect 4268 10684 4564 10704
rect 4324 10682 4348 10684
rect 4404 10682 4428 10684
rect 4484 10682 4508 10684
rect 4346 10630 4348 10682
rect 4410 10630 4422 10682
rect 4484 10630 4486 10682
rect 4324 10628 4348 10630
rect 4404 10628 4428 10630
rect 4484 10628 4508 10630
rect 4268 10608 4564 10628
rect 4268 9352 4564 9372
rect 4324 9350 4348 9352
rect 4404 9350 4428 9352
rect 4484 9350 4508 9352
rect 4346 9298 4348 9350
rect 4410 9298 4422 9350
rect 4484 9298 4486 9350
rect 4324 9296 4348 9298
rect 4404 9296 4428 9298
rect 4484 9296 4508 9298
rect 4268 9276 4564 9296
rect 4268 8020 4564 8040
rect 4324 8018 4348 8020
rect 4404 8018 4428 8020
rect 4484 8018 4508 8020
rect 4346 7966 4348 8018
rect 4410 7966 4422 8018
rect 4484 7966 4486 8018
rect 4324 7964 4348 7966
rect 4404 7964 4428 7966
rect 4484 7964 4508 7966
rect 4268 7944 4564 7964
rect 4054 7759 4106 7765
rect 4054 7701 4106 7707
rect 3286 7463 3338 7469
rect 3286 7405 3338 7411
rect 3382 7463 3434 7469
rect 3382 7405 3434 7411
rect 4054 7463 4106 7469
rect 4054 7405 4106 7411
rect 3190 6353 3242 6359
rect 3190 6295 3242 6301
rect 3094 5021 3146 5027
rect 3094 4963 3146 4969
rect 3106 3843 3134 4963
rect 3094 3837 3146 3843
rect 3094 3779 3146 3785
rect 3094 3541 3146 3547
rect 3094 3483 3146 3489
rect 2914 2724 3038 2752
rect 2914 800 2942 2724
rect 3106 1864 3134 3483
rect 3010 1836 3134 1864
rect 3010 800 3038 1836
rect 3202 800 3230 6295
rect 3298 3917 3326 7405
rect 3286 3911 3338 3917
rect 3286 3853 3338 3859
rect 3394 3788 3422 7405
rect 3670 7019 3722 7025
rect 3670 6961 3722 6967
rect 3478 4207 3530 4213
rect 3478 4149 3530 4155
rect 3298 3760 3422 3788
rect 3298 800 3326 3760
rect 3382 3467 3434 3473
rect 3382 3409 3434 3415
rect 3394 800 3422 3409
rect 3490 800 3518 4149
rect 3682 800 3710 6961
rect 3862 6353 3914 6359
rect 3862 6295 3914 6301
rect 3766 4281 3818 4287
rect 3766 4223 3818 4229
rect 3778 800 3806 4223
rect 3874 800 3902 6295
rect 3958 4133 4010 4139
rect 3958 4075 4010 4081
rect 3970 2585 3998 4075
rect 3958 2579 4010 2585
rect 3958 2521 4010 2527
rect 4066 800 4094 7405
rect 4268 6688 4564 6708
rect 4324 6686 4348 6688
rect 4404 6686 4428 6688
rect 4484 6686 4508 6688
rect 4346 6634 4348 6686
rect 4410 6634 4422 6686
rect 4484 6634 4486 6686
rect 4324 6632 4348 6634
rect 4404 6632 4428 6634
rect 4484 6632 4508 6634
rect 4268 6612 4564 6632
rect 4630 6353 4682 6359
rect 4630 6295 4682 6301
rect 4268 5356 4564 5376
rect 4324 5354 4348 5356
rect 4404 5354 4428 5356
rect 4484 5354 4508 5356
rect 4346 5302 4348 5354
rect 4410 5302 4422 5354
rect 4484 5302 4486 5354
rect 4324 5300 4348 5302
rect 4404 5300 4428 5302
rect 4484 5300 4508 5302
rect 4268 5280 4564 5300
rect 4150 5021 4202 5027
rect 4150 4963 4202 4969
rect 4162 800 4190 4963
rect 4268 4024 4564 4044
rect 4324 4022 4348 4024
rect 4404 4022 4428 4024
rect 4484 4022 4508 4024
rect 4346 3970 4348 4022
rect 4410 3970 4422 4022
rect 4484 3970 4486 4022
rect 4324 3968 4348 3970
rect 4404 3968 4428 3970
rect 4484 3968 4508 3970
rect 4268 3948 4564 3968
rect 4268 2692 4564 2712
rect 4324 2690 4348 2692
rect 4404 2690 4428 2692
rect 4484 2690 4508 2692
rect 4346 2638 4348 2690
rect 4410 2638 4422 2690
rect 4484 2638 4486 2690
rect 4324 2636 4348 2638
rect 4404 2636 4428 2638
rect 4484 2636 4508 2638
rect 4268 2616 4564 2636
rect 4246 2579 4298 2585
rect 4246 2521 4298 2527
rect 4342 2579 4394 2585
rect 4342 2521 4394 2527
rect 4258 800 4286 2521
rect 4354 800 4382 2521
rect 4642 2456 4670 6295
rect 4738 5249 4766 12946
rect 4822 8203 4874 8209
rect 4822 8145 4874 8151
rect 4726 5243 4778 5249
rect 4726 5185 4778 5191
rect 4726 4355 4778 4361
rect 4726 4297 4778 4303
rect 4450 2428 4670 2456
rect 4450 2012 4478 2428
rect 4738 2160 4766 4297
rect 4834 2585 4862 8145
rect 4916 7798 4972 7807
rect 4916 7733 4918 7742
rect 4970 7733 4972 7742
rect 4918 7701 4970 7707
rect 5026 5767 5054 25906
rect 5218 17607 5246 56171
rect 6070 37433 6122 37439
rect 6070 37375 6122 37381
rect 5206 17601 5258 17607
rect 5206 17543 5258 17549
rect 6082 9837 6110 37375
rect 6262 29441 6314 29447
rect 6262 29383 6314 29389
rect 6070 9831 6122 9837
rect 6070 9773 6122 9779
rect 6274 9763 6302 29383
rect 6370 27005 6398 56171
rect 6466 31667 6494 56763
rect 7042 56531 7070 59200
rect 7030 56525 7082 56531
rect 7030 56467 7082 56473
rect 7522 55717 7550 59200
rect 8098 56975 8126 59200
rect 8086 56969 8138 56975
rect 8086 56911 8138 56917
rect 8278 56895 8330 56901
rect 8278 56837 8330 56843
rect 7510 55711 7562 55717
rect 7510 55653 7562 55659
rect 7318 55415 7370 55421
rect 7318 55357 7370 55363
rect 7222 49051 7274 49057
rect 7222 48993 7274 48999
rect 6454 31661 6506 31667
rect 6454 31603 6506 31609
rect 6358 26999 6410 27005
rect 6358 26941 6410 26947
rect 6838 26851 6890 26857
rect 6838 26793 6890 26799
rect 6262 9757 6314 9763
rect 6262 9699 6314 9705
rect 5686 9683 5738 9689
rect 5686 9625 5738 9631
rect 5590 8573 5642 8579
rect 5590 8515 5642 8521
rect 5602 7765 5630 8515
rect 5590 7759 5642 7765
rect 5590 7701 5642 7707
rect 5302 7463 5354 7469
rect 5302 7405 5354 7411
rect 5206 6797 5258 6803
rect 5206 6739 5258 6745
rect 5014 5761 5066 5767
rect 5014 5703 5066 5709
rect 4918 5687 4970 5693
rect 4918 5629 4970 5635
rect 5110 5687 5162 5693
rect 5110 5629 5162 5635
rect 4930 4213 4958 5629
rect 5014 4281 5066 4287
rect 5014 4223 5066 4229
rect 4918 4207 4970 4213
rect 4918 4149 4970 4155
rect 4918 3023 4970 3029
rect 4918 2965 4970 2971
rect 4822 2579 4874 2585
rect 4822 2521 4874 2527
rect 4738 2132 4862 2160
rect 4726 2061 4778 2067
rect 4450 1984 4670 2012
rect 4726 2003 4778 2009
rect 4534 1913 4586 1919
rect 4534 1855 4586 1861
rect 4546 800 4574 1855
rect 4642 800 4670 1984
rect 4738 800 4766 2003
rect 4834 1919 4862 2132
rect 4822 1913 4874 1919
rect 4822 1855 4874 1861
rect 4930 800 4958 2965
rect 5026 800 5054 4223
rect 5122 4139 5150 5629
rect 5110 4133 5162 4139
rect 5110 4075 5162 4081
rect 5218 3769 5246 6739
rect 5206 3763 5258 3769
rect 5206 3705 5258 3711
rect 5206 3023 5258 3029
rect 5206 2965 5258 2971
rect 5110 2801 5162 2807
rect 5110 2743 5162 2749
rect 5122 800 5150 2743
rect 5218 800 5246 2965
rect 5314 2067 5342 7405
rect 5698 6433 5726 9625
rect 6166 8129 6218 8135
rect 6166 8071 6218 8077
rect 5782 6945 5834 6951
rect 5782 6887 5834 6893
rect 5878 6945 5930 6951
rect 5878 6887 5930 6893
rect 5686 6427 5738 6433
rect 5686 6369 5738 6375
rect 5494 6131 5546 6137
rect 5494 6073 5546 6079
rect 5398 5021 5450 5027
rect 5398 4963 5450 4969
rect 5302 2061 5354 2067
rect 5302 2003 5354 2009
rect 5410 800 5438 4963
rect 5506 800 5534 6073
rect 5794 5915 5822 6887
rect 5782 5909 5834 5915
rect 5782 5851 5834 5857
rect 5782 5539 5834 5545
rect 5782 5481 5834 5487
rect 5686 4281 5738 4287
rect 5686 4223 5738 4229
rect 5590 3689 5642 3695
rect 5590 3631 5642 3637
rect 5602 800 5630 3631
rect 5698 800 5726 4223
rect 5794 2807 5822 5481
rect 5782 2801 5834 2807
rect 5782 2743 5834 2749
rect 5890 800 5918 6887
rect 6178 5471 6206 8071
rect 6850 7099 6878 26793
rect 7126 24187 7178 24193
rect 7126 24129 7178 24135
rect 7030 7611 7082 7617
rect 7030 7553 7082 7559
rect 6838 7093 6890 7099
rect 6838 7035 6890 7041
rect 6550 6945 6602 6951
rect 6550 6887 6602 6893
rect 6934 6945 6986 6951
rect 6934 6887 6986 6893
rect 6262 6131 6314 6137
rect 6262 6073 6314 6079
rect 6166 5465 6218 5471
rect 6166 5407 6218 5413
rect 6070 5021 6122 5027
rect 6070 4963 6122 4969
rect 5974 3023 6026 3029
rect 5974 2965 6026 2971
rect 5986 800 6014 2965
rect 6082 800 6110 4963
rect 6274 800 6302 6073
rect 6454 4207 6506 4213
rect 6454 4149 6506 4155
rect 6358 3689 6410 3695
rect 6358 3631 6410 3637
rect 6370 800 6398 3631
rect 6466 800 6494 4149
rect 6562 800 6590 6887
rect 6838 5687 6890 5693
rect 6838 5629 6890 5635
rect 6742 2949 6794 2955
rect 6742 2891 6794 2897
rect 6754 800 6782 2891
rect 6850 800 6878 5629
rect 6946 800 6974 6887
rect 7042 5767 7070 7553
rect 7138 6433 7166 24129
rect 7234 8357 7262 48993
rect 7330 14869 7358 55357
rect 8086 31661 8138 31667
rect 8086 31603 8138 31609
rect 7990 21449 8042 21455
rect 7990 21391 8042 21397
rect 8002 21104 8030 21391
rect 7954 21076 8030 21104
rect 7954 21011 7982 21076
rect 7942 21005 7994 21011
rect 7942 20947 7994 20953
rect 7942 19525 7994 19531
rect 7942 19467 7994 19473
rect 7954 19328 7982 19467
rect 7954 19300 8030 19328
rect 8002 19235 8030 19300
rect 7990 19229 8042 19235
rect 7990 19171 8042 19177
rect 7942 18193 7994 18199
rect 7942 18135 7994 18141
rect 7954 17996 7982 18135
rect 7954 17968 8030 17996
rect 8002 17681 8030 17968
rect 7990 17675 8042 17681
rect 7990 17617 8042 17623
rect 7318 14863 7370 14869
rect 7318 14805 7370 14811
rect 7604 14458 7660 14467
rect 7604 14393 7606 14402
rect 7658 14393 7660 14402
rect 7606 14361 7658 14367
rect 7798 12199 7850 12205
rect 7798 12141 7850 12147
rect 7810 11835 7838 12141
rect 7798 11829 7850 11835
rect 7798 11771 7850 11777
rect 7942 8943 7994 8949
rect 7942 8885 7994 8891
rect 7954 8843 7982 8885
rect 7940 8834 7996 8843
rect 7940 8769 7996 8778
rect 7222 8351 7274 8357
rect 7222 8293 7274 8299
rect 7702 8277 7754 8283
rect 7702 8219 7754 8225
rect 7606 8129 7658 8135
rect 7606 8071 7658 8077
rect 7618 7099 7646 8071
rect 7606 7093 7658 7099
rect 7606 7035 7658 7041
rect 7318 6871 7370 6877
rect 7318 6813 7370 6819
rect 7126 6427 7178 6433
rect 7126 6369 7178 6375
rect 7030 5761 7082 5767
rect 7030 5703 7082 5709
rect 7222 5687 7274 5693
rect 7222 5629 7274 5635
rect 7030 3689 7082 3695
rect 7030 3631 7082 3637
rect 7042 800 7070 3631
rect 7234 800 7262 5629
rect 7330 800 7358 6813
rect 7606 5539 7658 5545
rect 7606 5481 7658 5487
rect 7414 4355 7466 4361
rect 7414 4297 7466 4303
rect 7426 800 7454 4297
rect 7618 800 7646 5481
rect 7714 800 7742 8219
rect 7798 8129 7850 8135
rect 7798 8071 7850 8077
rect 7810 7839 7838 8071
rect 7940 7946 7996 7955
rect 7940 7881 7996 7890
rect 7798 7833 7850 7839
rect 7798 7775 7850 7781
rect 7954 7765 7982 7881
rect 7942 7759 7994 7765
rect 7942 7701 7994 7707
rect 7798 7241 7850 7247
rect 7798 7183 7850 7189
rect 7810 4972 7838 7183
rect 8098 6211 8126 31603
rect 8290 20956 8318 56837
rect 8578 56531 8606 59200
rect 8566 56525 8618 56531
rect 8566 56467 8618 56473
rect 8566 56229 8618 56235
rect 8566 56171 8618 56177
rect 8578 27374 8606 56171
rect 9154 55717 9182 59200
rect 9634 57049 9662 59200
rect 9622 57043 9674 57049
rect 9622 56985 9674 56991
rect 9814 56747 9866 56753
rect 9814 56689 9866 56695
rect 9142 55711 9194 55717
rect 9142 55653 9194 55659
rect 8950 55415 9002 55421
rect 8950 55357 9002 55363
rect 8482 27346 8606 27374
rect 8374 21523 8426 21529
rect 8374 21465 8426 21471
rect 8386 21085 8414 21465
rect 8374 21079 8426 21085
rect 8374 21021 8426 21027
rect 8290 20928 8414 20956
rect 8278 19821 8330 19827
rect 8278 19763 8330 19769
rect 8290 19087 8318 19763
rect 8278 19081 8330 19087
rect 8278 19023 8330 19029
rect 8386 18734 8414 20928
rect 8482 19328 8510 27346
rect 8566 22929 8618 22935
rect 8566 22871 8618 22877
rect 8578 22491 8606 22871
rect 8854 22559 8906 22565
rect 8854 22501 8906 22507
rect 8566 22485 8618 22491
rect 8566 22427 8618 22433
rect 8758 22115 8810 22121
rect 8758 22057 8810 22063
rect 8770 21696 8798 22057
rect 8674 21668 8798 21696
rect 8482 19300 8606 19328
rect 8386 18706 8510 18734
rect 8182 18489 8234 18495
rect 8182 18431 8234 18437
rect 8194 18125 8222 18431
rect 8374 18193 8426 18199
rect 8374 18135 8426 18141
rect 8182 18119 8234 18125
rect 8182 18061 8234 18067
rect 8386 17755 8414 18135
rect 8374 17749 8426 17755
rect 8374 17691 8426 17697
rect 8182 16787 8234 16793
rect 8182 16729 8234 16735
rect 8194 16423 8222 16729
rect 8182 16417 8234 16423
rect 8182 16359 8234 16365
rect 8278 16121 8330 16127
rect 8278 16063 8330 16069
rect 8182 14493 8234 14499
rect 8180 14458 8182 14467
rect 8234 14458 8236 14467
rect 8180 14393 8236 14402
rect 8182 14197 8234 14203
rect 8182 14139 8234 14145
rect 8194 13833 8222 14139
rect 8182 13827 8234 13833
rect 8182 13769 8234 13775
rect 8290 12974 8318 16063
rect 8374 15603 8426 15609
rect 8374 15545 8426 15551
rect 8386 15165 8414 15545
rect 8374 15159 8426 15165
rect 8374 15101 8426 15107
rect 8194 12946 8318 12974
rect 8194 8672 8222 12946
rect 8278 9461 8330 9467
rect 8278 9403 8330 9409
rect 8290 8843 8318 9403
rect 8276 8834 8332 8843
rect 8276 8769 8332 8778
rect 8194 8644 8414 8672
rect 8228 7650 8284 7659
rect 8228 7585 8230 7594
rect 8282 7585 8284 7594
rect 8230 7553 8282 7559
rect 8386 7099 8414 8644
rect 8374 7093 8426 7099
rect 8374 7035 8426 7041
rect 8182 6797 8234 6803
rect 8182 6739 8234 6745
rect 8086 6205 8138 6211
rect 8086 6147 8138 6153
rect 8194 4972 8222 6739
rect 8482 6304 8510 18706
rect 8578 17533 8606 19300
rect 8674 19013 8702 21668
rect 8758 21597 8810 21603
rect 8758 21539 8810 21545
rect 8770 21159 8798 21539
rect 8758 21153 8810 21159
rect 8758 21095 8810 21101
rect 8662 19007 8714 19013
rect 8662 18949 8714 18955
rect 8566 17527 8618 17533
rect 8566 17469 8618 17475
rect 8758 15455 8810 15461
rect 8758 15397 8810 15403
rect 8770 15239 8798 15397
rect 8758 15233 8810 15239
rect 8758 15175 8810 15181
rect 8566 13087 8618 13093
rect 8566 13029 8618 13035
rect 8578 8135 8606 13029
rect 8566 8129 8618 8135
rect 8566 8071 8618 8077
rect 8578 8006 8606 8071
rect 8566 7907 8618 7913
rect 8566 7849 8618 7855
rect 8578 7807 8606 7849
rect 8564 7798 8620 7807
rect 8564 7733 8620 7742
rect 8758 7463 8810 7469
rect 8758 7405 8810 7411
rect 8770 7340 8798 7405
rect 8386 6276 8510 6304
rect 8578 7312 8798 7340
rect 8386 6211 8414 6276
rect 8374 6205 8426 6211
rect 8578 6156 8606 7312
rect 8374 6147 8426 6153
rect 8482 6128 8606 6156
rect 8374 5835 8426 5841
rect 8374 5777 8426 5783
rect 7810 4953 7982 4972
rect 7810 4947 7994 4953
rect 7810 4944 7942 4947
rect 7942 4889 7994 4895
rect 8098 4944 8222 4972
rect 7894 3911 7946 3917
rect 7894 3853 7946 3859
rect 7798 3689 7850 3695
rect 7798 3631 7850 3637
rect 7810 800 7838 3631
rect 7906 800 7934 3853
rect 8098 800 8126 4944
rect 8386 4879 8414 5777
rect 8374 4873 8426 4879
rect 8374 4815 8426 4821
rect 8278 3837 8330 3843
rect 8278 3779 8330 3785
rect 8182 3023 8234 3029
rect 8182 2965 8234 2971
rect 8194 800 8222 2965
rect 8290 800 8318 3779
rect 8482 800 8510 6128
rect 8866 6008 8894 22501
rect 8962 6507 8990 55357
rect 9826 15854 9854 56689
rect 10210 56531 10238 59200
rect 10690 56531 10718 59200
rect 11266 57049 11294 59200
rect 11254 57043 11306 57049
rect 11254 56985 11306 56991
rect 11254 56895 11306 56901
rect 11254 56837 11306 56843
rect 10198 56525 10250 56531
rect 10198 56467 10250 56473
rect 10678 56525 10730 56531
rect 10678 56467 10730 56473
rect 10390 56229 10442 56235
rect 10390 56171 10442 56177
rect 10774 56229 10826 56235
rect 10774 56171 10826 56177
rect 10402 32777 10430 56171
rect 10678 38765 10730 38771
rect 10678 38707 10730 38713
rect 10582 33437 10634 33443
rect 10582 33379 10634 33385
rect 10390 32771 10442 32777
rect 10390 32713 10442 32719
rect 10006 16565 10058 16571
rect 10006 16507 10058 16513
rect 9538 15826 9854 15854
rect 9430 8351 9482 8357
rect 9430 8293 9482 8299
rect 9442 7691 9470 8293
rect 9430 7685 9482 7691
rect 9538 7659 9566 15826
rect 9910 13457 9962 13463
rect 9910 13399 9962 13405
rect 9922 13241 9950 13399
rect 9910 13235 9962 13241
rect 9910 13177 9962 13183
rect 9622 8277 9674 8283
rect 9622 8219 9674 8225
rect 9718 8277 9770 8283
rect 9718 8219 9770 8225
rect 9910 8277 9962 8283
rect 9910 8219 9962 8225
rect 9634 8135 9662 8219
rect 9622 8129 9674 8135
rect 9622 8071 9674 8077
rect 9430 7627 9482 7633
rect 9524 7650 9580 7659
rect 9524 7585 9580 7594
rect 9142 7537 9194 7543
rect 9142 7479 9194 7485
rect 8950 6501 9002 6507
rect 8950 6443 9002 6449
rect 8866 5980 8990 6008
rect 8854 5835 8906 5841
rect 8854 5777 8906 5783
rect 8758 5687 8810 5693
rect 8758 5629 8810 5635
rect 8566 3689 8618 3695
rect 8566 3631 8618 3637
rect 8578 800 8606 3631
rect 8770 2894 8798 5629
rect 8674 2866 8798 2894
rect 8674 800 8702 2866
rect 8758 2801 8810 2807
rect 8758 2743 8810 2749
rect 8770 2585 8798 2743
rect 8758 2579 8810 2585
rect 8758 2521 8810 2527
rect 8866 2456 8894 5777
rect 8962 3103 8990 5980
rect 9046 4133 9098 4139
rect 9046 4075 9098 4081
rect 8950 3097 9002 3103
rect 8950 3039 9002 3045
rect 8950 2949 9002 2955
rect 8950 2891 9002 2897
rect 8770 2428 8894 2456
rect 8770 800 8798 2428
rect 8962 800 8990 2891
rect 9058 800 9086 4075
rect 9154 800 9182 7479
rect 9430 6353 9482 6359
rect 9430 6295 9482 6301
rect 9238 5021 9290 5027
rect 9238 4963 9290 4969
rect 9250 3917 9278 4963
rect 9238 3911 9290 3917
rect 9238 3853 9290 3859
rect 9334 3689 9386 3695
rect 9334 3631 9386 3637
rect 9346 2894 9374 3631
rect 9250 2866 9374 2894
rect 9250 800 9278 2866
rect 9442 800 9470 6295
rect 9730 4417 9758 8219
rect 9814 8203 9866 8209
rect 9922 8191 9950 8219
rect 9866 8163 9950 8191
rect 9814 8145 9866 8151
rect 9910 7463 9962 7469
rect 9910 7405 9962 7411
rect 9814 6945 9866 6951
rect 9814 6887 9866 6893
rect 9826 5841 9854 6887
rect 9814 5835 9866 5841
rect 9814 5777 9866 5783
rect 9538 4389 9758 4417
rect 9538 800 9566 4389
rect 9622 4355 9674 4361
rect 9622 4297 9674 4303
rect 9634 800 9662 4297
rect 9814 4281 9866 4287
rect 9814 4223 9866 4229
rect 9826 800 9854 4223
rect 9922 800 9950 7405
rect 10018 7099 10046 16507
rect 10198 8795 10250 8801
rect 10198 8737 10250 8743
rect 10210 7765 10238 8737
rect 10594 8431 10622 33379
rect 10690 9615 10718 38707
rect 10786 25934 10814 56171
rect 10786 25906 11102 25934
rect 10870 20339 10922 20345
rect 10870 20281 10922 20287
rect 10678 9609 10730 9615
rect 10678 9551 10730 9557
rect 10582 8425 10634 8431
rect 10582 8367 10634 8373
rect 10294 8277 10346 8283
rect 10294 8219 10346 8225
rect 10582 8277 10634 8283
rect 10582 8219 10634 8225
rect 10198 7759 10250 7765
rect 10198 7701 10250 7707
rect 10006 7093 10058 7099
rect 10006 7035 10058 7041
rect 10102 6353 10154 6359
rect 10102 6295 10154 6301
rect 10006 5021 10058 5027
rect 10006 4963 10058 4969
rect 10018 3843 10046 4963
rect 10006 3837 10058 3843
rect 10006 3779 10058 3785
rect 10006 3541 10058 3547
rect 10006 3483 10058 3489
rect 10018 800 10046 3483
rect 10114 800 10142 6295
rect 10198 5687 10250 5693
rect 10198 5629 10250 5635
rect 10210 4287 10238 5629
rect 10198 4281 10250 4287
rect 10198 4223 10250 4229
rect 10306 800 10334 8219
rect 10486 5687 10538 5693
rect 10486 5629 10538 5635
rect 10390 4355 10442 4361
rect 10390 4297 10442 4303
rect 10402 800 10430 4297
rect 10498 800 10526 5629
rect 10594 800 10622 8219
rect 10882 7099 10910 20281
rect 10966 19599 11018 19605
rect 10966 19541 11018 19547
rect 10978 7765 11006 19541
rect 11074 17015 11102 25906
rect 11062 17009 11114 17015
rect 11062 16951 11114 16957
rect 11266 7839 11294 56837
rect 11746 56531 11774 59200
rect 12214 56895 12266 56901
rect 12214 56837 12266 56843
rect 11734 56525 11786 56531
rect 11734 56467 11786 56473
rect 11926 56229 11978 56235
rect 11926 56171 11978 56177
rect 11938 50907 11966 56171
rect 11926 50901 11978 50907
rect 11926 50843 11978 50849
rect 12118 44907 12170 44913
rect 12118 44849 12170 44855
rect 11446 42835 11498 42841
rect 11446 42777 11498 42783
rect 11350 42761 11402 42767
rect 11350 42703 11402 42709
rect 11362 42545 11390 42703
rect 11350 42539 11402 42545
rect 11350 42481 11402 42487
rect 11458 27374 11486 42777
rect 11362 27346 11486 27374
rect 11362 8431 11390 27346
rect 12022 18193 12074 18199
rect 12022 18135 12074 18141
rect 12034 17829 12062 18135
rect 12022 17823 12074 17829
rect 12022 17765 12074 17771
rect 12022 16861 12074 16867
rect 12022 16803 12074 16809
rect 12034 16497 12062 16803
rect 12022 16491 12074 16497
rect 12022 16433 12074 16439
rect 11446 13457 11498 13463
rect 11446 13399 11498 13405
rect 11458 10503 11486 13399
rect 11446 10497 11498 10503
rect 11446 10439 11498 10445
rect 12130 8431 12158 44849
rect 11350 8425 11402 8431
rect 11350 8367 11402 8373
rect 12118 8425 12170 8431
rect 12118 8367 12170 8373
rect 11350 8277 11402 8283
rect 11350 8219 11402 8225
rect 12118 8277 12170 8283
rect 12118 8219 12170 8225
rect 11254 7833 11306 7839
rect 11254 7775 11306 7781
rect 10966 7759 11018 7765
rect 10966 7701 11018 7707
rect 10966 7463 11018 7469
rect 10966 7405 11018 7411
rect 10870 7093 10922 7099
rect 10870 7035 10922 7041
rect 10870 6353 10922 6359
rect 10870 6295 10922 6301
rect 10678 5021 10730 5027
rect 10678 4963 10730 4969
rect 10690 4139 10718 4963
rect 10774 4355 10826 4361
rect 10774 4297 10826 4303
rect 10678 4133 10730 4139
rect 10678 4075 10730 4081
rect 10786 800 10814 4297
rect 10882 800 10910 6295
rect 10978 800 11006 7405
rect 11254 7019 11306 7025
rect 11254 6961 11306 6967
rect 11158 4207 11210 4213
rect 11158 4149 11210 4155
rect 11170 800 11198 4149
rect 11266 800 11294 6961
rect 11362 800 11390 8219
rect 11734 7537 11786 7543
rect 11734 7479 11786 7485
rect 11638 6353 11690 6359
rect 11638 6295 11690 6301
rect 11446 4133 11498 4139
rect 11446 4075 11498 4081
rect 11458 800 11486 4075
rect 11650 800 11678 6295
rect 11746 800 11774 7479
rect 11830 5021 11882 5027
rect 11830 4963 11882 4969
rect 11842 800 11870 4963
rect 12022 3245 12074 3251
rect 12022 3187 12074 3193
rect 12034 800 12062 3187
rect 12130 800 12158 8219
rect 12226 7955 12254 56837
rect 12322 56531 12350 59200
rect 12802 56975 12830 59200
rect 12790 56969 12842 56975
rect 12790 56911 12842 56917
rect 12406 56821 12458 56827
rect 12406 56763 12458 56769
rect 12310 56525 12362 56531
rect 12310 56467 12362 56473
rect 12418 47534 12446 56763
rect 13378 56531 13406 59200
rect 13366 56525 13418 56531
rect 13366 56467 13418 56473
rect 12502 56303 12554 56309
rect 12502 56245 12554 56251
rect 13750 56303 13802 56309
rect 13750 56245 13802 56251
rect 12514 51203 12542 56245
rect 12694 56229 12746 56235
rect 12694 56171 12746 56177
rect 13558 56229 13610 56235
rect 13558 56171 13610 56177
rect 12502 51197 12554 51203
rect 12502 51139 12554 51145
rect 12322 47506 12446 47534
rect 12322 10429 12350 47506
rect 12706 38253 12734 56171
rect 12694 38247 12746 38253
rect 12694 38189 12746 38195
rect 12502 36101 12554 36107
rect 12502 36043 12554 36049
rect 12406 17453 12458 17459
rect 12406 17395 12458 17401
rect 12310 10423 12362 10429
rect 12310 10365 12362 10371
rect 12212 7946 12268 7955
rect 12212 7881 12268 7890
rect 12418 7765 12446 17395
rect 12514 9171 12542 36043
rect 12598 30773 12650 30779
rect 12598 30715 12650 30721
rect 12502 9165 12554 9171
rect 12502 9107 12554 9113
rect 12610 8875 12638 30715
rect 13570 27523 13598 56171
rect 13654 43575 13706 43581
rect 13654 43517 13706 43523
rect 13558 27517 13610 27523
rect 13558 27459 13610 27465
rect 13558 22781 13610 22787
rect 13558 22723 13610 22729
rect 13570 22565 13598 22723
rect 13558 22559 13610 22565
rect 13558 22501 13610 22507
rect 13462 19007 13514 19013
rect 13462 18949 13514 18955
rect 12982 15455 13034 15461
rect 12982 15397 13034 15403
rect 12994 15239 13022 15397
rect 12982 15233 13034 15239
rect 12982 15175 13034 15181
rect 12886 13013 12938 13019
rect 12886 12955 12938 12961
rect 12598 8869 12650 8875
rect 12598 8811 12650 8817
rect 12790 8573 12842 8579
rect 12790 8515 12842 8521
rect 12406 7759 12458 7765
rect 12406 7701 12458 7707
rect 12502 7759 12554 7765
rect 12502 7701 12554 7707
rect 12310 6353 12362 6359
rect 12310 6295 12362 6301
rect 12214 3171 12266 3177
rect 12214 3113 12266 3119
rect 12226 800 12254 3113
rect 12322 800 12350 6295
rect 12514 800 12542 7701
rect 12694 7019 12746 7025
rect 12694 6961 12746 6967
rect 12598 5687 12650 5693
rect 12598 5629 12650 5635
rect 12610 800 12638 5629
rect 12706 800 12734 6961
rect 12802 800 12830 8515
rect 12898 8431 12926 12955
rect 12886 8425 12938 8431
rect 12886 8367 12938 8373
rect 13474 7099 13502 18949
rect 13666 8431 13694 43517
rect 13762 13093 13790 56245
rect 13858 55717 13886 59200
rect 14434 56975 14462 59200
rect 14422 56969 14474 56975
rect 14422 56911 14474 56917
rect 14038 56895 14090 56901
rect 14038 56837 14090 56843
rect 13846 55711 13898 55717
rect 13846 55653 13898 55659
rect 13846 38173 13898 38179
rect 13846 38115 13898 38121
rect 13750 13087 13802 13093
rect 13750 13029 13802 13035
rect 13858 9689 13886 38115
rect 13942 28923 13994 28929
rect 13942 28865 13994 28871
rect 13954 16127 13982 28865
rect 13942 16121 13994 16127
rect 13942 16063 13994 16069
rect 13846 9683 13898 9689
rect 13846 9625 13898 9631
rect 13942 9683 13994 9689
rect 13942 9625 13994 9631
rect 13654 8425 13706 8431
rect 13654 8367 13706 8373
rect 13462 7093 13514 7099
rect 13462 7035 13514 7041
rect 13462 6945 13514 6951
rect 13462 6887 13514 6893
rect 13078 6131 13130 6137
rect 13078 6073 13130 6079
rect 12982 5021 13034 5027
rect 12982 4963 13034 4969
rect 12994 3177 13022 4963
rect 12982 3171 13034 3177
rect 12982 3113 13034 3119
rect 12982 3023 13034 3029
rect 12982 2965 13034 2971
rect 12994 800 13022 2965
rect 13090 800 13118 6073
rect 13366 5687 13418 5693
rect 13366 5629 13418 5635
rect 13174 3689 13226 3695
rect 13174 3631 13226 3637
rect 13186 800 13214 3631
rect 13378 3251 13406 5629
rect 13366 3245 13418 3251
rect 13366 3187 13418 3193
rect 13366 3023 13418 3029
rect 13366 2965 13418 2971
rect 13378 800 13406 2965
rect 13474 800 13502 6887
rect 13954 6433 13982 9625
rect 13942 6427 13994 6433
rect 13942 6369 13994 6375
rect 13942 6131 13994 6137
rect 13942 6073 13994 6079
rect 13954 5120 13982 6073
rect 13858 5092 13982 5120
rect 13558 4355 13610 4361
rect 13558 4297 13610 4303
rect 13570 800 13598 4297
rect 13654 3689 13706 3695
rect 13654 3631 13706 3637
rect 13666 800 13694 3631
rect 13858 800 13886 5092
rect 13942 5021 13994 5027
rect 13942 4963 13994 4969
rect 13954 800 13982 4963
rect 14050 4435 14078 56837
rect 14914 56531 14942 59200
rect 14902 56525 14954 56531
rect 14902 56467 14954 56473
rect 15190 56229 15242 56235
rect 15190 56171 15242 56177
rect 14134 55563 14186 55569
rect 14134 55505 14186 55511
rect 14146 42323 14174 55505
rect 15094 55119 15146 55125
rect 15094 55061 15146 55067
rect 14998 52899 15050 52905
rect 14998 52841 15050 52847
rect 14134 42317 14186 42323
rect 14134 42259 14186 42265
rect 14902 36915 14954 36921
rect 14902 36857 14954 36863
rect 14914 36551 14942 36857
rect 14902 36545 14954 36551
rect 14902 36487 14954 36493
rect 14902 26777 14954 26783
rect 14902 26719 14954 26725
rect 14710 9757 14762 9763
rect 14710 9699 14762 9705
rect 14230 7611 14282 7617
rect 14230 7553 14282 7559
rect 14134 6205 14186 6211
rect 14134 6147 14186 6153
rect 14038 4429 14090 4435
rect 14038 4371 14090 4377
rect 14038 3689 14090 3695
rect 14038 3631 14090 3637
rect 14050 800 14078 3631
rect 14146 800 14174 6147
rect 14242 2881 14270 7553
rect 14614 6945 14666 6951
rect 14614 6887 14666 6893
rect 14422 5021 14474 5027
rect 14422 4963 14474 4969
rect 14434 2900 14462 4963
rect 14518 3023 14570 3029
rect 14518 2965 14570 2971
rect 14230 2875 14282 2881
rect 14230 2817 14282 2823
rect 14338 2872 14462 2900
rect 14338 800 14366 2872
rect 14530 1568 14558 2965
rect 14434 1540 14558 1568
rect 14434 800 14462 1540
rect 14626 1420 14654 6887
rect 14722 6433 14750 9699
rect 14914 8801 14942 26719
rect 14902 8795 14954 8801
rect 14902 8737 14954 8743
rect 15010 7099 15038 52841
rect 14998 7093 15050 7099
rect 14998 7035 15050 7041
rect 15106 6581 15134 55061
rect 15202 9023 15230 56171
rect 15394 56161 15422 59200
rect 15970 56975 15998 59200
rect 16450 57049 16478 59200
rect 16438 57043 16490 57049
rect 16438 56985 16490 56991
rect 15958 56969 16010 56975
rect 15958 56911 16010 56917
rect 16150 56895 16202 56901
rect 16150 56837 16202 56843
rect 15382 56155 15434 56161
rect 15382 56097 15434 56103
rect 15286 54749 15338 54755
rect 15286 54691 15338 54697
rect 15298 24267 15326 54691
rect 16054 26777 16106 26783
rect 16054 26719 16106 26725
rect 15286 24261 15338 24267
rect 15286 24203 15338 24209
rect 15958 23817 16010 23823
rect 15958 23759 16010 23765
rect 15862 9831 15914 9837
rect 15862 9773 15914 9779
rect 15190 9017 15242 9023
rect 15190 8959 15242 8965
rect 15670 7463 15722 7469
rect 15670 7405 15722 7411
rect 15382 6945 15434 6951
rect 15382 6887 15434 6893
rect 15094 6575 15146 6581
rect 15094 6517 15146 6523
rect 14710 6427 14762 6433
rect 14710 6369 14762 6375
rect 14902 6353 14954 6359
rect 14902 6295 14954 6301
rect 14806 5021 14858 5027
rect 14530 1392 14654 1420
rect 14722 4981 14806 5009
rect 14530 800 14558 1392
rect 14722 800 14750 4981
rect 14806 4963 14858 4969
rect 14806 3689 14858 3695
rect 14806 3631 14858 3637
rect 14818 800 14846 3631
rect 14914 800 14942 6295
rect 14998 5687 15050 5693
rect 14998 5629 15050 5635
rect 15010 800 15038 5629
rect 15286 3689 15338 3695
rect 15202 3649 15286 3677
rect 15202 800 15230 3649
rect 15286 3631 15338 3637
rect 15394 3492 15422 6887
rect 15478 4355 15530 4361
rect 15478 4297 15530 4303
rect 15298 3464 15422 3492
rect 15298 800 15326 3464
rect 15382 2949 15434 2955
rect 15382 2891 15434 2897
rect 15394 800 15422 2891
rect 15490 800 15518 4297
rect 15682 800 15710 7405
rect 15874 6581 15902 9773
rect 15970 7765 15998 23759
rect 15958 7759 16010 7765
rect 15958 7701 16010 7707
rect 15958 7611 16010 7617
rect 15958 7553 16010 7559
rect 15970 7025 15998 7553
rect 16066 7099 16094 26719
rect 16162 9467 16190 56837
rect 17026 56531 17054 59200
rect 17506 56975 17534 59200
rect 18082 57049 18110 59200
rect 18562 57614 18590 59200
rect 18562 57586 18782 57614
rect 18070 57043 18122 57049
rect 18070 56985 18122 56991
rect 17494 56969 17546 56975
rect 17494 56911 17546 56917
rect 18754 56531 18782 57586
rect 19138 56975 19166 59200
rect 19618 57614 19646 59200
rect 19618 57586 20030 57614
rect 19126 56969 19178 56975
rect 19126 56911 19178 56917
rect 19628 56638 19924 56658
rect 19684 56636 19708 56638
rect 19764 56636 19788 56638
rect 19844 56636 19868 56638
rect 19706 56584 19708 56636
rect 19770 56584 19782 56636
rect 19844 56584 19846 56636
rect 19684 56582 19708 56584
rect 19764 56582 19788 56584
rect 19844 56582 19868 56584
rect 19628 56562 19924 56582
rect 20002 56531 20030 57586
rect 17014 56525 17066 56531
rect 17014 56467 17066 56473
rect 18742 56525 18794 56531
rect 18742 56467 18794 56473
rect 19990 56525 20042 56531
rect 19990 56467 20042 56473
rect 16822 56229 16874 56235
rect 16822 56171 16874 56177
rect 18646 56229 18698 56235
rect 18646 56171 18698 56177
rect 16630 46831 16682 46837
rect 16630 46773 16682 46779
rect 16534 42243 16586 42249
rect 16534 42185 16586 42191
rect 16546 22417 16574 42185
rect 16642 25229 16670 46773
rect 16834 26931 16862 56171
rect 17398 55415 17450 55421
rect 17398 55357 17450 55363
rect 16822 26925 16874 26931
rect 16822 26867 16874 26873
rect 16630 25223 16682 25229
rect 16630 25165 16682 25171
rect 17410 23897 17438 55357
rect 17974 44093 18026 44099
rect 17974 44035 18026 44041
rect 17878 36101 17930 36107
rect 17878 36043 17930 36049
rect 17398 23891 17450 23897
rect 17398 23833 17450 23839
rect 17782 22781 17834 22787
rect 17782 22723 17834 22729
rect 16534 22411 16586 22417
rect 16534 22353 16586 22359
rect 17794 19753 17822 22723
rect 17782 19747 17834 19753
rect 17782 19689 17834 19695
rect 17302 18267 17354 18273
rect 17302 18209 17354 18215
rect 16630 15899 16682 15905
rect 16630 15841 16682 15847
rect 16150 9461 16202 9467
rect 16150 9403 16202 9409
rect 16246 9461 16298 9467
rect 16246 9403 16298 9409
rect 16258 8357 16286 9403
rect 16246 8351 16298 8357
rect 16246 8293 16298 8299
rect 16150 8277 16202 8283
rect 16150 8219 16202 8225
rect 16342 8277 16394 8283
rect 16342 8219 16394 8225
rect 16054 7093 16106 7099
rect 16054 7035 16106 7041
rect 15958 7019 16010 7025
rect 15958 6961 16010 6967
rect 15862 6575 15914 6581
rect 15862 6517 15914 6523
rect 15862 5687 15914 5693
rect 15862 5629 15914 5635
rect 15874 2900 15902 5629
rect 15958 4355 16010 4361
rect 15958 4297 16010 4303
rect 15778 2872 15902 2900
rect 15778 800 15806 2872
rect 15970 2160 15998 4297
rect 16162 3640 16190 8219
rect 16246 5687 16298 5693
rect 16246 5629 16298 5635
rect 15874 2132 15998 2160
rect 16066 3612 16190 3640
rect 15874 800 15902 2132
rect 16066 800 16094 3612
rect 16258 2900 16286 5629
rect 16162 2872 16286 2900
rect 16162 800 16190 2872
rect 16246 2209 16298 2215
rect 16246 2151 16298 2157
rect 16258 800 16286 2151
rect 16354 800 16382 8219
rect 16642 7099 16670 15841
rect 17014 11015 17066 11021
rect 17014 10957 17066 10963
rect 17026 8357 17054 10957
rect 17014 8351 17066 8357
rect 17014 8293 17066 8299
rect 17110 8351 17162 8357
rect 17110 8293 17162 8299
rect 17122 7839 17150 8293
rect 17110 7833 17162 7839
rect 17110 7775 17162 7781
rect 17314 7099 17342 18209
rect 17590 10275 17642 10281
rect 17590 10217 17642 10223
rect 16630 7093 16682 7099
rect 16630 7035 16682 7041
rect 17302 7093 17354 7099
rect 17302 7035 17354 7041
rect 17110 6945 17162 6951
rect 17110 6887 17162 6893
rect 16822 6205 16874 6211
rect 16822 6147 16874 6153
rect 16534 5021 16586 5027
rect 16534 4963 16586 4969
rect 16438 4355 16490 4361
rect 16438 4297 16490 4303
rect 16450 2215 16478 4297
rect 16546 2955 16574 4963
rect 16726 3837 16778 3843
rect 16726 3779 16778 3785
rect 16630 3023 16682 3029
rect 16630 2965 16682 2971
rect 16534 2949 16586 2955
rect 16534 2891 16586 2897
rect 16438 2209 16490 2215
rect 16438 2151 16490 2157
rect 16534 1987 16586 1993
rect 16534 1929 16586 1935
rect 16546 800 16574 1929
rect 16642 800 16670 2965
rect 16738 1993 16766 3779
rect 16726 1987 16778 1993
rect 16726 1929 16778 1935
rect 16834 1864 16862 6147
rect 16918 4281 16970 4287
rect 16918 4223 16970 4229
rect 16738 1836 16862 1864
rect 16738 800 16766 1836
rect 16930 800 16958 4223
rect 17014 3023 17066 3029
rect 17014 2965 17066 2971
rect 17026 800 17054 2965
rect 17122 800 17150 6887
rect 17602 5915 17630 10217
rect 17686 9535 17738 9541
rect 17686 9477 17738 9483
rect 17698 6433 17726 9477
rect 17782 8129 17834 8135
rect 17782 8071 17834 8077
rect 17686 6427 17738 6433
rect 17686 6369 17738 6375
rect 17590 5909 17642 5915
rect 17590 5851 17642 5857
rect 17302 5687 17354 5693
rect 17302 5629 17354 5635
rect 17314 3843 17342 5629
rect 17794 5471 17822 8071
rect 17890 7173 17918 36043
rect 17986 20345 18014 44035
rect 18454 36767 18506 36773
rect 18454 36709 18506 36715
rect 17974 20339 18026 20345
rect 17974 20281 18026 20287
rect 17878 7167 17930 7173
rect 17878 7109 17930 7115
rect 17878 6945 17930 6951
rect 17878 6887 17930 6893
rect 17782 5465 17834 5471
rect 17782 5407 17834 5413
rect 17494 5021 17546 5027
rect 17494 4963 17546 4969
rect 17302 3837 17354 3843
rect 17302 3779 17354 3785
rect 17398 3689 17450 3695
rect 17398 3631 17450 3637
rect 17302 3541 17354 3547
rect 17302 3483 17354 3489
rect 17314 2900 17342 3483
rect 17218 2872 17342 2900
rect 17218 800 17246 2872
rect 17410 800 17438 3631
rect 17506 3547 17534 4963
rect 17590 4281 17642 4287
rect 17590 4223 17642 4229
rect 17494 3541 17546 3547
rect 17494 3483 17546 3489
rect 17494 3245 17546 3251
rect 17494 3187 17546 3193
rect 17506 800 17534 3187
rect 17602 800 17630 4223
rect 17686 2949 17738 2955
rect 17686 2891 17738 2897
rect 17698 800 17726 2891
rect 17890 800 17918 6887
rect 18466 6433 18494 36709
rect 18658 36181 18686 56171
rect 20194 55717 20222 59200
rect 20674 56975 20702 59200
rect 20662 56969 20714 56975
rect 20662 56911 20714 56917
rect 21250 56531 21278 59200
rect 21622 56895 21674 56901
rect 21622 56837 21674 56843
rect 21238 56525 21290 56531
rect 21238 56467 21290 56473
rect 20854 56229 20906 56235
rect 20854 56171 20906 56177
rect 21430 56229 21482 56235
rect 21430 56171 21482 56177
rect 20182 55711 20234 55717
rect 20182 55653 20234 55659
rect 20566 55637 20618 55643
rect 20566 55579 20618 55585
rect 20086 55415 20138 55421
rect 20086 55357 20138 55363
rect 19628 55306 19924 55326
rect 19684 55304 19708 55306
rect 19764 55304 19788 55306
rect 19844 55304 19868 55306
rect 19706 55252 19708 55304
rect 19770 55252 19782 55304
rect 19844 55252 19846 55304
rect 19684 55250 19708 55252
rect 19764 55250 19788 55252
rect 19844 55250 19868 55252
rect 19628 55230 19924 55250
rect 19628 53974 19924 53994
rect 19684 53972 19708 53974
rect 19764 53972 19788 53974
rect 19844 53972 19868 53974
rect 19706 53920 19708 53972
rect 19770 53920 19782 53972
rect 19844 53920 19846 53972
rect 19684 53918 19708 53920
rect 19764 53918 19788 53920
rect 19844 53918 19868 53920
rect 19628 53898 19924 53918
rect 19628 52642 19924 52662
rect 19684 52640 19708 52642
rect 19764 52640 19788 52642
rect 19844 52640 19868 52642
rect 19706 52588 19708 52640
rect 19770 52588 19782 52640
rect 19844 52588 19846 52640
rect 19684 52586 19708 52588
rect 19764 52586 19788 52588
rect 19844 52586 19868 52588
rect 19628 52566 19924 52586
rect 19414 51567 19466 51573
rect 19414 51509 19466 51515
rect 18646 36175 18698 36181
rect 18646 36117 18698 36123
rect 19030 30773 19082 30779
rect 19030 30715 19082 30721
rect 19042 30483 19070 30715
rect 19030 30477 19082 30483
rect 19030 30419 19082 30425
rect 19426 26117 19454 51509
rect 19628 51310 19924 51330
rect 19684 51308 19708 51310
rect 19764 51308 19788 51310
rect 19844 51308 19868 51310
rect 19706 51256 19708 51308
rect 19770 51256 19782 51308
rect 19844 51256 19846 51308
rect 19684 51254 19708 51256
rect 19764 51254 19788 51256
rect 19844 51254 19868 51256
rect 19628 51234 19924 51254
rect 19628 49978 19924 49998
rect 19684 49976 19708 49978
rect 19764 49976 19788 49978
rect 19844 49976 19868 49978
rect 19706 49924 19708 49976
rect 19770 49924 19782 49976
rect 19844 49924 19846 49976
rect 19684 49922 19708 49924
rect 19764 49922 19788 49924
rect 19844 49922 19868 49924
rect 19628 49902 19924 49922
rect 19628 48646 19924 48666
rect 19684 48644 19708 48646
rect 19764 48644 19788 48646
rect 19844 48644 19868 48646
rect 19706 48592 19708 48644
rect 19770 48592 19782 48644
rect 19844 48592 19846 48644
rect 19684 48590 19708 48592
rect 19764 48590 19788 48592
rect 19844 48590 19868 48592
rect 19628 48570 19924 48590
rect 19628 47314 19924 47334
rect 19684 47312 19708 47314
rect 19764 47312 19788 47314
rect 19844 47312 19868 47314
rect 19706 47260 19708 47312
rect 19770 47260 19782 47312
rect 19844 47260 19846 47312
rect 19684 47258 19708 47260
rect 19764 47258 19788 47260
rect 19844 47258 19868 47260
rect 19628 47238 19924 47258
rect 19990 46757 20042 46763
rect 19990 46699 20042 46705
rect 19628 45982 19924 46002
rect 19684 45980 19708 45982
rect 19764 45980 19788 45982
rect 19844 45980 19868 45982
rect 19706 45928 19708 45980
rect 19770 45928 19782 45980
rect 19844 45928 19846 45980
rect 19684 45926 19708 45928
rect 19764 45926 19788 45928
rect 19844 45926 19868 45928
rect 19628 45906 19924 45926
rect 19628 44650 19924 44670
rect 19684 44648 19708 44650
rect 19764 44648 19788 44650
rect 19844 44648 19868 44650
rect 19706 44596 19708 44648
rect 19770 44596 19782 44648
rect 19844 44596 19846 44648
rect 19684 44594 19708 44596
rect 19764 44594 19788 44596
rect 19844 44594 19868 44596
rect 19628 44574 19924 44594
rect 19628 43318 19924 43338
rect 19684 43316 19708 43318
rect 19764 43316 19788 43318
rect 19844 43316 19868 43318
rect 19706 43264 19708 43316
rect 19770 43264 19782 43316
rect 19844 43264 19846 43316
rect 19684 43262 19708 43264
rect 19764 43262 19788 43264
rect 19844 43262 19868 43264
rect 19628 43242 19924 43262
rect 19628 41986 19924 42006
rect 19684 41984 19708 41986
rect 19764 41984 19788 41986
rect 19844 41984 19868 41986
rect 19706 41932 19708 41984
rect 19770 41932 19782 41984
rect 19844 41932 19846 41984
rect 19684 41930 19708 41932
rect 19764 41930 19788 41932
rect 19844 41930 19868 41932
rect 19628 41910 19924 41930
rect 19628 40654 19924 40674
rect 19684 40652 19708 40654
rect 19764 40652 19788 40654
rect 19844 40652 19868 40654
rect 19706 40600 19708 40652
rect 19770 40600 19782 40652
rect 19844 40600 19846 40652
rect 19684 40598 19708 40600
rect 19764 40598 19788 40600
rect 19844 40598 19868 40600
rect 19628 40578 19924 40598
rect 19628 39322 19924 39342
rect 19684 39320 19708 39322
rect 19764 39320 19788 39322
rect 19844 39320 19868 39322
rect 19706 39268 19708 39320
rect 19770 39268 19782 39320
rect 19844 39268 19846 39320
rect 19684 39266 19708 39268
rect 19764 39266 19788 39268
rect 19844 39266 19868 39268
rect 19628 39246 19924 39266
rect 19628 37990 19924 38010
rect 19684 37988 19708 37990
rect 19764 37988 19788 37990
rect 19844 37988 19868 37990
rect 19706 37936 19708 37988
rect 19770 37936 19782 37988
rect 19844 37936 19846 37988
rect 19684 37934 19708 37936
rect 19764 37934 19788 37936
rect 19844 37934 19868 37936
rect 19628 37914 19924 37934
rect 19628 36658 19924 36678
rect 19684 36656 19708 36658
rect 19764 36656 19788 36658
rect 19844 36656 19868 36658
rect 19706 36604 19708 36656
rect 19770 36604 19782 36656
rect 19844 36604 19846 36656
rect 19684 36602 19708 36604
rect 19764 36602 19788 36604
rect 19844 36602 19868 36604
rect 19628 36582 19924 36602
rect 19510 36249 19562 36255
rect 19510 36191 19562 36197
rect 19414 26111 19466 26117
rect 19414 26053 19466 26059
rect 19522 22343 19550 36191
rect 19628 35326 19924 35346
rect 19684 35324 19708 35326
rect 19764 35324 19788 35326
rect 19844 35324 19868 35326
rect 19706 35272 19708 35324
rect 19770 35272 19782 35324
rect 19844 35272 19846 35324
rect 19684 35270 19708 35272
rect 19764 35270 19788 35272
rect 19844 35270 19868 35272
rect 19628 35250 19924 35270
rect 19628 33994 19924 34014
rect 19684 33992 19708 33994
rect 19764 33992 19788 33994
rect 19844 33992 19868 33994
rect 19706 33940 19708 33992
rect 19770 33940 19782 33992
rect 19844 33940 19846 33992
rect 19684 33938 19708 33940
rect 19764 33938 19788 33940
rect 19844 33938 19868 33940
rect 19628 33918 19924 33938
rect 19628 32662 19924 32682
rect 19684 32660 19708 32662
rect 19764 32660 19788 32662
rect 19844 32660 19868 32662
rect 19706 32608 19708 32660
rect 19770 32608 19782 32660
rect 19844 32608 19846 32660
rect 19684 32606 19708 32608
rect 19764 32606 19788 32608
rect 19844 32606 19868 32608
rect 19628 32586 19924 32606
rect 19628 31330 19924 31350
rect 19684 31328 19708 31330
rect 19764 31328 19788 31330
rect 19844 31328 19868 31330
rect 19706 31276 19708 31328
rect 19770 31276 19782 31328
rect 19844 31276 19846 31328
rect 19684 31274 19708 31276
rect 19764 31274 19788 31276
rect 19844 31274 19868 31276
rect 19628 31254 19924 31274
rect 19628 29998 19924 30018
rect 19684 29996 19708 29998
rect 19764 29996 19788 29998
rect 19844 29996 19868 29998
rect 19706 29944 19708 29996
rect 19770 29944 19782 29996
rect 19844 29944 19846 29996
rect 19684 29942 19708 29944
rect 19764 29942 19788 29944
rect 19844 29942 19868 29944
rect 19628 29922 19924 29942
rect 19628 28666 19924 28686
rect 19684 28664 19708 28666
rect 19764 28664 19788 28666
rect 19844 28664 19868 28666
rect 19706 28612 19708 28664
rect 19770 28612 19782 28664
rect 19844 28612 19846 28664
rect 19684 28610 19708 28612
rect 19764 28610 19788 28612
rect 19844 28610 19868 28612
rect 19628 28590 19924 28610
rect 19628 27334 19924 27354
rect 19684 27332 19708 27334
rect 19764 27332 19788 27334
rect 19844 27332 19868 27334
rect 19706 27280 19708 27332
rect 19770 27280 19782 27332
rect 19844 27280 19846 27332
rect 19684 27278 19708 27280
rect 19764 27278 19788 27280
rect 19844 27278 19868 27280
rect 19628 27258 19924 27278
rect 19628 26002 19924 26022
rect 19684 26000 19708 26002
rect 19764 26000 19788 26002
rect 19844 26000 19868 26002
rect 19706 25948 19708 26000
rect 19770 25948 19782 26000
rect 19844 25948 19846 26000
rect 19684 25946 19708 25948
rect 19764 25946 19788 25948
rect 19844 25946 19868 25948
rect 19628 25926 19924 25946
rect 19628 24670 19924 24690
rect 19684 24668 19708 24670
rect 19764 24668 19788 24670
rect 19844 24668 19868 24670
rect 19706 24616 19708 24668
rect 19770 24616 19782 24668
rect 19844 24616 19846 24668
rect 19684 24614 19708 24616
rect 19764 24614 19788 24616
rect 19844 24614 19868 24616
rect 19628 24594 19924 24614
rect 19628 23338 19924 23358
rect 19684 23336 19708 23338
rect 19764 23336 19788 23338
rect 19844 23336 19868 23338
rect 19706 23284 19708 23336
rect 19770 23284 19782 23336
rect 19844 23284 19846 23336
rect 19684 23282 19708 23284
rect 19764 23282 19788 23284
rect 19844 23282 19868 23284
rect 19628 23262 19924 23282
rect 19510 22337 19562 22343
rect 19510 22279 19562 22285
rect 19628 22006 19924 22026
rect 19684 22004 19708 22006
rect 19764 22004 19788 22006
rect 19844 22004 19868 22006
rect 19706 21952 19708 22004
rect 19770 21952 19782 22004
rect 19844 21952 19846 22004
rect 19684 21950 19708 21952
rect 19764 21950 19788 21952
rect 19844 21950 19868 21952
rect 19628 21930 19924 21950
rect 19628 20674 19924 20694
rect 19684 20672 19708 20674
rect 19764 20672 19788 20674
rect 19844 20672 19868 20674
rect 19706 20620 19708 20672
rect 19770 20620 19782 20672
rect 19844 20620 19846 20672
rect 19684 20618 19708 20620
rect 19764 20618 19788 20620
rect 19844 20618 19868 20620
rect 19628 20598 19924 20618
rect 19628 19342 19924 19362
rect 19684 19340 19708 19342
rect 19764 19340 19788 19342
rect 19844 19340 19868 19342
rect 19706 19288 19708 19340
rect 19770 19288 19782 19340
rect 19844 19288 19846 19340
rect 19684 19286 19708 19288
rect 19764 19286 19788 19288
rect 19844 19286 19868 19288
rect 19628 19266 19924 19286
rect 19628 18010 19924 18030
rect 19684 18008 19708 18010
rect 19764 18008 19788 18010
rect 19844 18008 19868 18010
rect 19706 17956 19708 18008
rect 19770 17956 19782 18008
rect 19844 17956 19846 18008
rect 19684 17954 19708 17956
rect 19764 17954 19788 17956
rect 19844 17954 19868 17956
rect 19628 17934 19924 17954
rect 19628 16678 19924 16698
rect 19684 16676 19708 16678
rect 19764 16676 19788 16678
rect 19844 16676 19868 16678
rect 19706 16624 19708 16676
rect 19770 16624 19782 16676
rect 19844 16624 19846 16676
rect 19684 16622 19708 16624
rect 19764 16622 19788 16624
rect 19844 16622 19868 16624
rect 19628 16602 19924 16622
rect 19628 15346 19924 15366
rect 19684 15344 19708 15346
rect 19764 15344 19788 15346
rect 19844 15344 19868 15346
rect 19706 15292 19708 15344
rect 19770 15292 19782 15344
rect 19844 15292 19846 15344
rect 19684 15290 19708 15292
rect 19764 15290 19788 15292
rect 19844 15290 19868 15292
rect 19628 15270 19924 15290
rect 19628 14014 19924 14034
rect 19684 14012 19708 14014
rect 19764 14012 19788 14014
rect 19844 14012 19868 14014
rect 19706 13960 19708 14012
rect 19770 13960 19782 14012
rect 19844 13960 19846 14012
rect 19684 13958 19708 13960
rect 19764 13958 19788 13960
rect 19844 13958 19868 13960
rect 19628 13938 19924 13958
rect 19628 12682 19924 12702
rect 19684 12680 19708 12682
rect 19764 12680 19788 12682
rect 19844 12680 19868 12682
rect 19706 12628 19708 12680
rect 19770 12628 19782 12680
rect 19844 12628 19846 12680
rect 19684 12626 19708 12628
rect 19764 12626 19788 12628
rect 19844 12626 19868 12628
rect 19628 12606 19924 12626
rect 19628 11350 19924 11370
rect 19684 11348 19708 11350
rect 19764 11348 19788 11350
rect 19844 11348 19868 11350
rect 19706 11296 19708 11348
rect 19770 11296 19782 11348
rect 19844 11296 19846 11348
rect 19684 11294 19708 11296
rect 19764 11294 19788 11296
rect 19844 11294 19868 11296
rect 19628 11274 19924 11294
rect 19628 10018 19924 10038
rect 19684 10016 19708 10018
rect 19764 10016 19788 10018
rect 19844 10016 19868 10018
rect 19706 9964 19708 10016
rect 19770 9964 19782 10016
rect 19844 9964 19846 10016
rect 19684 9962 19708 9964
rect 19764 9962 19788 9964
rect 19844 9962 19868 9964
rect 19628 9942 19924 9962
rect 19222 9757 19274 9763
rect 19222 9699 19274 9705
rect 18838 8795 18890 8801
rect 18838 8737 18890 8743
rect 18850 7099 18878 8737
rect 18838 7093 18890 7099
rect 18838 7035 18890 7041
rect 18550 6945 18602 6951
rect 18550 6887 18602 6893
rect 18454 6427 18506 6433
rect 18454 6369 18506 6375
rect 18262 6205 18314 6211
rect 18262 6147 18314 6153
rect 17974 5021 18026 5027
rect 17974 4963 18026 4969
rect 17986 800 18014 4963
rect 18070 3689 18122 3695
rect 18070 3631 18122 3637
rect 18082 800 18110 3631
rect 18274 800 18302 6147
rect 18358 6131 18410 6137
rect 18358 6073 18410 6079
rect 18370 3251 18398 6073
rect 18454 3689 18506 3695
rect 18454 3631 18506 3637
rect 18358 3245 18410 3251
rect 18358 3187 18410 3193
rect 18358 3097 18410 3103
rect 18358 3039 18410 3045
rect 18370 800 18398 3039
rect 18466 800 18494 3631
rect 18562 800 18590 6887
rect 19234 6433 19262 9699
rect 19628 8686 19924 8706
rect 19684 8684 19708 8686
rect 19764 8684 19788 8686
rect 19844 8684 19868 8686
rect 19706 8632 19708 8684
rect 19770 8632 19782 8684
rect 19844 8632 19846 8684
rect 19684 8630 19708 8632
rect 19764 8630 19788 8632
rect 19844 8630 19868 8632
rect 19628 8610 19924 8630
rect 19628 7354 19924 7374
rect 19684 7352 19708 7354
rect 19764 7352 19788 7354
rect 19844 7352 19868 7354
rect 19706 7300 19708 7352
rect 19770 7300 19782 7352
rect 19844 7300 19846 7352
rect 19684 7298 19708 7300
rect 19764 7298 19788 7300
rect 19844 7298 19868 7300
rect 19628 7278 19924 7298
rect 20002 7173 20030 46699
rect 20098 15905 20126 55357
rect 20470 54749 20522 54755
rect 20470 54691 20522 54697
rect 20482 45431 20510 54691
rect 20470 45425 20522 45431
rect 20470 45367 20522 45373
rect 20086 15899 20138 15905
rect 20086 15841 20138 15847
rect 20470 14789 20522 14795
rect 20470 14731 20522 14737
rect 20278 12569 20330 12575
rect 20278 12511 20330 12517
rect 20290 9467 20318 12511
rect 20374 12125 20426 12131
rect 20374 12067 20426 12073
rect 20386 11835 20414 12067
rect 20374 11829 20426 11835
rect 20374 11771 20426 11777
rect 20278 9461 20330 9467
rect 20278 9403 20330 9409
rect 19990 7167 20042 7173
rect 19990 7109 20042 7115
rect 20374 6945 20426 6951
rect 20374 6887 20426 6893
rect 19222 6427 19274 6433
rect 19222 6369 19274 6375
rect 19318 6353 19370 6359
rect 19318 6295 19370 6301
rect 18934 6205 18986 6211
rect 18934 6147 18986 6153
rect 18742 5687 18794 5693
rect 18742 5629 18794 5635
rect 18754 800 18782 5629
rect 18838 3023 18890 3029
rect 18838 2965 18890 2971
rect 18850 800 18878 2965
rect 18946 800 18974 6147
rect 19030 5021 19082 5027
rect 19030 4963 19082 4969
rect 19126 5021 19178 5027
rect 19126 4963 19178 4969
rect 19042 3103 19070 4963
rect 19030 3097 19082 3103
rect 19030 3039 19082 3045
rect 19138 2604 19166 4963
rect 19222 3689 19274 3695
rect 19222 3631 19274 3637
rect 19042 2576 19166 2604
rect 19042 800 19070 2576
rect 19234 800 19262 3631
rect 19330 800 19358 6295
rect 19628 6022 19924 6042
rect 19684 6020 19708 6022
rect 19764 6020 19788 6022
rect 19844 6020 19868 6022
rect 19706 5968 19708 6020
rect 19770 5968 19782 6020
rect 19844 5968 19846 6020
rect 19684 5966 19708 5968
rect 19764 5966 19788 5968
rect 19844 5966 19868 5968
rect 19628 5946 19924 5966
rect 20182 5687 20234 5693
rect 20182 5629 20234 5635
rect 19628 4690 19924 4710
rect 19684 4688 19708 4690
rect 19764 4688 19788 4690
rect 19844 4688 19868 4690
rect 19706 4636 19708 4688
rect 19770 4636 19782 4688
rect 19844 4636 19846 4688
rect 19684 4634 19708 4636
rect 19764 4634 19788 4636
rect 19844 4634 19868 4636
rect 19628 4614 19924 4634
rect 19414 3837 19466 3843
rect 19414 3779 19466 3785
rect 19426 800 19454 3779
rect 19990 3689 20042 3695
rect 19990 3631 20042 3637
rect 19628 3358 19924 3378
rect 19684 3356 19708 3358
rect 19764 3356 19788 3358
rect 19844 3356 19868 3358
rect 19706 3304 19708 3356
rect 19770 3304 19782 3356
rect 19844 3304 19846 3356
rect 19684 3302 19708 3304
rect 19764 3302 19788 3304
rect 19844 3302 19868 3304
rect 19628 3282 19924 3302
rect 19702 3245 19754 3251
rect 19702 3187 19754 3193
rect 19606 2949 19658 2955
rect 19606 2891 19658 2897
rect 19618 800 19646 2891
rect 19714 800 19742 3187
rect 19798 3097 19850 3103
rect 19798 3039 19850 3045
rect 19810 800 19838 3039
rect 20002 1864 20030 3631
rect 20086 3171 20138 3177
rect 20086 3113 20138 3119
rect 19906 1836 20030 1864
rect 19906 800 19934 1836
rect 20098 800 20126 3113
rect 20194 3103 20222 5629
rect 20278 4355 20330 4361
rect 20278 4297 20330 4303
rect 20182 3097 20234 3103
rect 20182 3039 20234 3045
rect 20182 2505 20234 2511
rect 20182 2447 20234 2453
rect 20194 800 20222 2447
rect 20290 800 20318 4297
rect 20386 3251 20414 6887
rect 20482 6433 20510 14731
rect 20578 6581 20606 55579
rect 20758 55415 20810 55421
rect 20758 55357 20810 55363
rect 20662 35583 20714 35589
rect 20662 35525 20714 35531
rect 20674 12427 20702 35525
rect 20662 12421 20714 12427
rect 20662 12363 20714 12369
rect 20770 12224 20798 55357
rect 20866 20567 20894 56171
rect 21442 24119 21470 56171
rect 21430 24113 21482 24119
rect 21430 24055 21482 24061
rect 20950 22337 21002 22343
rect 20950 22279 21002 22285
rect 20854 20561 20906 20567
rect 20854 20503 20906 20509
rect 20854 19451 20906 19457
rect 20854 19393 20906 19399
rect 20866 12575 20894 19393
rect 20854 12569 20906 12575
rect 20854 12511 20906 12517
rect 20854 12421 20906 12427
rect 20854 12363 20906 12369
rect 20674 12196 20798 12224
rect 20674 7025 20702 12196
rect 20866 11539 20894 12363
rect 20854 11533 20906 11539
rect 20854 11475 20906 11481
rect 20962 7765 20990 22279
rect 21634 20937 21662 56837
rect 21730 56531 21758 59200
rect 22306 56975 22334 59200
rect 22294 56969 22346 56975
rect 22294 56911 22346 56917
rect 22786 56531 22814 59200
rect 23362 57614 23390 59200
rect 23362 57586 23486 57614
rect 23350 56895 23402 56901
rect 23350 56837 23402 56843
rect 21718 56525 21770 56531
rect 21718 56467 21770 56473
rect 22774 56525 22826 56531
rect 22774 56467 22826 56473
rect 22102 56229 22154 56235
rect 22102 56171 22154 56177
rect 22966 56229 23018 56235
rect 22966 56171 23018 56177
rect 21718 35583 21770 35589
rect 21718 35525 21770 35531
rect 21730 33887 21758 35525
rect 21718 33881 21770 33887
rect 21718 33823 21770 33829
rect 21622 20931 21674 20937
rect 21622 20873 21674 20879
rect 21526 20117 21578 20123
rect 21526 20059 21578 20065
rect 21538 17089 21566 20059
rect 21526 17083 21578 17089
rect 21526 17025 21578 17031
rect 21526 16935 21578 16941
rect 21526 16877 21578 16883
rect 21238 14789 21290 14795
rect 21238 14731 21290 14737
rect 20950 7759 21002 7765
rect 20950 7701 21002 7707
rect 20758 7463 20810 7469
rect 20758 7405 20810 7411
rect 20662 7019 20714 7025
rect 20662 6961 20714 6967
rect 20662 6871 20714 6877
rect 20662 6813 20714 6819
rect 20566 6575 20618 6581
rect 20566 6517 20618 6523
rect 20470 6427 20522 6433
rect 20470 6369 20522 6375
rect 20674 5860 20702 6813
rect 20482 5832 20702 5860
rect 20374 3245 20426 3251
rect 20374 3187 20426 3193
rect 20482 800 20510 5832
rect 20566 5687 20618 5693
rect 20566 5629 20618 5635
rect 20578 800 20606 5629
rect 20662 5021 20714 5027
rect 20662 4963 20714 4969
rect 20674 3843 20702 4963
rect 20662 3837 20714 3843
rect 20662 3779 20714 3785
rect 20662 3689 20714 3695
rect 20662 3631 20714 3637
rect 20674 800 20702 3631
rect 20770 800 20798 7405
rect 21250 7099 21278 14731
rect 21538 10947 21566 16877
rect 21526 10941 21578 10947
rect 21526 10883 21578 10889
rect 22114 10133 22142 56171
rect 22390 54749 22442 54755
rect 22390 54691 22442 54697
rect 22294 43427 22346 43433
rect 22294 43369 22346 43375
rect 22102 10127 22154 10133
rect 22102 10069 22154 10075
rect 21910 9831 21962 9837
rect 21910 9773 21962 9779
rect 21526 9239 21578 9245
rect 21526 9181 21578 9187
rect 21238 7093 21290 7099
rect 21238 7035 21290 7041
rect 21142 6945 21194 6951
rect 21142 6887 21194 6893
rect 20854 5021 20906 5027
rect 20854 4963 20906 4969
rect 20866 2511 20894 4963
rect 21046 4355 21098 4361
rect 21046 4297 21098 4303
rect 20950 2949 21002 2955
rect 20950 2891 21002 2897
rect 20854 2505 20906 2511
rect 20854 2447 20906 2453
rect 20962 800 20990 2891
rect 21058 800 21086 4297
rect 21154 800 21182 6887
rect 21538 6433 21566 9181
rect 21922 7099 21950 9773
rect 22102 8129 22154 8135
rect 22102 8071 22154 8077
rect 22114 7913 22142 8071
rect 22102 7907 22154 7913
rect 22102 7849 22154 7855
rect 22306 7173 22334 43369
rect 22402 10355 22430 54691
rect 22978 41805 23006 56171
rect 22966 41799 23018 41805
rect 22966 41741 23018 41747
rect 23254 24335 23306 24341
rect 23254 24277 23306 24283
rect 22390 10349 22442 10355
rect 22390 10291 22442 10297
rect 22966 9905 23018 9911
rect 22966 9847 23018 9853
rect 22294 7167 22346 7173
rect 22294 7109 22346 7115
rect 21910 7093 21962 7099
rect 21910 7035 21962 7041
rect 21910 6945 21962 6951
rect 21910 6887 21962 6893
rect 21526 6427 21578 6433
rect 21526 6369 21578 6375
rect 21430 6131 21482 6137
rect 21430 6073 21482 6079
rect 21526 6131 21578 6137
rect 21526 6073 21578 6079
rect 21238 3911 21290 3917
rect 21238 3853 21290 3859
rect 21250 800 21278 3853
rect 21442 3177 21470 6073
rect 21430 3171 21482 3177
rect 21430 3113 21482 3119
rect 21430 3023 21482 3029
rect 21430 2965 21482 2971
rect 21442 800 21470 2965
rect 21538 800 21566 6073
rect 21814 5687 21866 5693
rect 21634 5647 21814 5675
rect 21634 800 21662 5647
rect 21814 5629 21866 5635
rect 21718 5539 21770 5545
rect 21718 5481 21770 5487
rect 21730 2955 21758 5481
rect 21814 4355 21866 4361
rect 21814 4297 21866 4303
rect 21718 2949 21770 2955
rect 21718 2891 21770 2897
rect 21826 800 21854 4297
rect 21922 800 21950 6887
rect 22978 6433 23006 9847
rect 23158 7537 23210 7543
rect 23158 7479 23210 7485
rect 23170 7025 23198 7479
rect 23266 7173 23294 24277
rect 23362 11613 23390 56837
rect 23458 55717 23486 57586
rect 23842 56975 23870 59200
rect 23830 56969 23882 56975
rect 23830 56911 23882 56917
rect 24418 56531 24446 59200
rect 24406 56525 24458 56531
rect 24406 56467 24458 56473
rect 24406 56229 24458 56235
rect 24406 56171 24458 56177
rect 23446 55711 23498 55717
rect 23446 55653 23498 55659
rect 24310 55563 24362 55569
rect 24310 55505 24362 55511
rect 23734 39875 23786 39881
rect 23734 39817 23786 39823
rect 23638 25223 23690 25229
rect 23638 25165 23690 25171
rect 23350 11607 23402 11613
rect 23350 11549 23402 11555
rect 23254 7167 23306 7173
rect 23254 7109 23306 7115
rect 23158 7019 23210 7025
rect 23158 6961 23210 6967
rect 23350 6945 23402 6951
rect 23350 6887 23402 6893
rect 22966 6427 23018 6433
rect 22966 6369 23018 6375
rect 23062 5687 23114 5693
rect 23062 5629 23114 5635
rect 22774 5021 22826 5027
rect 22774 4963 22826 4969
rect 22006 4281 22058 4287
rect 22006 4223 22058 4229
rect 22018 800 22046 4223
rect 22786 3917 22814 4963
rect 22774 3911 22826 3917
rect 22774 3853 22826 3859
rect 22294 3837 22346 3843
rect 23074 3788 23102 5629
rect 23158 4947 23210 4953
rect 23158 4889 23210 4895
rect 22294 3779 22346 3785
rect 22102 3689 22154 3695
rect 22102 3631 22154 3637
rect 22114 800 22142 3631
rect 22306 800 22334 3779
rect 22786 3760 23102 3788
rect 22582 3541 22634 3547
rect 22582 3483 22634 3489
rect 22390 3097 22442 3103
rect 22390 3039 22442 3045
rect 22402 800 22430 3039
rect 22486 2949 22538 2955
rect 22486 2891 22538 2897
rect 22498 800 22526 2891
rect 22594 800 22622 3483
rect 22786 800 22814 3760
rect 22870 3689 22922 3695
rect 22870 3631 22922 3637
rect 22882 800 22910 3631
rect 22966 3171 23018 3177
rect 22966 3113 23018 3119
rect 22978 800 23006 3113
rect 23170 800 23198 4889
rect 23254 4355 23306 4361
rect 23254 4297 23306 4303
rect 23266 800 23294 4297
rect 23362 3547 23390 6887
rect 23650 6433 23678 25165
rect 23746 9763 23774 39817
rect 24022 30773 24074 30779
rect 24022 30715 24074 30721
rect 23830 26111 23882 26117
rect 23830 26053 23882 26059
rect 23734 9757 23786 9763
rect 23734 9699 23786 9705
rect 23734 7463 23786 7469
rect 23734 7405 23786 7411
rect 23638 6427 23690 6433
rect 23638 6369 23690 6375
rect 23638 6131 23690 6137
rect 23638 6073 23690 6079
rect 23446 5687 23498 5693
rect 23446 5629 23498 5635
rect 23350 3541 23402 3547
rect 23350 3483 23402 3489
rect 23350 3245 23402 3251
rect 23350 3187 23402 3193
rect 23362 800 23390 3187
rect 23458 800 23486 5629
rect 23542 5021 23594 5027
rect 23542 4963 23594 4969
rect 23554 3103 23582 4963
rect 23650 3843 23678 6073
rect 23638 3837 23690 3843
rect 23638 3779 23690 3785
rect 23638 3689 23690 3695
rect 23638 3631 23690 3637
rect 23542 3097 23594 3103
rect 23542 3039 23594 3045
rect 23650 800 23678 3631
rect 23746 800 23774 7405
rect 23842 7173 23870 26053
rect 24034 9911 24062 30715
rect 24322 27893 24350 55505
rect 24418 34331 24446 56171
rect 24898 55717 24926 59200
rect 25474 56975 25502 59200
rect 25462 56969 25514 56975
rect 25462 56911 25514 56917
rect 25954 56531 25982 59200
rect 26326 56895 26378 56901
rect 26326 56837 26378 56843
rect 25942 56525 25994 56531
rect 25942 56467 25994 56473
rect 26134 56229 26186 56235
rect 26134 56171 26186 56177
rect 24886 55711 24938 55717
rect 24886 55653 24938 55659
rect 26146 55643 26174 56171
rect 26134 55637 26186 55643
rect 26134 55579 26186 55585
rect 24982 55563 25034 55569
rect 24982 55505 25034 55511
rect 24406 34325 24458 34331
rect 24406 34267 24458 34273
rect 24502 32105 24554 32111
rect 24502 32047 24554 32053
rect 24514 31815 24542 32047
rect 24502 31809 24554 31815
rect 24502 31751 24554 31757
rect 24310 27887 24362 27893
rect 24310 27829 24362 27835
rect 24994 12205 25022 55505
rect 25654 43871 25706 43877
rect 25654 43813 25706 43819
rect 25174 41429 25226 41435
rect 25174 41371 25226 41377
rect 25078 40097 25130 40103
rect 25078 40039 25130 40045
rect 24982 12199 25034 12205
rect 24982 12141 25034 12147
rect 24502 11755 24554 11761
rect 24502 11697 24554 11703
rect 24118 11533 24170 11539
rect 24118 11475 24170 11481
rect 24022 9905 24074 9911
rect 24022 9847 24074 9853
rect 23926 9091 23978 9097
rect 23926 9033 23978 9039
rect 23938 7765 23966 9033
rect 23926 7759 23978 7765
rect 23926 7701 23978 7707
rect 23830 7167 23882 7173
rect 23830 7109 23882 7115
rect 24130 6581 24158 11475
rect 24514 9689 24542 11697
rect 24502 9683 24554 9689
rect 24502 9625 24554 9631
rect 24310 9609 24362 9615
rect 24310 9551 24362 9557
rect 24322 7839 24350 9551
rect 25090 7839 25118 40039
rect 25186 9837 25214 41371
rect 25462 24927 25514 24933
rect 25462 24869 25514 24875
rect 25174 9831 25226 9837
rect 25174 9773 25226 9779
rect 24310 7833 24362 7839
rect 24310 7775 24362 7781
rect 25078 7833 25130 7839
rect 25078 7775 25130 7781
rect 24790 7759 24842 7765
rect 24790 7701 24842 7707
rect 24694 7463 24746 7469
rect 24694 7405 24746 7411
rect 24214 6945 24266 6951
rect 24214 6887 24266 6893
rect 24502 6945 24554 6951
rect 24502 6887 24554 6893
rect 24118 6575 24170 6581
rect 24118 6517 24170 6523
rect 23926 6131 23978 6137
rect 23926 6073 23978 6079
rect 23938 3177 23966 6073
rect 24118 3763 24170 3769
rect 24118 3705 24170 3711
rect 23926 3171 23978 3177
rect 23926 3113 23978 3119
rect 23830 3097 23882 3103
rect 23830 3039 23882 3045
rect 23842 800 23870 3039
rect 24022 3023 24074 3029
rect 24022 2965 24074 2971
rect 24034 800 24062 2965
rect 24130 800 24158 3705
rect 24226 3251 24254 6887
rect 24406 3689 24458 3695
rect 24406 3631 24458 3637
rect 24214 3245 24266 3251
rect 24214 3187 24266 3193
rect 24214 2949 24266 2955
rect 24214 2891 24266 2897
rect 24226 800 24254 2891
rect 24418 1864 24446 3631
rect 24322 1836 24446 1864
rect 24322 800 24350 1836
rect 24514 800 24542 6887
rect 24598 5687 24650 5693
rect 24598 5629 24650 5635
rect 24610 800 24638 5629
rect 24706 3769 24734 7405
rect 24694 3763 24746 3769
rect 24694 3705 24746 3711
rect 24694 3615 24746 3621
rect 24694 3557 24746 3563
rect 24706 800 24734 3557
rect 24802 800 24830 7701
rect 25474 7617 25502 24869
rect 25462 7611 25514 7617
rect 25462 7553 25514 7559
rect 25666 7099 25694 43813
rect 25942 42761 25994 42767
rect 25942 42703 25994 42709
rect 25954 18865 25982 42703
rect 26134 42539 26186 42545
rect 26134 42481 26186 42487
rect 25942 18859 25994 18865
rect 25942 18801 25994 18807
rect 26038 13679 26090 13685
rect 26038 13621 26090 13627
rect 25942 7463 25994 7469
rect 25942 7405 25994 7411
rect 25654 7093 25706 7099
rect 25654 7035 25706 7041
rect 25174 6871 25226 6877
rect 25174 6813 25226 6819
rect 25078 5021 25130 5027
rect 25078 4963 25130 4969
rect 24886 4947 24938 4953
rect 24886 4889 24938 4895
rect 24898 2955 24926 4889
rect 24982 3171 25034 3177
rect 24982 3113 25034 3119
rect 24886 2949 24938 2955
rect 24886 2891 24938 2897
rect 24994 800 25022 3113
rect 25090 3103 25118 4963
rect 25078 3097 25130 3103
rect 25078 3039 25130 3045
rect 25078 2949 25130 2955
rect 25078 2891 25130 2897
rect 25090 800 25118 2891
rect 25186 800 25214 6813
rect 25654 6353 25706 6359
rect 25654 6295 25706 6301
rect 25462 4355 25514 4361
rect 25462 4297 25514 4303
rect 25366 3097 25418 3103
rect 25366 3039 25418 3045
rect 25378 800 25406 3039
rect 25474 800 25502 4297
rect 25558 3615 25610 3621
rect 25558 3557 25610 3563
rect 25570 800 25598 3557
rect 25666 800 25694 6295
rect 25954 3621 25982 7405
rect 26050 7173 26078 13621
rect 26146 7765 26174 42481
rect 26338 12871 26366 56837
rect 26530 56531 26558 59200
rect 27010 56975 27038 59200
rect 26998 56969 27050 56975
rect 26998 56911 27050 56917
rect 27586 56531 27614 59200
rect 28066 56531 28094 59200
rect 28642 56975 28670 59200
rect 29122 57049 29150 59200
rect 29110 57043 29162 57049
rect 29110 56985 29162 56991
rect 28630 56969 28682 56975
rect 28630 56911 28682 56917
rect 28822 56895 28874 56901
rect 28822 56837 28874 56843
rect 26518 56525 26570 56531
rect 26518 56467 26570 56473
rect 27574 56525 27626 56531
rect 27574 56467 27626 56473
rect 28054 56525 28106 56531
rect 28054 56467 28106 56473
rect 26902 56229 26954 56235
rect 26902 56171 26954 56177
rect 27766 56229 27818 56235
rect 27766 56171 27818 56177
rect 28150 56229 28202 56235
rect 28150 56171 28202 56177
rect 26914 52905 26942 56171
rect 26902 52899 26954 52905
rect 26902 52841 26954 52847
rect 26806 34769 26858 34775
rect 26806 34711 26858 34717
rect 26326 12865 26378 12871
rect 26326 12807 26378 12813
rect 26134 7759 26186 7765
rect 26134 7701 26186 7707
rect 26710 7463 26762 7469
rect 26710 7405 26762 7411
rect 26038 7167 26090 7173
rect 26038 7109 26090 7115
rect 26326 6131 26378 6137
rect 26326 6073 26378 6079
rect 26230 5687 26282 5693
rect 26230 5629 26282 5635
rect 26038 5539 26090 5545
rect 26038 5481 26090 5487
rect 25942 3615 25994 3621
rect 25942 3557 25994 3563
rect 25846 3541 25898 3547
rect 25846 3483 25898 3489
rect 25858 800 25886 3483
rect 25942 3245 25994 3251
rect 25942 3187 25994 3193
rect 25954 800 25982 3187
rect 26050 800 26078 5481
rect 26134 4355 26186 4361
rect 26134 4297 26186 4303
rect 26146 800 26174 4297
rect 26242 3103 26270 5629
rect 26230 3097 26282 3103
rect 26230 3039 26282 3045
rect 26338 800 26366 6073
rect 26614 5021 26666 5027
rect 26614 4963 26666 4969
rect 26518 4355 26570 4361
rect 26518 4297 26570 4303
rect 26422 3837 26474 3843
rect 26422 3779 26474 3785
rect 26434 800 26462 3779
rect 26530 800 26558 4297
rect 26626 3177 26654 4963
rect 26614 3171 26666 3177
rect 26614 3113 26666 3119
rect 26722 800 26750 7405
rect 26818 7173 26846 34711
rect 27382 32105 27434 32111
rect 27382 32047 27434 32053
rect 27394 31889 27422 32047
rect 27382 31883 27434 31889
rect 27382 31825 27434 31831
rect 26902 22781 26954 22787
rect 26902 22723 26954 22729
rect 26914 21899 26942 22723
rect 26902 21893 26954 21899
rect 26902 21835 26954 21841
rect 27778 15905 27806 56171
rect 27958 46165 28010 46171
rect 27958 46107 28010 46113
rect 27862 18859 27914 18865
rect 27862 18801 27914 18807
rect 27766 15899 27818 15905
rect 27766 15841 27818 15847
rect 27574 13901 27626 13907
rect 27574 13843 27626 13849
rect 27586 7173 27614 13843
rect 26806 7167 26858 7173
rect 26806 7109 26858 7115
rect 27574 7167 27626 7173
rect 27574 7109 27626 7115
rect 26902 6945 26954 6951
rect 26902 6887 26954 6893
rect 26806 6353 26858 6359
rect 26806 6295 26858 6301
rect 26818 800 26846 6295
rect 26914 3251 26942 6887
rect 26998 6871 27050 6877
rect 26998 6813 27050 6819
rect 27766 6871 27818 6877
rect 27766 6813 27818 6819
rect 26902 3245 26954 3251
rect 26902 3187 26954 3193
rect 26902 3023 26954 3029
rect 26902 2965 26954 2971
rect 26914 800 26942 2965
rect 27010 800 27038 6813
rect 27382 5687 27434 5693
rect 27382 5629 27434 5635
rect 27394 3788 27422 5629
rect 27202 3760 27422 3788
rect 27202 800 27230 3760
rect 27286 3689 27338 3695
rect 27286 3631 27338 3637
rect 27298 800 27326 3631
rect 27382 3245 27434 3251
rect 27382 3187 27434 3193
rect 27394 800 27422 3187
rect 27478 3097 27530 3103
rect 27478 3039 27530 3045
rect 27490 800 27518 3039
rect 27670 2949 27722 2955
rect 27670 2891 27722 2897
rect 27682 800 27710 2891
rect 27778 800 27806 6813
rect 27874 6581 27902 18801
rect 27970 11687 27998 46107
rect 28162 13167 28190 56171
rect 28834 13833 28862 56837
rect 29698 56531 29726 59200
rect 30178 56975 30206 59200
rect 30166 56969 30218 56975
rect 30166 56911 30218 56917
rect 30658 56531 30686 59200
rect 29686 56525 29738 56531
rect 29686 56467 29738 56473
rect 30646 56525 30698 56531
rect 30646 56467 30698 56473
rect 29590 56229 29642 56235
rect 29590 56171 29642 56177
rect 30934 56229 30986 56235
rect 30934 56171 30986 56177
rect 28918 40911 28970 40917
rect 28918 40853 28970 40859
rect 28822 13827 28874 13833
rect 28822 13769 28874 13775
rect 28150 13161 28202 13167
rect 28150 13103 28202 13109
rect 27958 11681 28010 11687
rect 27958 11623 28010 11629
rect 28054 8129 28106 8135
rect 28054 8071 28106 8077
rect 28066 7099 28094 8071
rect 28930 7913 28958 40853
rect 29494 30551 29546 30557
rect 29494 30493 29546 30499
rect 29014 13161 29066 13167
rect 29014 13103 29066 13109
rect 28918 7907 28970 7913
rect 28918 7849 28970 7855
rect 28930 7765 28958 7849
rect 28918 7759 28970 7765
rect 28918 7701 28970 7707
rect 28150 7463 28202 7469
rect 28150 7405 28202 7411
rect 28054 7093 28106 7099
rect 28054 7035 28106 7041
rect 27862 6575 27914 6581
rect 27862 6517 27914 6523
rect 27862 5687 27914 5693
rect 27862 5629 27914 5635
rect 27874 800 27902 5629
rect 28054 5021 28106 5027
rect 28054 4963 28106 4969
rect 28066 3843 28094 4963
rect 28054 3837 28106 3843
rect 28054 3779 28106 3785
rect 28054 3541 28106 3547
rect 28054 3483 28106 3489
rect 28066 800 28094 3483
rect 28162 800 28190 7405
rect 29026 6433 29054 13103
rect 29206 7463 29258 7469
rect 29206 7405 29258 7411
rect 29014 6427 29066 6433
rect 29014 6369 29066 6375
rect 28438 6131 28490 6137
rect 28438 6073 28490 6079
rect 28342 4355 28394 4361
rect 28342 4297 28394 4303
rect 28246 3171 28298 3177
rect 28246 3113 28298 3119
rect 28258 800 28286 3113
rect 28354 800 28382 4297
rect 28450 3251 28478 6073
rect 28822 5687 28874 5693
rect 28822 5629 28874 5635
rect 28834 3936 28862 5629
rect 28918 5021 28970 5027
rect 28918 4963 28970 4969
rect 28642 3908 28862 3936
rect 28438 3245 28490 3251
rect 28438 3187 28490 3193
rect 28534 3245 28586 3251
rect 28534 3187 28586 3193
rect 28546 800 28574 3187
rect 28642 800 28670 3908
rect 28822 3837 28874 3843
rect 28822 3779 28874 3785
rect 28726 3763 28778 3769
rect 28726 3705 28778 3711
rect 28738 800 28766 3705
rect 28834 2937 28862 3779
rect 28930 3103 28958 4963
rect 29110 4355 29162 4361
rect 29110 4297 29162 4303
rect 29014 3837 29066 3843
rect 29014 3779 29066 3785
rect 28918 3097 28970 3103
rect 28918 3039 28970 3045
rect 28834 2909 28958 2937
rect 28930 800 28958 2909
rect 29026 800 29054 3779
rect 29122 800 29150 4297
rect 29218 800 29246 7405
rect 29506 7099 29534 30493
rect 29602 13537 29630 56171
rect 29686 48903 29738 48909
rect 29686 48845 29738 48851
rect 29590 13531 29642 13537
rect 29590 13473 29642 13479
rect 29698 9097 29726 48845
rect 30550 38765 30602 38771
rect 30550 38707 30602 38713
rect 30166 13013 30218 13019
rect 30166 12955 30218 12961
rect 30178 11021 30206 12955
rect 30166 11015 30218 11021
rect 30166 10957 30218 10963
rect 30358 9609 30410 9615
rect 30358 9551 30410 9557
rect 30370 9097 30398 9551
rect 29686 9091 29738 9097
rect 29686 9033 29738 9039
rect 30358 9091 30410 9097
rect 30358 9033 30410 9039
rect 30166 7759 30218 7765
rect 30166 7701 30218 7707
rect 30178 7543 30206 7701
rect 30166 7537 30218 7543
rect 30166 7479 30218 7485
rect 29590 7463 29642 7469
rect 29590 7405 29642 7411
rect 29494 7093 29546 7099
rect 29494 7035 29546 7041
rect 29398 6945 29450 6951
rect 29398 6887 29450 6893
rect 29302 5021 29354 5027
rect 29302 4963 29354 4969
rect 29314 3177 29342 4963
rect 29410 3251 29438 6887
rect 29494 3615 29546 3621
rect 29494 3557 29546 3563
rect 29398 3245 29450 3251
rect 29398 3187 29450 3193
rect 29302 3171 29354 3177
rect 29302 3113 29354 3119
rect 29398 3097 29450 3103
rect 29398 3039 29450 3045
rect 29410 800 29438 3039
rect 29506 800 29534 3557
rect 29602 800 29630 7405
rect 30562 7173 30590 38707
rect 30946 37439 30974 56171
rect 31234 56161 31262 59200
rect 31714 56975 31742 59200
rect 31702 56969 31754 56975
rect 31702 56911 31754 56917
rect 31894 56895 31946 56901
rect 31894 56837 31946 56843
rect 31318 56229 31370 56235
rect 31318 56171 31370 56177
rect 31222 56155 31274 56161
rect 31222 56097 31274 56103
rect 30934 37433 30986 37439
rect 30934 37375 30986 37381
rect 30934 22781 30986 22787
rect 30934 22723 30986 22729
rect 30838 18267 30890 18273
rect 30838 18209 30890 18215
rect 30850 14203 30878 18209
rect 30838 14197 30890 14203
rect 30838 14139 30890 14145
rect 30946 9171 30974 22723
rect 31330 14499 31358 56171
rect 31606 45425 31658 45431
rect 31606 45367 31658 45373
rect 31510 38765 31562 38771
rect 31510 38707 31562 38713
rect 31414 34769 31466 34775
rect 31414 34711 31466 34717
rect 31426 24193 31454 34711
rect 31414 24187 31466 24193
rect 31414 24129 31466 24135
rect 31318 14493 31370 14499
rect 31318 14435 31370 14441
rect 31030 12125 31082 12131
rect 31030 12067 31082 12073
rect 31042 11761 31070 12067
rect 31030 11755 31082 11761
rect 31030 11697 31082 11703
rect 31522 11613 31550 38707
rect 31510 11607 31562 11613
rect 31510 11549 31562 11555
rect 30934 9165 30986 9171
rect 30934 9107 30986 9113
rect 30646 7611 30698 7617
rect 30646 7553 30698 7559
rect 30550 7167 30602 7173
rect 30550 7109 30602 7115
rect 29974 6945 30026 6951
rect 29974 6887 30026 6893
rect 29686 6353 29738 6359
rect 29686 6295 29738 6301
rect 29698 800 29726 6295
rect 29782 6131 29834 6137
rect 29782 6073 29834 6079
rect 29794 3917 29822 6073
rect 29782 3911 29834 3917
rect 29782 3853 29834 3859
rect 29782 3171 29834 3177
rect 29782 3113 29834 3119
rect 29794 2585 29822 3113
rect 29878 3023 29930 3029
rect 29878 2965 29930 2971
rect 29782 2579 29834 2585
rect 29782 2521 29834 2527
rect 29890 800 29918 2965
rect 29986 800 30014 6887
rect 30658 6452 30686 7553
rect 31030 7463 31082 7469
rect 31030 7405 31082 7411
rect 30562 6424 30686 6452
rect 30262 5687 30314 5693
rect 30262 5629 30314 5635
rect 30274 2900 30302 5629
rect 30358 5021 30410 5027
rect 30358 4963 30410 4969
rect 30370 3843 30398 4963
rect 30358 3837 30410 3843
rect 30358 3779 30410 3785
rect 30454 3689 30506 3695
rect 30082 2872 30302 2900
rect 30370 3649 30454 3677
rect 30082 800 30110 2872
rect 30370 1864 30398 3649
rect 30454 3631 30506 3637
rect 30454 3245 30506 3251
rect 30454 3187 30506 3193
rect 30274 1836 30398 1864
rect 30274 800 30302 1836
rect 30358 1765 30410 1771
rect 30358 1707 30410 1713
rect 30370 800 30398 1707
rect 30466 800 30494 3187
rect 30562 3177 30590 6424
rect 30646 6279 30698 6285
rect 30646 6221 30698 6227
rect 30658 5471 30686 6221
rect 30742 6131 30794 6137
rect 30742 6073 30794 6079
rect 30646 5465 30698 5471
rect 30646 5407 30698 5413
rect 30754 3677 30782 6073
rect 30838 5687 30890 5693
rect 30838 5629 30890 5635
rect 30658 3649 30782 3677
rect 30550 3171 30602 3177
rect 30550 3113 30602 3119
rect 30550 2949 30602 2955
rect 30550 2891 30602 2897
rect 30562 800 30590 2891
rect 30658 1771 30686 3649
rect 30742 3615 30794 3621
rect 30742 3557 30794 3563
rect 30646 1765 30698 1771
rect 30646 1707 30698 1713
rect 30754 800 30782 3557
rect 30850 800 30878 5629
rect 30934 4355 30986 4361
rect 30934 4297 30986 4303
rect 30946 800 30974 4297
rect 31042 800 31070 7405
rect 31618 7099 31646 45367
rect 31906 15165 31934 56837
rect 32290 56531 32318 59200
rect 32770 57614 32798 59200
rect 32770 57586 32894 57614
rect 32758 56895 32810 56901
rect 32758 56837 32810 56843
rect 32278 56525 32330 56531
rect 32278 56467 32330 56473
rect 32470 56229 32522 56235
rect 32470 56171 32522 56177
rect 32482 49575 32510 56171
rect 32470 49569 32522 49575
rect 32470 49511 32522 49517
rect 32770 39215 32798 56837
rect 32866 56531 32894 57586
rect 33346 56975 33374 59200
rect 33334 56969 33386 56975
rect 33334 56911 33386 56917
rect 33826 56531 33854 59200
rect 34102 56895 34154 56901
rect 34102 56837 34154 56843
rect 32854 56525 32906 56531
rect 32854 56467 32906 56473
rect 33814 56525 33866 56531
rect 33814 56467 33866 56473
rect 34006 56229 34058 56235
rect 34006 56171 34058 56177
rect 33910 40763 33962 40769
rect 33910 40705 33962 40711
rect 32758 39209 32810 39215
rect 32758 39151 32810 39157
rect 32662 38099 32714 38105
rect 32662 38041 32714 38047
rect 32374 36545 32426 36551
rect 32374 36487 32426 36493
rect 31894 15159 31946 15165
rect 31894 15101 31946 15107
rect 32386 9911 32414 36487
rect 32566 35583 32618 35589
rect 32566 35525 32618 35531
rect 32470 24853 32522 24859
rect 32470 24795 32522 24801
rect 32374 9905 32426 9911
rect 32374 9847 32426 9853
rect 32374 7611 32426 7617
rect 32374 7553 32426 7559
rect 32386 7247 32414 7553
rect 32374 7241 32426 7247
rect 32374 7183 32426 7189
rect 32482 7099 32510 24795
rect 32578 9541 32606 35525
rect 32674 13167 32702 38041
rect 32758 22559 32810 22565
rect 32758 22501 32810 22507
rect 32662 13161 32714 13167
rect 32662 13103 32714 13109
rect 32770 9837 32798 22501
rect 33814 13753 33866 13759
rect 33814 13695 33866 13701
rect 33142 9905 33194 9911
rect 33142 9847 33194 9853
rect 32758 9831 32810 9837
rect 32758 9773 32810 9779
rect 32566 9535 32618 9541
rect 32566 9477 32618 9483
rect 31606 7093 31658 7099
rect 31606 7035 31658 7041
rect 32470 7093 32522 7099
rect 32470 7035 32522 7041
rect 31798 6945 31850 6951
rect 31798 6887 31850 6893
rect 32374 6945 32426 6951
rect 32374 6887 32426 6893
rect 31222 6353 31274 6359
rect 31222 6295 31274 6301
rect 31126 5021 31178 5027
rect 31126 4963 31178 4969
rect 31138 3103 31166 4963
rect 31126 3097 31178 3103
rect 31126 3039 31178 3045
rect 31234 800 31262 6295
rect 31702 5687 31754 5693
rect 31702 5629 31754 5635
rect 31714 4528 31742 5629
rect 31618 4500 31742 4528
rect 31318 3689 31370 3695
rect 31318 3631 31370 3637
rect 31330 800 31358 3631
rect 31414 3541 31466 3547
rect 31414 3483 31466 3489
rect 31426 800 31454 3483
rect 31618 800 31646 4500
rect 31702 4355 31754 4361
rect 31702 4297 31754 4303
rect 31714 800 31742 4297
rect 31810 3621 31838 6887
rect 32182 6871 32234 6877
rect 32182 6813 32234 6819
rect 31894 5021 31946 5027
rect 31894 4963 31946 4969
rect 31798 3615 31850 3621
rect 31798 3557 31850 3563
rect 31906 3251 31934 4963
rect 31990 3911 32042 3917
rect 31990 3853 32042 3859
rect 31894 3245 31946 3251
rect 31894 3187 31946 3193
rect 32002 3177 32030 3853
rect 31798 3171 31850 3177
rect 31798 3113 31850 3119
rect 31990 3171 32042 3177
rect 31990 3113 32042 3119
rect 31810 800 31838 3113
rect 31894 3097 31946 3103
rect 31894 3039 31946 3045
rect 31906 800 31934 3039
rect 32086 3023 32138 3029
rect 32086 2965 32138 2971
rect 32098 800 32126 2965
rect 32194 800 32222 6813
rect 32386 3547 32414 6887
rect 32950 6797 33002 6803
rect 32950 6739 33002 6745
rect 32758 4355 32810 4361
rect 32758 4297 32810 4303
rect 32470 3689 32522 3695
rect 32470 3631 32522 3637
rect 32374 3541 32426 3547
rect 32374 3483 32426 3489
rect 32278 2949 32330 2955
rect 32278 2891 32330 2897
rect 32290 800 32318 2891
rect 32482 800 32510 3631
rect 32662 3245 32714 3251
rect 32662 3187 32714 3193
rect 32566 3171 32618 3177
rect 32566 3113 32618 3119
rect 32578 800 32606 3113
rect 32674 800 32702 3187
rect 32770 800 32798 4297
rect 32962 800 32990 6739
rect 33154 6581 33182 9847
rect 33826 7765 33854 13695
rect 33922 8431 33950 40705
rect 34018 30927 34046 56171
rect 34006 30921 34058 30927
rect 34006 30863 34058 30869
rect 34114 15535 34142 56837
rect 34402 56531 34430 59200
rect 34882 56975 34910 59200
rect 34988 57304 35284 57324
rect 35044 57302 35068 57304
rect 35124 57302 35148 57304
rect 35204 57302 35228 57304
rect 35066 57250 35068 57302
rect 35130 57250 35142 57302
rect 35204 57250 35206 57302
rect 35044 57248 35068 57250
rect 35124 57248 35148 57250
rect 35204 57248 35228 57250
rect 34988 57228 35284 57248
rect 34870 56969 34922 56975
rect 34870 56911 34922 56917
rect 34870 56821 34922 56827
rect 34870 56763 34922 56769
rect 34390 56525 34442 56531
rect 34390 56467 34442 56473
rect 34774 56229 34826 56235
rect 34774 56171 34826 56177
rect 34786 25007 34814 56171
rect 34774 25001 34826 25007
rect 34774 24943 34826 24949
rect 34678 18785 34730 18791
rect 34678 18727 34730 18733
rect 34102 15529 34154 15535
rect 34102 15471 34154 15477
rect 34390 14123 34442 14129
rect 34390 14065 34442 14071
rect 34006 9831 34058 9837
rect 34006 9773 34058 9779
rect 33910 8425 33962 8431
rect 33910 8367 33962 8373
rect 33814 7759 33866 7765
rect 33814 7701 33866 7707
rect 33622 7463 33674 7469
rect 33622 7405 33674 7411
rect 33142 6575 33194 6581
rect 33142 6517 33194 6523
rect 33526 6131 33578 6137
rect 33526 6073 33578 6079
rect 33142 5687 33194 5693
rect 33142 5629 33194 5635
rect 33238 5687 33290 5693
rect 33238 5629 33290 5635
rect 33154 2955 33182 5629
rect 33142 2949 33194 2955
rect 33142 2891 33194 2897
rect 33250 2752 33278 5629
rect 33334 5021 33386 5027
rect 33334 4963 33386 4969
rect 33346 3103 33374 4963
rect 33538 3917 33566 6073
rect 33526 3911 33578 3917
rect 33526 3853 33578 3859
rect 33430 3837 33482 3843
rect 33430 3779 33482 3785
rect 33334 3097 33386 3103
rect 33334 3039 33386 3045
rect 33334 2949 33386 2955
rect 33334 2891 33386 2897
rect 33058 2724 33278 2752
rect 33058 800 33086 2724
rect 33346 1420 33374 2891
rect 33154 1392 33374 1420
rect 33154 800 33182 1392
rect 33238 1321 33290 1327
rect 33238 1263 33290 1269
rect 33250 800 33278 1263
rect 33442 800 33470 3779
rect 33526 3689 33578 3695
rect 33526 3631 33578 3637
rect 33538 800 33566 3631
rect 33634 800 33662 7405
rect 34018 7099 34046 9773
rect 34294 9757 34346 9763
rect 34294 9699 34346 9705
rect 34006 7093 34058 7099
rect 34006 7035 34058 7041
rect 34306 6433 34334 9699
rect 34402 8431 34430 14065
rect 34582 10941 34634 10947
rect 34582 10883 34634 10889
rect 34390 8425 34442 8431
rect 34390 8367 34442 8373
rect 34594 7765 34622 10883
rect 34582 7759 34634 7765
rect 34582 7701 34634 7707
rect 34390 7463 34442 7469
rect 34390 7405 34442 7411
rect 34294 6427 34346 6433
rect 34294 6369 34346 6375
rect 33814 6353 33866 6359
rect 33814 6295 33866 6301
rect 33718 6131 33770 6137
rect 33718 6073 33770 6079
rect 33730 3177 33758 6073
rect 33718 3171 33770 3177
rect 33718 3113 33770 3119
rect 33826 3085 33854 6295
rect 34102 5021 34154 5027
rect 34102 4963 34154 4969
rect 33910 4355 33962 4361
rect 33910 4297 33962 4303
rect 33730 3057 33854 3085
rect 33730 1327 33758 3057
rect 33814 2801 33866 2807
rect 33814 2743 33866 2749
rect 33826 2511 33854 2743
rect 33814 2505 33866 2511
rect 33814 2447 33866 2453
rect 33814 2357 33866 2363
rect 33814 2299 33866 2305
rect 33718 1321 33770 1327
rect 33718 1263 33770 1269
rect 33826 800 33854 2299
rect 33922 800 33950 4297
rect 34114 3251 34142 4963
rect 34198 4281 34250 4287
rect 34198 4223 34250 4229
rect 34102 3245 34154 3251
rect 34102 3187 34154 3193
rect 34006 3097 34058 3103
rect 34006 3039 34058 3045
rect 34018 800 34046 3039
rect 34210 1420 34238 4223
rect 34294 3689 34346 3695
rect 34294 3631 34346 3637
rect 34114 1392 34238 1420
rect 34114 800 34142 1392
rect 34306 800 34334 3631
rect 34402 800 34430 7405
rect 34582 6945 34634 6951
rect 34582 6887 34634 6893
rect 34594 4528 34622 6887
rect 34690 6581 34718 18727
rect 34882 15461 34910 56763
rect 35458 56531 35486 59200
rect 35938 57614 35966 59200
rect 35938 57586 36062 57614
rect 35446 56525 35498 56531
rect 35446 56467 35498 56473
rect 36034 56457 36062 57586
rect 36514 56975 36542 59200
rect 36502 56969 36554 56975
rect 36502 56911 36554 56917
rect 36022 56451 36074 56457
rect 36022 56393 36074 56399
rect 35350 56229 35402 56235
rect 35350 56171 35402 56177
rect 36886 56229 36938 56235
rect 36886 56171 36938 56177
rect 34988 55972 35284 55992
rect 35044 55970 35068 55972
rect 35124 55970 35148 55972
rect 35204 55970 35228 55972
rect 35066 55918 35068 55970
rect 35130 55918 35142 55970
rect 35204 55918 35206 55970
rect 35044 55916 35068 55918
rect 35124 55916 35148 55918
rect 35204 55916 35228 55918
rect 34988 55896 35284 55916
rect 34988 54640 35284 54660
rect 35044 54638 35068 54640
rect 35124 54638 35148 54640
rect 35204 54638 35228 54640
rect 35066 54586 35068 54638
rect 35130 54586 35142 54638
rect 35204 54586 35206 54638
rect 35044 54584 35068 54586
rect 35124 54584 35148 54586
rect 35204 54584 35228 54586
rect 34988 54564 35284 54584
rect 34988 53308 35284 53328
rect 35044 53306 35068 53308
rect 35124 53306 35148 53308
rect 35204 53306 35228 53308
rect 35066 53254 35068 53306
rect 35130 53254 35142 53306
rect 35204 53254 35206 53306
rect 35044 53252 35068 53254
rect 35124 53252 35148 53254
rect 35204 53252 35228 53254
rect 34988 53232 35284 53252
rect 35362 53053 35390 56171
rect 35350 53047 35402 53053
rect 35350 52989 35402 52995
rect 34988 51976 35284 51996
rect 35044 51974 35068 51976
rect 35124 51974 35148 51976
rect 35204 51974 35228 51976
rect 35066 51922 35068 51974
rect 35130 51922 35142 51974
rect 35204 51922 35206 51974
rect 35044 51920 35068 51922
rect 35124 51920 35148 51922
rect 35204 51920 35228 51922
rect 34988 51900 35284 51920
rect 34988 50644 35284 50664
rect 35044 50642 35068 50644
rect 35124 50642 35148 50644
rect 35204 50642 35228 50644
rect 35066 50590 35068 50642
rect 35130 50590 35142 50642
rect 35204 50590 35206 50642
rect 35044 50588 35068 50590
rect 35124 50588 35148 50590
rect 35204 50588 35228 50590
rect 34988 50568 35284 50588
rect 34988 49312 35284 49332
rect 35044 49310 35068 49312
rect 35124 49310 35148 49312
rect 35204 49310 35228 49312
rect 35066 49258 35068 49310
rect 35130 49258 35142 49310
rect 35204 49258 35206 49310
rect 35044 49256 35068 49258
rect 35124 49256 35148 49258
rect 35204 49256 35228 49258
rect 34988 49236 35284 49256
rect 34988 47980 35284 48000
rect 35044 47978 35068 47980
rect 35124 47978 35148 47980
rect 35204 47978 35228 47980
rect 35066 47926 35068 47978
rect 35130 47926 35142 47978
rect 35204 47926 35206 47978
rect 35044 47924 35068 47926
rect 35124 47924 35148 47926
rect 35204 47924 35228 47926
rect 34988 47904 35284 47924
rect 34988 46648 35284 46668
rect 35044 46646 35068 46648
rect 35124 46646 35148 46648
rect 35204 46646 35228 46648
rect 35066 46594 35068 46646
rect 35130 46594 35142 46646
rect 35204 46594 35206 46646
rect 35044 46592 35068 46594
rect 35124 46592 35148 46594
rect 35204 46592 35228 46594
rect 34988 46572 35284 46592
rect 34988 45316 35284 45336
rect 35044 45314 35068 45316
rect 35124 45314 35148 45316
rect 35204 45314 35228 45316
rect 35066 45262 35068 45314
rect 35130 45262 35142 45314
rect 35204 45262 35206 45314
rect 35044 45260 35068 45262
rect 35124 45260 35148 45262
rect 35204 45260 35228 45262
rect 34988 45240 35284 45260
rect 34988 43984 35284 44004
rect 35044 43982 35068 43984
rect 35124 43982 35148 43984
rect 35204 43982 35228 43984
rect 35066 43930 35068 43982
rect 35130 43930 35142 43982
rect 35204 43930 35206 43982
rect 35044 43928 35068 43930
rect 35124 43928 35148 43930
rect 35204 43928 35228 43930
rect 34988 43908 35284 43928
rect 34988 42652 35284 42672
rect 35044 42650 35068 42652
rect 35124 42650 35148 42652
rect 35204 42650 35228 42652
rect 35066 42598 35068 42650
rect 35130 42598 35142 42650
rect 35204 42598 35206 42650
rect 35044 42596 35068 42598
rect 35124 42596 35148 42598
rect 35204 42596 35228 42598
rect 34988 42576 35284 42596
rect 34988 41320 35284 41340
rect 35044 41318 35068 41320
rect 35124 41318 35148 41320
rect 35204 41318 35228 41320
rect 35066 41266 35068 41318
rect 35130 41266 35142 41318
rect 35204 41266 35206 41318
rect 35044 41264 35068 41266
rect 35124 41264 35148 41266
rect 35204 41264 35228 41266
rect 34988 41244 35284 41264
rect 34988 39988 35284 40008
rect 35044 39986 35068 39988
rect 35124 39986 35148 39988
rect 35204 39986 35228 39988
rect 35066 39934 35068 39986
rect 35130 39934 35142 39986
rect 35204 39934 35206 39986
rect 35044 39932 35068 39934
rect 35124 39932 35148 39934
rect 35204 39932 35228 39934
rect 34988 39912 35284 39932
rect 34988 38656 35284 38676
rect 35044 38654 35068 38656
rect 35124 38654 35148 38656
rect 35204 38654 35228 38656
rect 35066 38602 35068 38654
rect 35130 38602 35142 38654
rect 35204 38602 35206 38654
rect 35044 38600 35068 38602
rect 35124 38600 35148 38602
rect 35204 38600 35228 38602
rect 34988 38580 35284 38600
rect 34988 37324 35284 37344
rect 35044 37322 35068 37324
rect 35124 37322 35148 37324
rect 35204 37322 35228 37324
rect 35066 37270 35068 37322
rect 35130 37270 35142 37322
rect 35204 37270 35206 37322
rect 35044 37268 35068 37270
rect 35124 37268 35148 37270
rect 35204 37268 35228 37270
rect 34988 37248 35284 37268
rect 34988 35992 35284 36012
rect 35044 35990 35068 35992
rect 35124 35990 35148 35992
rect 35204 35990 35228 35992
rect 35066 35938 35068 35990
rect 35130 35938 35142 35990
rect 35204 35938 35206 35990
rect 35044 35936 35068 35938
rect 35124 35936 35148 35938
rect 35204 35936 35228 35938
rect 34988 35916 35284 35936
rect 34988 34660 35284 34680
rect 35044 34658 35068 34660
rect 35124 34658 35148 34660
rect 35204 34658 35228 34660
rect 35066 34606 35068 34658
rect 35130 34606 35142 34658
rect 35204 34606 35206 34658
rect 35044 34604 35068 34606
rect 35124 34604 35148 34606
rect 35204 34604 35228 34606
rect 34988 34584 35284 34604
rect 34988 33328 35284 33348
rect 35044 33326 35068 33328
rect 35124 33326 35148 33328
rect 35204 33326 35228 33328
rect 35066 33274 35068 33326
rect 35130 33274 35142 33326
rect 35204 33274 35206 33326
rect 35044 33272 35068 33274
rect 35124 33272 35148 33274
rect 35204 33272 35228 33274
rect 34988 33252 35284 33272
rect 34988 31996 35284 32016
rect 35044 31994 35068 31996
rect 35124 31994 35148 31996
rect 35204 31994 35228 31996
rect 35066 31942 35068 31994
rect 35130 31942 35142 31994
rect 35204 31942 35206 31994
rect 35044 31940 35068 31942
rect 35124 31940 35148 31942
rect 35204 31940 35228 31942
rect 34988 31920 35284 31940
rect 35446 31809 35498 31815
rect 35446 31751 35498 31757
rect 35350 31735 35402 31741
rect 35350 31677 35402 31683
rect 34988 30664 35284 30684
rect 35044 30662 35068 30664
rect 35124 30662 35148 30664
rect 35204 30662 35228 30664
rect 35066 30610 35068 30662
rect 35130 30610 35142 30662
rect 35204 30610 35206 30662
rect 35044 30608 35068 30610
rect 35124 30608 35148 30610
rect 35204 30608 35228 30610
rect 34988 30588 35284 30608
rect 34988 29332 35284 29352
rect 35044 29330 35068 29332
rect 35124 29330 35148 29332
rect 35204 29330 35228 29332
rect 35066 29278 35068 29330
rect 35130 29278 35142 29330
rect 35204 29278 35206 29330
rect 35044 29276 35068 29278
rect 35124 29276 35148 29278
rect 35204 29276 35228 29278
rect 34988 29256 35284 29276
rect 34988 28000 35284 28020
rect 35044 27998 35068 28000
rect 35124 27998 35148 28000
rect 35204 27998 35228 28000
rect 35066 27946 35068 27998
rect 35130 27946 35142 27998
rect 35204 27946 35206 27998
rect 35044 27944 35068 27946
rect 35124 27944 35148 27946
rect 35204 27944 35228 27946
rect 34988 27924 35284 27944
rect 34988 26668 35284 26688
rect 35044 26666 35068 26668
rect 35124 26666 35148 26668
rect 35204 26666 35228 26668
rect 35066 26614 35068 26666
rect 35130 26614 35142 26666
rect 35204 26614 35206 26666
rect 35044 26612 35068 26614
rect 35124 26612 35148 26614
rect 35204 26612 35228 26614
rect 34988 26592 35284 26612
rect 34988 25336 35284 25356
rect 35044 25334 35068 25336
rect 35124 25334 35148 25336
rect 35204 25334 35228 25336
rect 35066 25282 35068 25334
rect 35130 25282 35142 25334
rect 35204 25282 35206 25334
rect 35044 25280 35068 25282
rect 35124 25280 35148 25282
rect 35204 25280 35228 25282
rect 34988 25260 35284 25280
rect 34988 24004 35284 24024
rect 35044 24002 35068 24004
rect 35124 24002 35148 24004
rect 35204 24002 35228 24004
rect 35066 23950 35068 24002
rect 35130 23950 35142 24002
rect 35204 23950 35206 24002
rect 35044 23948 35068 23950
rect 35124 23948 35148 23950
rect 35204 23948 35228 23950
rect 34988 23928 35284 23948
rect 34988 22672 35284 22692
rect 35044 22670 35068 22672
rect 35124 22670 35148 22672
rect 35204 22670 35228 22672
rect 35066 22618 35068 22670
rect 35130 22618 35142 22670
rect 35204 22618 35206 22670
rect 35044 22616 35068 22618
rect 35124 22616 35148 22618
rect 35204 22616 35228 22618
rect 34988 22596 35284 22616
rect 34988 21340 35284 21360
rect 35044 21338 35068 21340
rect 35124 21338 35148 21340
rect 35204 21338 35228 21340
rect 35066 21286 35068 21338
rect 35130 21286 35142 21338
rect 35204 21286 35206 21338
rect 35044 21284 35068 21286
rect 35124 21284 35148 21286
rect 35204 21284 35228 21286
rect 34988 21264 35284 21284
rect 34988 20008 35284 20028
rect 35044 20006 35068 20008
rect 35124 20006 35148 20008
rect 35204 20006 35228 20008
rect 35066 19954 35068 20006
rect 35130 19954 35142 20006
rect 35204 19954 35206 20006
rect 35044 19952 35068 19954
rect 35124 19952 35148 19954
rect 35204 19952 35228 19954
rect 34988 19932 35284 19952
rect 34988 18676 35284 18696
rect 35044 18674 35068 18676
rect 35124 18674 35148 18676
rect 35204 18674 35228 18676
rect 35066 18622 35068 18674
rect 35130 18622 35142 18674
rect 35204 18622 35206 18674
rect 35044 18620 35068 18622
rect 35124 18620 35148 18622
rect 35204 18620 35228 18622
rect 34988 18600 35284 18620
rect 34988 17344 35284 17364
rect 35044 17342 35068 17344
rect 35124 17342 35148 17344
rect 35204 17342 35228 17344
rect 35066 17290 35068 17342
rect 35130 17290 35142 17342
rect 35204 17290 35206 17342
rect 35044 17288 35068 17290
rect 35124 17288 35148 17290
rect 35204 17288 35228 17290
rect 34988 17268 35284 17288
rect 34988 16012 35284 16032
rect 35044 16010 35068 16012
rect 35124 16010 35148 16012
rect 35204 16010 35228 16012
rect 35066 15958 35068 16010
rect 35130 15958 35142 16010
rect 35204 15958 35206 16010
rect 35044 15956 35068 15958
rect 35124 15956 35148 15958
rect 35204 15956 35228 15958
rect 34988 15936 35284 15956
rect 34870 15455 34922 15461
rect 34870 15397 34922 15403
rect 34988 14680 35284 14700
rect 35044 14678 35068 14680
rect 35124 14678 35148 14680
rect 35204 14678 35228 14680
rect 35066 14626 35068 14678
rect 35130 14626 35142 14678
rect 35204 14626 35206 14678
rect 35044 14624 35068 14626
rect 35124 14624 35148 14626
rect 35204 14624 35228 14626
rect 34988 14604 35284 14624
rect 34988 13348 35284 13368
rect 35044 13346 35068 13348
rect 35124 13346 35148 13348
rect 35204 13346 35228 13348
rect 35066 13294 35068 13346
rect 35130 13294 35142 13346
rect 35204 13294 35206 13346
rect 35044 13292 35068 13294
rect 35124 13292 35148 13294
rect 35204 13292 35228 13294
rect 34988 13272 35284 13292
rect 34988 12016 35284 12036
rect 35044 12014 35068 12016
rect 35124 12014 35148 12016
rect 35204 12014 35228 12016
rect 35066 11962 35068 12014
rect 35130 11962 35142 12014
rect 35204 11962 35206 12014
rect 35044 11960 35068 11962
rect 35124 11960 35148 11962
rect 35204 11960 35228 11962
rect 34988 11940 35284 11960
rect 34988 10684 35284 10704
rect 35044 10682 35068 10684
rect 35124 10682 35148 10684
rect 35204 10682 35228 10684
rect 35066 10630 35068 10682
rect 35130 10630 35142 10682
rect 35204 10630 35206 10682
rect 35044 10628 35068 10630
rect 35124 10628 35148 10630
rect 35204 10628 35228 10630
rect 34988 10608 35284 10628
rect 34988 9352 35284 9372
rect 35044 9350 35068 9352
rect 35124 9350 35148 9352
rect 35204 9350 35228 9352
rect 35066 9298 35068 9350
rect 35130 9298 35142 9350
rect 35204 9298 35206 9350
rect 35044 9296 35068 9298
rect 35124 9296 35148 9298
rect 35204 9296 35228 9298
rect 34988 9276 35284 9296
rect 35062 8869 35114 8875
rect 35062 8811 35114 8817
rect 35074 8431 35102 8811
rect 35062 8425 35114 8431
rect 35062 8367 35114 8373
rect 34988 8020 35284 8040
rect 35044 8018 35068 8020
rect 35124 8018 35148 8020
rect 35204 8018 35228 8020
rect 35066 7966 35068 8018
rect 35130 7966 35142 8018
rect 35204 7966 35206 8018
rect 35044 7964 35068 7966
rect 35124 7964 35148 7966
rect 35204 7964 35228 7966
rect 34988 7944 35284 7964
rect 35362 7765 35390 31677
rect 35458 9837 35486 31751
rect 35542 27665 35594 27671
rect 35542 27607 35594 27613
rect 35554 10133 35582 27607
rect 36898 22491 36926 56171
rect 36994 56087 37022 59200
rect 37570 56531 37598 59200
rect 38050 56901 38078 59200
rect 38038 56895 38090 56901
rect 38038 56837 38090 56843
rect 37942 56747 37994 56753
rect 37942 56689 37994 56695
rect 37558 56525 37610 56531
rect 37558 56467 37610 56473
rect 37462 56229 37514 56235
rect 37462 56171 37514 56177
rect 36982 56081 37034 56087
rect 36982 56023 37034 56029
rect 37078 29441 37130 29447
rect 37078 29383 37130 29389
rect 37090 29225 37118 29383
rect 37078 29219 37130 29225
rect 37078 29161 37130 29167
rect 36886 22485 36938 22491
rect 36886 22427 36938 22433
rect 35638 22189 35690 22195
rect 35638 22131 35690 22137
rect 35542 10127 35594 10133
rect 35542 10069 35594 10075
rect 35650 9911 35678 22131
rect 35734 15899 35786 15905
rect 35734 15841 35786 15847
rect 35638 9905 35690 9911
rect 35638 9847 35690 9853
rect 35446 9831 35498 9837
rect 35446 9773 35498 9779
rect 35746 9763 35774 15841
rect 37474 15831 37502 56171
rect 37954 16497 37982 56689
rect 38626 56531 38654 59200
rect 38614 56525 38666 56531
rect 38614 56467 38666 56473
rect 38422 56229 38474 56235
rect 38422 56171 38474 56177
rect 38134 33437 38186 33443
rect 38134 33379 38186 33385
rect 37942 16491 37994 16497
rect 37942 16433 37994 16439
rect 37462 15825 37514 15831
rect 37462 15767 37514 15773
rect 36598 14863 36650 14869
rect 36598 14805 36650 14811
rect 36610 14573 36638 14805
rect 36598 14567 36650 14573
rect 36598 14509 36650 14515
rect 37750 13827 37802 13833
rect 37750 13769 37802 13775
rect 36502 11607 36554 11613
rect 36502 11549 36554 11555
rect 36118 10127 36170 10133
rect 36118 10069 36170 10075
rect 35734 9757 35786 9763
rect 35734 9699 35786 9705
rect 36130 7765 36158 10069
rect 36214 9905 36266 9911
rect 36214 9847 36266 9853
rect 35350 7759 35402 7765
rect 35350 7701 35402 7707
rect 36118 7759 36170 7765
rect 36118 7701 36170 7707
rect 34774 7463 34826 7469
rect 34774 7405 34826 7411
rect 35830 7463 35882 7469
rect 35830 7405 35882 7411
rect 34678 6575 34730 6581
rect 34678 6517 34730 6523
rect 34678 5687 34730 5693
rect 34678 5629 34730 5635
rect 34498 4500 34622 4528
rect 34498 3103 34526 4500
rect 34582 4355 34634 4361
rect 34582 4297 34634 4303
rect 34486 3097 34538 3103
rect 34486 3039 34538 3045
rect 34484 2914 34540 2923
rect 34484 2849 34540 2858
rect 34498 800 34526 2849
rect 34594 800 34622 4297
rect 34690 2363 34718 5629
rect 34678 2357 34730 2363
rect 34678 2299 34730 2305
rect 34786 800 34814 7405
rect 35734 6945 35786 6951
rect 35734 6887 35786 6893
rect 34988 6688 35284 6708
rect 35044 6686 35068 6688
rect 35124 6686 35148 6688
rect 35204 6686 35228 6688
rect 35066 6634 35068 6686
rect 35130 6634 35142 6686
rect 35204 6634 35206 6686
rect 35044 6632 35068 6634
rect 35124 6632 35148 6634
rect 35204 6632 35228 6634
rect 34988 6612 35284 6632
rect 35746 6581 35774 6887
rect 35734 6575 35786 6581
rect 35734 6517 35786 6523
rect 35446 6427 35498 6433
rect 35446 6369 35498 6375
rect 34988 5356 35284 5376
rect 35044 5354 35068 5356
rect 35124 5354 35148 5356
rect 35204 5354 35228 5356
rect 35066 5302 35068 5354
rect 35130 5302 35142 5354
rect 35204 5302 35206 5354
rect 35044 5300 35068 5302
rect 35124 5300 35148 5302
rect 35204 5300 35228 5302
rect 34988 5280 35284 5300
rect 34870 5021 34922 5027
rect 34870 4963 34922 4969
rect 35350 5021 35402 5027
rect 35350 4963 35402 4969
rect 34882 3843 34910 4963
rect 34988 4024 35284 4044
rect 35044 4022 35068 4024
rect 35124 4022 35148 4024
rect 35204 4022 35228 4024
rect 35066 3970 35068 4022
rect 35130 3970 35142 4022
rect 35204 3970 35206 4022
rect 35044 3968 35068 3970
rect 35124 3968 35148 3970
rect 35204 3968 35228 3970
rect 34988 3948 35284 3968
rect 34870 3837 34922 3843
rect 34870 3779 34922 3785
rect 34966 3689 35018 3695
rect 34882 3649 34966 3677
rect 34882 1864 34910 3649
rect 34966 3631 35018 3637
rect 35362 3085 35390 4963
rect 35266 3057 35390 3085
rect 35266 2923 35294 3057
rect 35458 3048 35486 6369
rect 35542 3911 35594 3917
rect 35542 3853 35594 3859
rect 35554 3177 35582 3853
rect 35734 3689 35786 3695
rect 35734 3631 35786 3637
rect 35542 3171 35594 3177
rect 35542 3113 35594 3119
rect 35350 3023 35402 3029
rect 35458 3020 35678 3048
rect 35350 2965 35402 2971
rect 35252 2914 35308 2923
rect 35252 2849 35308 2858
rect 34988 2692 35284 2712
rect 35044 2690 35068 2692
rect 35124 2690 35148 2692
rect 35204 2690 35228 2692
rect 35066 2638 35068 2690
rect 35130 2638 35142 2690
rect 35204 2638 35206 2690
rect 35044 2636 35068 2638
rect 35124 2636 35148 2638
rect 35204 2636 35228 2638
rect 34988 2616 35284 2636
rect 35156 2470 35212 2479
rect 35156 2405 35212 2414
rect 34882 1836 35006 1864
rect 34870 1247 34922 1253
rect 34870 1189 34922 1195
rect 34882 800 34910 1189
rect 34978 800 35006 1836
rect 35170 800 35198 2405
rect 35362 1697 35390 2965
rect 35446 2949 35498 2955
rect 35446 2891 35498 2897
rect 35650 2894 35678 3020
rect 35350 1691 35402 1697
rect 35350 1633 35402 1639
rect 35458 1568 35486 2891
rect 35266 1540 35486 1568
rect 35554 2866 35678 2894
rect 35266 800 35294 1540
rect 35350 1395 35402 1401
rect 35350 1337 35402 1343
rect 35362 800 35390 1337
rect 35554 828 35582 2866
rect 35638 2579 35690 2585
rect 35638 2521 35690 2527
rect 35458 800 35582 828
rect 35650 800 35678 2521
rect 35746 800 35774 3631
rect 35842 800 35870 7405
rect 36226 7099 36254 9847
rect 36514 7913 36542 11549
rect 36982 9831 37034 9837
rect 36982 9773 37034 9779
rect 36790 9757 36842 9763
rect 36790 9699 36842 9705
rect 36802 9097 36830 9699
rect 36790 9091 36842 9097
rect 36790 9033 36842 9039
rect 36502 7907 36554 7913
rect 36502 7849 36554 7855
rect 36514 7765 36542 7849
rect 36502 7759 36554 7765
rect 36502 7701 36554 7707
rect 36598 7463 36650 7469
rect 36598 7405 36650 7411
rect 36214 7093 36266 7099
rect 36214 7035 36266 7041
rect 35926 6945 35978 6951
rect 35926 6887 35978 6893
rect 36406 6945 36458 6951
rect 36406 6887 36458 6893
rect 35938 3219 35966 6887
rect 36310 6353 36362 6359
rect 36310 6295 36362 6301
rect 36022 5687 36074 5693
rect 36022 5629 36074 5635
rect 36214 5687 36266 5693
rect 36214 5629 36266 5635
rect 35924 3210 35980 3219
rect 35924 3145 35980 3154
rect 35926 3097 35978 3103
rect 35926 3039 35978 3045
rect 35938 1253 35966 3039
rect 36034 2955 36062 5629
rect 36118 5021 36170 5027
rect 36118 4963 36170 4969
rect 36130 3103 36158 4963
rect 36118 3097 36170 3103
rect 36118 3039 36170 3045
rect 36022 2949 36074 2955
rect 36022 2891 36074 2897
rect 36226 2894 36254 5629
rect 36130 2866 36254 2894
rect 36130 1420 36158 2866
rect 36322 1697 36350 6295
rect 36310 1691 36362 1697
rect 36310 1633 36362 1639
rect 36418 1568 36446 6887
rect 36502 3689 36554 3695
rect 36502 3631 36554 3637
rect 36034 1392 36158 1420
rect 36226 1540 36446 1568
rect 35926 1247 35978 1253
rect 35926 1189 35978 1195
rect 36034 800 36062 1392
rect 36118 1321 36170 1327
rect 36118 1263 36170 1269
rect 36130 800 36158 1263
rect 36226 800 36254 1540
rect 36310 1395 36362 1401
rect 36310 1337 36362 1343
rect 36322 800 36350 1337
rect 36514 800 36542 3631
rect 36610 800 36638 7405
rect 36994 7099 37022 9773
rect 37462 7833 37514 7839
rect 37462 7775 37514 7781
rect 36982 7093 37034 7099
rect 36982 7035 37034 7041
rect 37474 7025 37502 7775
rect 37762 7099 37790 13769
rect 38038 7463 38090 7469
rect 38038 7405 38090 7411
rect 37750 7093 37802 7099
rect 37750 7035 37802 7041
rect 37462 7019 37514 7025
rect 37462 6961 37514 6967
rect 36982 6945 37034 6951
rect 36982 6887 37034 6893
rect 36886 6279 36938 6285
rect 36886 6221 36938 6227
rect 36898 6137 36926 6221
rect 36886 6131 36938 6137
rect 36886 6073 36938 6079
rect 36898 5619 36926 6073
rect 36886 5613 36938 5619
rect 36886 5555 36938 5561
rect 36886 5021 36938 5027
rect 36886 4963 36938 4969
rect 36790 4355 36842 4361
rect 36790 4297 36842 4303
rect 36694 3097 36746 3103
rect 36694 3039 36746 3045
rect 36706 800 36734 3039
rect 36802 800 36830 4297
rect 36898 2585 36926 4963
rect 36886 2579 36938 2585
rect 36886 2521 36938 2527
rect 36994 800 37022 6887
rect 37654 6797 37706 6803
rect 37654 6739 37706 6745
rect 37558 5687 37610 5693
rect 37558 5629 37610 5635
rect 37462 5613 37514 5619
rect 37462 5555 37514 5561
rect 37174 4281 37226 4287
rect 37174 4223 37226 4229
rect 37078 3171 37130 3177
rect 37078 3113 37130 3119
rect 37090 800 37118 3113
rect 37186 800 37214 4223
rect 37366 3541 37418 3547
rect 37366 3483 37418 3489
rect 37270 3023 37322 3029
rect 37270 2965 37322 2971
rect 37282 1327 37310 2965
rect 37270 1321 37322 1327
rect 37270 1263 37322 1269
rect 37378 800 37406 3483
rect 37474 800 37502 5555
rect 37570 3103 37598 5629
rect 37558 3097 37610 3103
rect 37558 3039 37610 3045
rect 37558 2949 37610 2955
rect 37558 2891 37610 2897
rect 37570 800 37598 2891
rect 37666 800 37694 6739
rect 37846 3837 37898 3843
rect 37846 3779 37898 3785
rect 37858 800 37886 3779
rect 37942 3689 37994 3695
rect 37942 3631 37994 3637
rect 37954 800 37982 3631
rect 38050 800 38078 7405
rect 38146 7173 38174 33379
rect 38230 30477 38282 30483
rect 38230 30419 38282 30425
rect 38242 19827 38270 30419
rect 38230 19821 38282 19827
rect 38230 19763 38282 19769
rect 38434 9615 38462 56171
rect 39106 55717 39134 59200
rect 39682 56901 39710 59200
rect 39670 56895 39722 56901
rect 39670 56837 39722 56843
rect 39766 56747 39818 56753
rect 39766 56689 39818 56695
rect 39574 56451 39626 56457
rect 39574 56393 39626 56399
rect 39094 55711 39146 55717
rect 39094 55653 39146 55659
rect 39190 55563 39242 55569
rect 39190 55505 39242 55511
rect 39094 24261 39146 24267
rect 39094 24203 39146 24209
rect 38422 9609 38474 9615
rect 38422 9551 38474 9557
rect 39106 7913 39134 24203
rect 39094 7907 39146 7913
rect 39094 7849 39146 7855
rect 38806 7759 38858 7765
rect 38806 7701 38858 7707
rect 38134 7167 38186 7173
rect 38134 7109 38186 7115
rect 38518 7167 38570 7173
rect 38518 7109 38570 7115
rect 38530 7044 38558 7109
rect 38434 7016 38558 7044
rect 38326 3097 38378 3103
rect 38326 3039 38378 3045
rect 38134 2949 38186 2955
rect 38134 2891 38186 2897
rect 38146 800 38174 2891
rect 38338 800 38366 3039
rect 38434 800 38462 7016
rect 38518 6945 38570 6951
rect 38518 6887 38570 6893
rect 38530 3547 38558 6887
rect 38614 5021 38666 5027
rect 38614 4963 38666 4969
rect 38518 3541 38570 3547
rect 38518 3483 38570 3489
rect 38518 3245 38570 3251
rect 38518 3187 38570 3193
rect 38530 800 38558 3187
rect 38626 3177 38654 4963
rect 38710 3689 38762 3695
rect 38710 3631 38762 3637
rect 38614 3171 38666 3177
rect 38614 3113 38666 3119
rect 38722 800 38750 3631
rect 38818 800 38846 7701
rect 39106 7691 39134 7849
rect 39094 7685 39146 7691
rect 39094 7627 39146 7633
rect 38998 7019 39050 7025
rect 38998 6961 39050 6967
rect 38902 6353 38954 6359
rect 38902 6295 38954 6301
rect 38914 800 38942 6295
rect 39010 5545 39038 6961
rect 39094 5687 39146 5693
rect 39094 5629 39146 5635
rect 38998 5539 39050 5545
rect 38998 5481 39050 5487
rect 38998 4355 39050 4361
rect 38998 4297 39050 4303
rect 39010 800 39038 4297
rect 39106 2955 39134 5629
rect 39202 3917 39230 55505
rect 39586 22935 39614 56393
rect 39670 47645 39722 47651
rect 39670 47587 39722 47593
rect 39574 22929 39626 22935
rect 39574 22871 39626 22877
rect 39478 7463 39530 7469
rect 39478 7405 39530 7411
rect 39286 5687 39338 5693
rect 39286 5629 39338 5635
rect 39190 3911 39242 3917
rect 39190 3853 39242 3859
rect 39094 2949 39146 2955
rect 39094 2891 39146 2897
rect 39190 2949 39242 2955
rect 39190 2891 39242 2897
rect 39202 800 39230 2891
rect 39298 800 39326 5629
rect 39382 5021 39434 5027
rect 39382 4963 39434 4969
rect 39394 3843 39422 4963
rect 39382 3837 39434 3843
rect 39382 3779 39434 3785
rect 39382 3541 39434 3547
rect 39382 3483 39434 3489
rect 39394 800 39422 3483
rect 39490 800 39518 7405
rect 39682 7173 39710 47587
rect 39778 16423 39806 56689
rect 40162 56531 40190 59200
rect 40438 56747 40490 56753
rect 40438 56689 40490 56695
rect 40150 56525 40202 56531
rect 40150 56467 40202 56473
rect 39862 56229 39914 56235
rect 39862 56171 39914 56177
rect 39766 16417 39818 16423
rect 39766 16359 39818 16365
rect 39874 15239 39902 56171
rect 40246 22411 40298 22417
rect 40246 22353 40298 22359
rect 39862 15233 39914 15239
rect 39862 15175 39914 15181
rect 40258 7932 40286 22353
rect 40450 10799 40478 56689
rect 40738 55717 40766 59200
rect 41218 56975 41246 59200
rect 41206 56969 41258 56975
rect 41206 56911 41258 56917
rect 40822 56747 40874 56753
rect 40822 56689 40874 56695
rect 40834 56087 40862 56689
rect 41794 56531 41822 59200
rect 42274 56531 42302 59200
rect 42850 56901 42878 59200
rect 42838 56895 42890 56901
rect 42838 56837 42890 56843
rect 42934 56747 42986 56753
rect 42934 56689 42986 56695
rect 41782 56525 41834 56531
rect 41782 56467 41834 56473
rect 42262 56525 42314 56531
rect 42262 56467 42314 56473
rect 42358 56377 42410 56383
rect 42358 56319 42410 56325
rect 42070 56229 42122 56235
rect 42070 56171 42122 56177
rect 40822 56081 40874 56087
rect 40822 56023 40874 56029
rect 40726 55711 40778 55717
rect 40726 55653 40778 55659
rect 40822 55563 40874 55569
rect 40822 55505 40874 55511
rect 40834 34849 40862 55505
rect 40918 50087 40970 50093
rect 40918 50029 40970 50035
rect 40822 34843 40874 34849
rect 40822 34785 40874 34791
rect 40930 13907 40958 50029
rect 42082 25229 42110 56171
rect 42370 55051 42398 56319
rect 42646 56229 42698 56235
rect 42646 56171 42698 56177
rect 42358 55045 42410 55051
rect 42358 54987 42410 54993
rect 42166 26925 42218 26931
rect 42166 26867 42218 26873
rect 42070 25223 42122 25229
rect 42070 25165 42122 25171
rect 41878 23891 41930 23897
rect 41878 23833 41930 23839
rect 40918 13901 40970 13907
rect 40918 13843 40970 13849
rect 41782 12125 41834 12131
rect 41782 12067 41834 12073
rect 41206 10867 41258 10873
rect 41206 10809 41258 10815
rect 40438 10793 40490 10799
rect 40438 10735 40490 10741
rect 40162 7913 40286 7932
rect 40162 7907 40298 7913
rect 40162 7904 40246 7907
rect 40162 7617 40190 7904
rect 40246 7849 40298 7855
rect 40246 7759 40298 7765
rect 40246 7701 40298 7707
rect 40150 7611 40202 7617
rect 40150 7553 40202 7559
rect 39670 7167 39722 7173
rect 39670 7109 39722 7115
rect 39862 6871 39914 6877
rect 39862 6813 39914 6819
rect 39574 5021 39626 5027
rect 39574 4963 39626 4969
rect 39586 3251 39614 4963
rect 39766 4355 39818 4361
rect 39766 4297 39818 4303
rect 39574 3245 39626 3251
rect 39574 3187 39626 3193
rect 39670 3171 39722 3177
rect 39670 3113 39722 3119
rect 39682 800 39710 3113
rect 39778 800 39806 4297
rect 39874 800 39902 6813
rect 39958 6131 40010 6137
rect 39958 6073 40010 6079
rect 39970 2955 39998 6073
rect 40054 3837 40106 3843
rect 40054 3779 40106 3785
rect 39958 2949 40010 2955
rect 39958 2891 40010 2897
rect 40066 800 40094 3779
rect 40150 3541 40202 3547
rect 40150 3483 40202 3489
rect 40162 800 40190 3483
rect 40258 800 40286 7701
rect 41110 6797 41162 6803
rect 41110 6739 41162 6745
rect 40342 6353 40394 6359
rect 40342 6295 40394 6301
rect 40354 800 40382 6295
rect 40630 6279 40682 6285
rect 40630 6221 40682 6227
rect 40534 3023 40586 3029
rect 40534 2965 40586 2971
rect 40546 800 40574 2965
rect 40642 800 40670 6221
rect 40822 6205 40874 6211
rect 40822 6147 40874 6153
rect 40726 5687 40778 5693
rect 40726 5629 40778 5635
rect 40738 800 40766 5629
rect 40834 3103 40862 6147
rect 40918 5021 40970 5027
rect 40918 4963 40970 4969
rect 40930 3177 40958 4963
rect 41014 3689 41066 3695
rect 41014 3631 41066 3637
rect 40918 3171 40970 3177
rect 40918 3113 40970 3119
rect 40822 3097 40874 3103
rect 40822 3039 40874 3045
rect 41026 2894 41054 3631
rect 41122 3344 41150 6739
rect 41218 6433 41246 10809
rect 41794 7765 41822 12067
rect 41782 7759 41834 7765
rect 41782 7701 41834 7707
rect 41782 7463 41834 7469
rect 41782 7405 41834 7411
rect 41302 6575 41354 6581
rect 41302 6517 41354 6523
rect 41206 6427 41258 6433
rect 41206 6369 41258 6375
rect 41122 3316 41246 3344
rect 41218 3251 41246 3316
rect 41206 3245 41258 3251
rect 41206 3187 41258 3193
rect 41110 3171 41162 3177
rect 41110 3113 41162 3119
rect 40822 2875 40874 2881
rect 40822 2817 40874 2823
rect 40930 2866 41054 2894
rect 40834 2511 40862 2817
rect 40822 2505 40874 2511
rect 40822 2447 40874 2453
rect 40930 800 40958 2866
rect 41014 1469 41066 1475
rect 41014 1411 41066 1417
rect 41026 800 41054 1411
rect 41122 800 41150 3113
rect 41206 3097 41258 3103
rect 41206 3039 41258 3045
rect 41218 800 41246 3039
rect 41314 1475 41342 6517
rect 41686 5021 41738 5027
rect 41686 4963 41738 4969
rect 41698 3843 41726 4963
rect 41686 3837 41738 3843
rect 41686 3779 41738 3785
rect 41794 3640 41822 7405
rect 41890 7173 41918 23833
rect 42178 8579 42206 26867
rect 42658 17163 42686 56171
rect 42742 27517 42794 27523
rect 42742 27459 42794 27465
rect 42646 17157 42698 17163
rect 42646 17099 42698 17105
rect 42166 8573 42218 8579
rect 42166 8515 42218 8521
rect 42178 8431 42206 8515
rect 42166 8425 42218 8431
rect 42166 8367 42218 8373
rect 42754 7765 42782 27459
rect 42838 18267 42890 18273
rect 42838 18209 42890 18215
rect 42850 16571 42878 18209
rect 42946 17829 42974 56689
rect 43330 56531 43358 59200
rect 43906 56531 43934 59200
rect 44386 56901 44414 59200
rect 44374 56895 44426 56901
rect 44374 56837 44426 56843
rect 44758 56747 44810 56753
rect 44758 56689 44810 56695
rect 43318 56525 43370 56531
rect 43318 56467 43370 56473
rect 43894 56525 43946 56531
rect 43894 56467 43946 56473
rect 43894 56303 43946 56309
rect 43894 56245 43946 56251
rect 43510 56229 43562 56235
rect 43510 56171 43562 56177
rect 43522 48761 43550 56171
rect 43510 48755 43562 48761
rect 43510 48697 43562 48703
rect 43906 46911 43934 56245
rect 44182 56229 44234 56235
rect 44182 56171 44234 56177
rect 43894 46905 43946 46911
rect 43894 46847 43946 46853
rect 44086 28923 44138 28929
rect 44086 28865 44138 28871
rect 43894 20117 43946 20123
rect 43894 20059 43946 20065
rect 42934 17823 42986 17829
rect 42934 17765 42986 17771
rect 42838 16565 42890 16571
rect 42838 16507 42890 16513
rect 42838 14197 42890 14203
rect 42838 14139 42890 14145
rect 42742 7759 42794 7765
rect 42742 7701 42794 7707
rect 42454 7463 42506 7469
rect 42454 7405 42506 7411
rect 41878 7167 41930 7173
rect 41878 7109 41930 7115
rect 42262 7167 42314 7173
rect 42262 7109 42314 7115
rect 41890 6951 41918 7109
rect 41878 6945 41930 6951
rect 41878 6887 41930 6893
rect 42274 6581 42302 7109
rect 42262 6575 42314 6581
rect 42262 6517 42314 6523
rect 41878 6353 41930 6359
rect 41878 6295 41930 6301
rect 41410 3612 41822 3640
rect 41302 1469 41354 1475
rect 41302 1411 41354 1417
rect 41410 800 41438 3612
rect 41590 3541 41642 3547
rect 41590 3483 41642 3489
rect 41494 2949 41546 2955
rect 41494 2891 41546 2897
rect 41506 800 41534 2891
rect 41602 800 41630 3483
rect 41686 3245 41738 3251
rect 41686 3187 41738 3193
rect 41698 800 41726 3187
rect 41890 800 41918 6295
rect 42070 5687 42122 5693
rect 42070 5629 42122 5635
rect 42262 5687 42314 5693
rect 42262 5629 42314 5635
rect 41974 4355 42026 4361
rect 41974 4297 42026 4303
rect 41986 800 42014 4297
rect 42082 2955 42110 5629
rect 42166 5021 42218 5027
rect 42166 4963 42218 4969
rect 42178 3177 42206 4963
rect 42166 3171 42218 3177
rect 42166 3113 42218 3119
rect 42166 3023 42218 3029
rect 42166 2965 42218 2971
rect 42070 2949 42122 2955
rect 42070 2891 42122 2897
rect 42178 976 42206 2965
rect 42082 948 42206 976
rect 42082 800 42110 948
rect 42274 800 42302 5629
rect 42358 4355 42410 4361
rect 42358 4297 42410 4303
rect 42370 800 42398 4297
rect 42466 800 42494 7405
rect 42850 6433 42878 14139
rect 43702 13235 43754 13241
rect 43702 13177 43754 13183
rect 43030 8943 43082 8949
rect 43030 8885 43082 8891
rect 43042 7099 43070 8885
rect 43510 7167 43562 7173
rect 43510 7109 43562 7115
rect 43030 7093 43082 7099
rect 43030 7035 43082 7041
rect 43414 7093 43466 7099
rect 43414 7035 43466 7041
rect 43426 6803 43454 7035
rect 43414 6797 43466 6803
rect 43414 6739 43466 6745
rect 42838 6427 42890 6433
rect 42838 6369 42890 6375
rect 42646 6205 42698 6211
rect 42646 6147 42698 6153
rect 42658 3029 42686 6147
rect 43426 5767 43454 6739
rect 43414 5761 43466 5767
rect 43414 5703 43466 5709
rect 43222 5687 43274 5693
rect 43222 5629 43274 5635
rect 42838 3763 42890 3769
rect 42838 3705 42890 3711
rect 42742 3689 42794 3695
rect 42742 3631 42794 3637
rect 42646 3023 42698 3029
rect 42646 2965 42698 2971
rect 42550 2949 42602 2955
rect 42550 2891 42602 2897
rect 42562 800 42590 2891
rect 42754 800 42782 3631
rect 42850 800 42878 3705
rect 43234 3159 43262 5629
rect 43318 5021 43370 5027
rect 43318 4963 43370 4969
rect 42946 3131 43262 3159
rect 42946 800 42974 3131
rect 43222 3097 43274 3103
rect 43222 3039 43274 3045
rect 43030 3023 43082 3029
rect 43030 2965 43082 2971
rect 43042 800 43070 2965
rect 43234 2752 43262 3039
rect 43330 2955 43358 4963
rect 43414 4355 43466 4361
rect 43414 4297 43466 4303
rect 43318 2949 43370 2955
rect 43318 2891 43370 2897
rect 43426 2752 43454 4297
rect 43522 4213 43550 7109
rect 43714 7044 43742 13177
rect 43906 7691 43934 20059
rect 43990 19747 44042 19753
rect 43990 19689 44042 19695
rect 44002 7765 44030 19689
rect 43990 7759 44042 7765
rect 43990 7701 44042 7707
rect 43894 7685 43946 7691
rect 43894 7627 43946 7633
rect 43894 7463 43946 7469
rect 43894 7405 43946 7411
rect 43798 7093 43850 7099
rect 43714 7041 43798 7044
rect 43714 7035 43850 7041
rect 43714 7016 43838 7035
rect 43798 6945 43850 6951
rect 43798 6887 43850 6893
rect 43606 6871 43658 6877
rect 43606 6813 43658 6819
rect 43510 4207 43562 4213
rect 43510 4149 43562 4155
rect 43234 2724 43358 2752
rect 43426 2724 43550 2752
rect 43222 2579 43274 2585
rect 43222 2521 43274 2527
rect 43234 800 43262 2521
rect 43330 800 43358 2724
rect 43522 2160 43550 2724
rect 43426 2132 43550 2160
rect 43426 800 43454 2132
rect 43618 800 43646 6813
rect 43702 5687 43754 5693
rect 43702 5629 43754 5635
rect 43714 800 43742 5629
rect 43810 3769 43838 6887
rect 43798 3763 43850 3769
rect 43798 3705 43850 3711
rect 43798 3615 43850 3621
rect 43798 3557 43850 3563
rect 43810 800 43838 3557
rect 43906 800 43934 7405
rect 44098 6433 44126 28865
rect 44194 12353 44222 56171
rect 44374 36101 44426 36107
rect 44374 36043 44426 36049
rect 44182 12347 44234 12353
rect 44182 12289 44234 12295
rect 44386 8505 44414 36043
rect 44662 20783 44714 20789
rect 44662 20725 44714 20731
rect 44374 8499 44426 8505
rect 44374 8441 44426 8447
rect 44278 6797 44330 6803
rect 44278 6739 44330 6745
rect 44086 6427 44138 6433
rect 44086 6369 44138 6375
rect 44086 6131 44138 6137
rect 44086 6073 44138 6079
rect 44098 3344 44126 6073
rect 44002 3316 44126 3344
rect 44002 2585 44030 3316
rect 44086 3245 44138 3251
rect 44086 3187 44138 3193
rect 43990 2579 44042 2585
rect 43990 2521 44042 2527
rect 44098 800 44126 3187
rect 44182 2949 44234 2955
rect 44182 2891 44234 2897
rect 44194 800 44222 2891
rect 44290 800 44318 6739
rect 44674 6433 44702 20725
rect 44770 17755 44798 56689
rect 44962 56531 44990 59200
rect 44950 56525 45002 56531
rect 44950 56467 45002 56473
rect 45442 55717 45470 59200
rect 45922 56901 45950 59200
rect 45910 56895 45962 56901
rect 45910 56837 45962 56843
rect 46102 56747 46154 56753
rect 46102 56689 46154 56695
rect 45430 55711 45482 55717
rect 45430 55653 45482 55659
rect 45334 55637 45386 55643
rect 45334 55579 45386 55585
rect 44854 49421 44906 49427
rect 44854 49363 44906 49369
rect 44758 17749 44810 17755
rect 44758 17691 44810 17697
rect 44758 12125 44810 12131
rect 44758 12067 44810 12073
rect 44770 11761 44798 12067
rect 44866 11761 44894 49363
rect 45046 19821 45098 19827
rect 45046 19763 45098 19769
rect 44758 11755 44810 11761
rect 44758 11697 44810 11703
rect 44854 11755 44906 11761
rect 44854 11697 44906 11703
rect 44758 10793 44810 10799
rect 44758 10735 44810 10741
rect 44770 7913 44798 10735
rect 44950 8795 45002 8801
rect 44950 8737 45002 8743
rect 44758 7907 44810 7913
rect 44758 7849 44810 7855
rect 44758 7463 44810 7469
rect 44758 7405 44810 7411
rect 44662 6427 44714 6433
rect 44662 6369 44714 6375
rect 44662 5687 44714 5693
rect 44662 5629 44714 5635
rect 44674 3936 44702 5629
rect 44482 3908 44702 3936
rect 44482 800 44510 3908
rect 44566 3763 44618 3769
rect 44566 3705 44618 3711
rect 44578 800 44606 3705
rect 44770 3529 44798 7405
rect 44962 7173 44990 8737
rect 45058 7765 45086 19763
rect 45346 12131 45374 55579
rect 45814 55415 45866 55421
rect 45814 55357 45866 55363
rect 45430 46757 45482 46763
rect 45430 46699 45482 46705
rect 45442 23823 45470 46699
rect 45622 28109 45674 28115
rect 45622 28051 45674 28057
rect 45430 23817 45482 23823
rect 45430 23759 45482 23765
rect 45334 12125 45386 12131
rect 45334 12067 45386 12073
rect 45634 7765 45662 28051
rect 45826 19679 45854 55357
rect 45814 19673 45866 19679
rect 45814 19615 45866 19621
rect 45814 18119 45866 18125
rect 45814 18061 45866 18067
rect 45826 17533 45854 18061
rect 46114 17681 46142 56689
rect 46498 56531 46526 59200
rect 46486 56525 46538 56531
rect 46486 56467 46538 56473
rect 46870 56303 46922 56309
rect 46870 56245 46922 56251
rect 46678 56229 46730 56235
rect 46678 56171 46730 56177
rect 46102 17675 46154 17681
rect 46102 17617 46154 17623
rect 45814 17527 45866 17533
rect 45814 17469 45866 17475
rect 46690 14129 46718 56171
rect 46882 40547 46910 56245
rect 46978 55717 47006 59200
rect 47554 56975 47582 59200
rect 47542 56969 47594 56975
rect 47542 56911 47594 56917
rect 48034 56531 48062 59200
rect 48610 56531 48638 59200
rect 49090 56901 49118 59200
rect 49078 56895 49130 56901
rect 49078 56837 49130 56843
rect 48694 56747 48746 56753
rect 48694 56689 48746 56695
rect 48022 56525 48074 56531
rect 48022 56467 48074 56473
rect 48598 56525 48650 56531
rect 48598 56467 48650 56473
rect 47062 56377 47114 56383
rect 47062 56319 47114 56325
rect 46966 55711 47018 55717
rect 46966 55653 47018 55659
rect 47074 47534 47102 56319
rect 48214 56229 48266 56235
rect 48214 56171 48266 56177
rect 48598 56229 48650 56235
rect 48598 56171 48650 56177
rect 48118 49421 48170 49427
rect 48118 49363 48170 49369
rect 46978 47506 47102 47534
rect 46978 46097 47006 47506
rect 46966 46091 47018 46097
rect 46966 46033 47018 46039
rect 47734 44093 47786 44099
rect 47734 44035 47786 44041
rect 47746 43877 47774 44035
rect 47734 43871 47786 43877
rect 47734 43813 47786 43819
rect 46870 40541 46922 40547
rect 46870 40483 46922 40489
rect 46678 14123 46730 14129
rect 46678 14065 46730 14071
rect 48022 8277 48074 8283
rect 48022 8219 48074 8225
rect 45046 7759 45098 7765
rect 45046 7701 45098 7707
rect 45622 7759 45674 7765
rect 45622 7701 45674 7707
rect 45814 7759 45866 7765
rect 45814 7701 45866 7707
rect 46486 7759 46538 7765
rect 46486 7701 46538 7707
rect 45046 7463 45098 7469
rect 45046 7405 45098 7411
rect 44950 7167 45002 7173
rect 44950 7109 45002 7115
rect 44854 5021 44906 5027
rect 44854 4963 44906 4969
rect 44674 3501 44798 3529
rect 44674 800 44702 3501
rect 44866 3177 44894 4963
rect 44950 4355 45002 4361
rect 44950 4297 45002 4303
rect 44854 3171 44906 3177
rect 44854 3113 44906 3119
rect 44758 3097 44810 3103
rect 44758 3039 44810 3045
rect 44770 800 44798 3039
rect 44962 800 44990 4297
rect 45058 800 45086 7405
rect 45430 6945 45482 6951
rect 45346 6905 45430 6933
rect 45238 3615 45290 3621
rect 45238 3557 45290 3563
rect 45142 3171 45194 3177
rect 45142 3113 45194 3119
rect 45154 800 45182 3113
rect 45250 800 45278 3557
rect 45346 3159 45374 6905
rect 45430 6887 45482 6893
rect 45526 6353 45578 6359
rect 45526 6295 45578 6301
rect 45430 5021 45482 5027
rect 45430 4963 45482 4969
rect 45442 3251 45470 4963
rect 45430 3245 45482 3251
rect 45430 3187 45482 3193
rect 45346 3131 45470 3159
rect 45442 800 45470 3131
rect 45538 800 45566 6295
rect 45622 3023 45674 3029
rect 45622 2965 45674 2971
rect 45634 800 45662 2965
rect 45826 800 45854 7701
rect 46102 5687 46154 5693
rect 46102 5629 46154 5635
rect 46114 3640 46142 5629
rect 46198 5021 46250 5027
rect 46198 4963 46250 4969
rect 46294 5021 46346 5027
rect 46294 4963 46346 4969
rect 45922 3612 46142 3640
rect 45922 800 45950 3612
rect 46006 3541 46058 3547
rect 46006 3483 46058 3489
rect 46018 800 46046 3483
rect 46210 3103 46238 4963
rect 46306 3177 46334 4963
rect 46294 3171 46346 3177
rect 46294 3113 46346 3119
rect 46198 3097 46250 3103
rect 46198 3039 46250 3045
rect 46390 3097 46442 3103
rect 46390 3039 46442 3045
rect 46294 2949 46346 2955
rect 46294 2891 46346 2897
rect 46102 2801 46154 2807
rect 46102 2743 46154 2749
rect 46114 800 46142 2743
rect 46306 800 46334 2891
rect 46402 800 46430 3039
rect 46498 800 46526 7701
rect 47926 7611 47978 7617
rect 47926 7553 47978 7559
rect 47254 7463 47306 7469
rect 47254 7405 47306 7411
rect 46774 6945 46826 6951
rect 46774 6887 46826 6893
rect 46678 5687 46730 5693
rect 46594 5647 46678 5675
rect 46594 800 46622 5647
rect 46678 5629 46730 5635
rect 46786 4528 46814 6887
rect 46870 6871 46922 6877
rect 46870 6813 46922 6819
rect 46690 4500 46814 4528
rect 46690 2807 46718 4500
rect 46774 4355 46826 4361
rect 46774 4297 46826 4303
rect 46678 2801 46730 2807
rect 46678 2743 46730 2749
rect 46786 800 46814 4297
rect 46882 800 46910 6813
rect 46966 6353 47018 6359
rect 46966 6295 47018 6301
rect 46978 800 47006 6295
rect 47158 3689 47210 3695
rect 47158 3631 47210 3637
rect 47170 800 47198 3631
rect 47266 800 47294 7405
rect 47938 7247 47966 7553
rect 47926 7241 47978 7247
rect 47926 7183 47978 7189
rect 47734 6353 47786 6359
rect 47734 6295 47786 6301
rect 47542 5687 47594 5693
rect 47542 5629 47594 5635
rect 47554 4380 47582 5629
rect 47638 5021 47690 5027
rect 47638 4963 47690 4969
rect 47362 4352 47582 4380
rect 47362 800 47390 4352
rect 47446 4281 47498 4287
rect 47446 4223 47498 4229
rect 47458 800 47486 4223
rect 47542 3541 47594 3547
rect 47542 3483 47594 3489
rect 47554 2752 47582 3483
rect 47650 2955 47678 4963
rect 47638 2949 47690 2955
rect 47638 2891 47690 2897
rect 47554 2724 47678 2752
rect 47650 800 47678 2724
rect 47746 800 47774 6295
rect 47830 4355 47882 4361
rect 47830 4297 47882 4303
rect 47842 800 47870 4297
rect 48034 800 48062 8219
rect 48130 7543 48158 49363
rect 48226 47577 48254 56171
rect 48214 47571 48266 47577
rect 48214 47513 48266 47519
rect 48310 40911 48362 40917
rect 48310 40853 48362 40859
rect 48118 7537 48170 7543
rect 48118 7479 48170 7485
rect 48322 7099 48350 40853
rect 48610 18495 48638 56171
rect 48706 19235 48734 56689
rect 49666 56531 49694 59200
rect 50146 56531 50174 59200
rect 50722 56901 50750 59200
rect 50710 56895 50762 56901
rect 50710 56837 50762 56843
rect 50806 56747 50858 56753
rect 50806 56689 50858 56695
rect 50348 56638 50644 56658
rect 50404 56636 50428 56638
rect 50484 56636 50508 56638
rect 50564 56636 50588 56638
rect 50426 56584 50428 56636
rect 50490 56584 50502 56636
rect 50564 56584 50566 56636
rect 50404 56582 50428 56584
rect 50484 56582 50508 56584
rect 50564 56582 50588 56584
rect 50348 56562 50644 56582
rect 49654 56525 49706 56531
rect 49654 56467 49706 56473
rect 50134 56525 50186 56531
rect 50134 56467 50186 56473
rect 50230 56229 50282 56235
rect 50230 56171 50282 56177
rect 48886 48089 48938 48095
rect 48886 48031 48938 48037
rect 48694 19229 48746 19235
rect 48694 19171 48746 19177
rect 48598 18489 48650 18495
rect 48598 18431 48650 18437
rect 48598 17083 48650 17089
rect 48598 17025 48650 17031
rect 48610 8579 48638 17025
rect 48790 10867 48842 10873
rect 48790 10809 48842 10815
rect 48694 10275 48746 10281
rect 48694 10217 48746 10223
rect 48706 9171 48734 10217
rect 48694 9165 48746 9171
rect 48694 9107 48746 9113
rect 48598 8573 48650 8579
rect 48598 8515 48650 8521
rect 48610 8283 48638 8515
rect 48802 8357 48830 10809
rect 48898 8431 48926 48031
rect 50134 31883 50186 31889
rect 50134 31825 50186 31831
rect 49078 29441 49130 29447
rect 49078 29383 49130 29389
rect 48886 8425 48938 8431
rect 48886 8367 48938 8373
rect 48790 8351 48842 8357
rect 48790 8293 48842 8299
rect 48598 8277 48650 8283
rect 48598 8219 48650 8225
rect 48694 8203 48746 8209
rect 48694 8145 48746 8151
rect 48406 7463 48458 7469
rect 48406 7405 48458 7411
rect 48310 7093 48362 7099
rect 48310 7035 48362 7041
rect 48310 6945 48362 6951
rect 48310 6887 48362 6893
rect 48214 3689 48266 3695
rect 48214 3631 48266 3637
rect 48118 3171 48170 3177
rect 48118 3113 48170 3119
rect 48130 800 48158 3113
rect 48226 800 48254 3631
rect 48322 3547 48350 6887
rect 48310 3541 48362 3547
rect 48310 3483 48362 3489
rect 48418 1864 48446 7405
rect 48598 4281 48650 4287
rect 48598 4223 48650 4229
rect 48502 3245 48554 3251
rect 48502 3187 48554 3193
rect 48322 1836 48446 1864
rect 48322 800 48350 1836
rect 48514 800 48542 3187
rect 48610 800 48638 4223
rect 48706 800 48734 8145
rect 49090 7099 49118 29383
rect 49366 29219 49418 29225
rect 49366 29161 49418 29167
rect 49378 7765 49406 29161
rect 49654 20117 49706 20123
rect 49654 20059 49706 20065
rect 49558 16121 49610 16127
rect 49558 16063 49610 16069
rect 49570 15905 49598 16063
rect 49558 15899 49610 15905
rect 49558 15841 49610 15847
rect 49666 9689 49694 20059
rect 49654 9683 49706 9689
rect 49654 9625 49706 9631
rect 49462 8277 49514 8283
rect 49462 8219 49514 8225
rect 49366 7759 49418 7765
rect 49366 7701 49418 7707
rect 49174 7537 49226 7543
rect 49174 7479 49226 7485
rect 49078 7093 49130 7099
rect 49078 7035 49130 7041
rect 48790 6353 48842 6359
rect 48790 6295 48842 6301
rect 48802 800 48830 6295
rect 48982 5687 49034 5693
rect 48982 5629 49034 5635
rect 48994 3177 49022 5629
rect 49186 3640 49214 7479
rect 49366 5021 49418 5027
rect 49366 4963 49418 4969
rect 49270 3837 49322 3843
rect 49270 3779 49322 3785
rect 49090 3612 49214 3640
rect 48982 3171 49034 3177
rect 48982 3113 49034 3119
rect 48982 2949 49034 2955
rect 48982 2891 49034 2897
rect 48994 800 49022 2891
rect 49090 800 49118 3612
rect 49282 2900 49310 3779
rect 49186 2872 49310 2900
rect 49186 800 49214 2872
rect 49378 800 49406 4963
rect 49474 800 49502 8219
rect 50146 7099 50174 31825
rect 50242 9541 50270 56171
rect 50348 55306 50644 55326
rect 50404 55304 50428 55306
rect 50484 55304 50508 55306
rect 50564 55304 50588 55306
rect 50426 55252 50428 55304
rect 50490 55252 50502 55304
rect 50564 55252 50566 55304
rect 50404 55250 50428 55252
rect 50484 55250 50508 55252
rect 50564 55250 50588 55252
rect 50348 55230 50644 55250
rect 50348 53974 50644 53994
rect 50404 53972 50428 53974
rect 50484 53972 50508 53974
rect 50564 53972 50588 53974
rect 50426 53920 50428 53972
rect 50490 53920 50502 53972
rect 50564 53920 50566 53972
rect 50404 53918 50428 53920
rect 50484 53918 50508 53920
rect 50564 53918 50588 53920
rect 50348 53898 50644 53918
rect 50348 52642 50644 52662
rect 50404 52640 50428 52642
rect 50484 52640 50508 52642
rect 50564 52640 50588 52642
rect 50426 52588 50428 52640
rect 50490 52588 50502 52640
rect 50564 52588 50566 52640
rect 50404 52586 50428 52588
rect 50484 52586 50508 52588
rect 50564 52586 50588 52588
rect 50348 52566 50644 52586
rect 50348 51310 50644 51330
rect 50404 51308 50428 51310
rect 50484 51308 50508 51310
rect 50564 51308 50588 51310
rect 50426 51256 50428 51308
rect 50490 51256 50502 51308
rect 50564 51256 50566 51308
rect 50404 51254 50428 51256
rect 50484 51254 50508 51256
rect 50564 51254 50588 51256
rect 50348 51234 50644 51254
rect 50348 49978 50644 49998
rect 50404 49976 50428 49978
rect 50484 49976 50508 49978
rect 50564 49976 50588 49978
rect 50426 49924 50428 49976
rect 50490 49924 50502 49976
rect 50564 49924 50566 49976
rect 50404 49922 50428 49924
rect 50484 49922 50508 49924
rect 50564 49922 50588 49924
rect 50348 49902 50644 49922
rect 50348 48646 50644 48666
rect 50404 48644 50428 48646
rect 50484 48644 50508 48646
rect 50564 48644 50588 48646
rect 50426 48592 50428 48644
rect 50490 48592 50502 48644
rect 50564 48592 50566 48644
rect 50404 48590 50428 48592
rect 50484 48590 50508 48592
rect 50564 48590 50588 48592
rect 50348 48570 50644 48590
rect 50348 47314 50644 47334
rect 50404 47312 50428 47314
rect 50484 47312 50508 47314
rect 50564 47312 50588 47314
rect 50426 47260 50428 47312
rect 50490 47260 50502 47312
rect 50564 47260 50566 47312
rect 50404 47258 50428 47260
rect 50484 47258 50508 47260
rect 50564 47258 50588 47260
rect 50348 47238 50644 47258
rect 50348 45982 50644 46002
rect 50404 45980 50428 45982
rect 50484 45980 50508 45982
rect 50564 45980 50588 45982
rect 50426 45928 50428 45980
rect 50490 45928 50502 45980
rect 50564 45928 50566 45980
rect 50404 45926 50428 45928
rect 50484 45926 50508 45928
rect 50564 45926 50588 45928
rect 50348 45906 50644 45926
rect 50348 44650 50644 44670
rect 50404 44648 50428 44650
rect 50484 44648 50508 44650
rect 50564 44648 50588 44650
rect 50426 44596 50428 44648
rect 50490 44596 50502 44648
rect 50564 44596 50566 44648
rect 50404 44594 50428 44596
rect 50484 44594 50508 44596
rect 50564 44594 50588 44596
rect 50348 44574 50644 44594
rect 50348 43318 50644 43338
rect 50404 43316 50428 43318
rect 50484 43316 50508 43318
rect 50564 43316 50588 43318
rect 50426 43264 50428 43316
rect 50490 43264 50502 43316
rect 50564 43264 50566 43316
rect 50404 43262 50428 43264
rect 50484 43262 50508 43264
rect 50564 43262 50588 43264
rect 50348 43242 50644 43262
rect 50348 41986 50644 42006
rect 50404 41984 50428 41986
rect 50484 41984 50508 41986
rect 50564 41984 50588 41986
rect 50426 41932 50428 41984
rect 50490 41932 50502 41984
rect 50564 41932 50566 41984
rect 50404 41930 50428 41932
rect 50484 41930 50508 41932
rect 50564 41930 50588 41932
rect 50348 41910 50644 41930
rect 50348 40654 50644 40674
rect 50404 40652 50428 40654
rect 50484 40652 50508 40654
rect 50564 40652 50588 40654
rect 50426 40600 50428 40652
rect 50490 40600 50502 40652
rect 50564 40600 50566 40652
rect 50404 40598 50428 40600
rect 50484 40598 50508 40600
rect 50564 40598 50588 40600
rect 50348 40578 50644 40598
rect 50348 39322 50644 39342
rect 50404 39320 50428 39322
rect 50484 39320 50508 39322
rect 50564 39320 50588 39322
rect 50426 39268 50428 39320
rect 50490 39268 50502 39320
rect 50564 39268 50566 39320
rect 50404 39266 50428 39268
rect 50484 39266 50508 39268
rect 50564 39266 50588 39268
rect 50348 39246 50644 39266
rect 50348 37990 50644 38010
rect 50404 37988 50428 37990
rect 50484 37988 50508 37990
rect 50564 37988 50588 37990
rect 50426 37936 50428 37988
rect 50490 37936 50502 37988
rect 50564 37936 50566 37988
rect 50404 37934 50428 37936
rect 50484 37934 50508 37936
rect 50564 37934 50588 37936
rect 50348 37914 50644 37934
rect 50348 36658 50644 36678
rect 50404 36656 50428 36658
rect 50484 36656 50508 36658
rect 50564 36656 50588 36658
rect 50426 36604 50428 36656
rect 50490 36604 50502 36656
rect 50564 36604 50566 36656
rect 50404 36602 50428 36604
rect 50484 36602 50508 36604
rect 50564 36602 50588 36604
rect 50348 36582 50644 36602
rect 50348 35326 50644 35346
rect 50404 35324 50428 35326
rect 50484 35324 50508 35326
rect 50564 35324 50588 35326
rect 50426 35272 50428 35324
rect 50490 35272 50502 35324
rect 50564 35272 50566 35324
rect 50404 35270 50428 35272
rect 50484 35270 50508 35272
rect 50564 35270 50588 35272
rect 50348 35250 50644 35270
rect 50348 33994 50644 34014
rect 50404 33992 50428 33994
rect 50484 33992 50508 33994
rect 50564 33992 50588 33994
rect 50426 33940 50428 33992
rect 50490 33940 50502 33992
rect 50564 33940 50566 33992
rect 50404 33938 50428 33940
rect 50484 33938 50508 33940
rect 50564 33938 50588 33940
rect 50348 33918 50644 33938
rect 50348 32662 50644 32682
rect 50404 32660 50428 32662
rect 50484 32660 50508 32662
rect 50564 32660 50588 32662
rect 50426 32608 50428 32660
rect 50490 32608 50502 32660
rect 50564 32608 50566 32660
rect 50404 32606 50428 32608
rect 50484 32606 50508 32608
rect 50564 32606 50588 32608
rect 50348 32586 50644 32606
rect 50348 31330 50644 31350
rect 50404 31328 50428 31330
rect 50484 31328 50508 31330
rect 50564 31328 50588 31330
rect 50426 31276 50428 31328
rect 50490 31276 50502 31328
rect 50564 31276 50566 31328
rect 50404 31274 50428 31276
rect 50484 31274 50508 31276
rect 50564 31274 50588 31276
rect 50348 31254 50644 31274
rect 50348 29998 50644 30018
rect 50404 29996 50428 29998
rect 50484 29996 50508 29998
rect 50564 29996 50588 29998
rect 50426 29944 50428 29996
rect 50490 29944 50502 29996
rect 50564 29944 50566 29996
rect 50404 29942 50428 29944
rect 50484 29942 50508 29944
rect 50564 29942 50588 29944
rect 50348 29922 50644 29942
rect 50348 28666 50644 28686
rect 50404 28664 50428 28666
rect 50484 28664 50508 28666
rect 50564 28664 50588 28666
rect 50426 28612 50428 28664
rect 50490 28612 50502 28664
rect 50564 28612 50566 28664
rect 50404 28610 50428 28612
rect 50484 28610 50508 28612
rect 50564 28610 50588 28612
rect 50348 28590 50644 28610
rect 50348 27334 50644 27354
rect 50404 27332 50428 27334
rect 50484 27332 50508 27334
rect 50564 27332 50588 27334
rect 50426 27280 50428 27332
rect 50490 27280 50502 27332
rect 50564 27280 50566 27332
rect 50404 27278 50428 27280
rect 50484 27278 50508 27280
rect 50564 27278 50588 27280
rect 50348 27258 50644 27278
rect 50348 26002 50644 26022
rect 50404 26000 50428 26002
rect 50484 26000 50508 26002
rect 50564 26000 50588 26002
rect 50426 25948 50428 26000
rect 50490 25948 50502 26000
rect 50564 25948 50566 26000
rect 50404 25946 50428 25948
rect 50484 25946 50508 25948
rect 50564 25946 50588 25948
rect 50348 25926 50644 25946
rect 50710 24927 50762 24933
rect 50710 24869 50762 24875
rect 50348 24670 50644 24690
rect 50404 24668 50428 24670
rect 50484 24668 50508 24670
rect 50564 24668 50588 24670
rect 50426 24616 50428 24668
rect 50490 24616 50502 24668
rect 50564 24616 50566 24668
rect 50404 24614 50428 24616
rect 50484 24614 50508 24616
rect 50564 24614 50588 24616
rect 50348 24594 50644 24614
rect 50348 23338 50644 23358
rect 50404 23336 50428 23338
rect 50484 23336 50508 23338
rect 50564 23336 50588 23338
rect 50426 23284 50428 23336
rect 50490 23284 50502 23336
rect 50564 23284 50566 23336
rect 50404 23282 50428 23284
rect 50484 23282 50508 23284
rect 50564 23282 50588 23284
rect 50348 23262 50644 23282
rect 50348 22006 50644 22026
rect 50404 22004 50428 22006
rect 50484 22004 50508 22006
rect 50564 22004 50588 22006
rect 50426 21952 50428 22004
rect 50490 21952 50502 22004
rect 50564 21952 50566 22004
rect 50404 21950 50428 21952
rect 50484 21950 50508 21952
rect 50564 21950 50588 21952
rect 50348 21930 50644 21950
rect 50348 20674 50644 20694
rect 50404 20672 50428 20674
rect 50484 20672 50508 20674
rect 50564 20672 50588 20674
rect 50426 20620 50428 20672
rect 50490 20620 50502 20672
rect 50564 20620 50566 20672
rect 50404 20618 50428 20620
rect 50484 20618 50508 20620
rect 50564 20618 50588 20620
rect 50348 20598 50644 20618
rect 50348 19342 50644 19362
rect 50404 19340 50428 19342
rect 50484 19340 50508 19342
rect 50564 19340 50588 19342
rect 50426 19288 50428 19340
rect 50490 19288 50502 19340
rect 50564 19288 50566 19340
rect 50404 19286 50428 19288
rect 50484 19286 50508 19288
rect 50564 19286 50588 19288
rect 50348 19266 50644 19286
rect 50348 18010 50644 18030
rect 50404 18008 50428 18010
rect 50484 18008 50508 18010
rect 50564 18008 50588 18010
rect 50426 17956 50428 18008
rect 50490 17956 50502 18008
rect 50564 17956 50566 18008
rect 50404 17954 50428 17956
rect 50484 17954 50508 17956
rect 50564 17954 50588 17956
rect 50348 17934 50644 17954
rect 50348 16678 50644 16698
rect 50404 16676 50428 16678
rect 50484 16676 50508 16678
rect 50564 16676 50588 16678
rect 50426 16624 50428 16676
rect 50490 16624 50502 16676
rect 50564 16624 50566 16676
rect 50404 16622 50428 16624
rect 50484 16622 50508 16624
rect 50564 16622 50588 16624
rect 50348 16602 50644 16622
rect 50348 15346 50644 15366
rect 50404 15344 50428 15346
rect 50484 15344 50508 15346
rect 50564 15344 50588 15346
rect 50426 15292 50428 15344
rect 50490 15292 50502 15344
rect 50564 15292 50566 15344
rect 50404 15290 50428 15292
rect 50484 15290 50508 15292
rect 50564 15290 50588 15292
rect 50348 15270 50644 15290
rect 50348 14014 50644 14034
rect 50404 14012 50428 14014
rect 50484 14012 50508 14014
rect 50564 14012 50588 14014
rect 50426 13960 50428 14012
rect 50490 13960 50502 14012
rect 50564 13960 50566 14012
rect 50404 13958 50428 13960
rect 50484 13958 50508 13960
rect 50564 13958 50588 13960
rect 50348 13938 50644 13958
rect 50348 12682 50644 12702
rect 50404 12680 50428 12682
rect 50484 12680 50508 12682
rect 50564 12680 50588 12682
rect 50426 12628 50428 12680
rect 50490 12628 50502 12680
rect 50564 12628 50566 12680
rect 50404 12626 50428 12628
rect 50484 12626 50508 12628
rect 50564 12626 50588 12628
rect 50348 12606 50644 12626
rect 50348 11350 50644 11370
rect 50404 11348 50428 11350
rect 50484 11348 50508 11350
rect 50564 11348 50588 11350
rect 50426 11296 50428 11348
rect 50490 11296 50502 11348
rect 50564 11296 50566 11348
rect 50404 11294 50428 11296
rect 50484 11294 50508 11296
rect 50564 11294 50588 11296
rect 50348 11274 50644 11294
rect 50348 10018 50644 10038
rect 50404 10016 50428 10018
rect 50484 10016 50508 10018
rect 50564 10016 50588 10018
rect 50426 9964 50428 10016
rect 50490 9964 50502 10016
rect 50564 9964 50566 10016
rect 50404 9962 50428 9964
rect 50484 9962 50508 9964
rect 50564 9962 50588 9964
rect 50348 9942 50644 9962
rect 50230 9535 50282 9541
rect 50230 9477 50282 9483
rect 50348 8686 50644 8706
rect 50404 8684 50428 8686
rect 50484 8684 50508 8686
rect 50564 8684 50588 8686
rect 50426 8632 50428 8684
rect 50490 8632 50502 8684
rect 50564 8632 50566 8684
rect 50404 8630 50428 8632
rect 50484 8630 50508 8632
rect 50564 8630 50588 8632
rect 50348 8610 50644 8630
rect 50722 8505 50750 24869
rect 50818 19087 50846 56689
rect 51202 56161 51230 59200
rect 51286 56229 51338 56235
rect 51286 56171 51338 56177
rect 51190 56155 51242 56161
rect 51190 56097 51242 56103
rect 51094 22855 51146 22861
rect 51094 22797 51146 22803
rect 50806 19081 50858 19087
rect 50806 19023 50858 19029
rect 51106 12427 51134 22797
rect 51094 12421 51146 12427
rect 51094 12363 51146 12369
rect 50806 11829 50858 11835
rect 50806 11771 50858 11777
rect 50710 8499 50762 8505
rect 50710 8441 50762 8447
rect 50348 7354 50644 7374
rect 50404 7352 50428 7354
rect 50484 7352 50508 7354
rect 50564 7352 50588 7354
rect 50426 7300 50428 7352
rect 50490 7300 50502 7352
rect 50564 7300 50566 7352
rect 50404 7298 50428 7300
rect 50484 7298 50508 7300
rect 50564 7298 50588 7300
rect 50348 7278 50644 7298
rect 50134 7093 50186 7099
rect 50134 7035 50186 7041
rect 50134 6945 50186 6951
rect 50134 6887 50186 6893
rect 49558 6353 49610 6359
rect 49558 6295 49610 6301
rect 49570 800 49598 6295
rect 49750 6131 49802 6137
rect 49750 6073 49802 6079
rect 49654 5687 49706 5693
rect 49654 5629 49706 5635
rect 49666 3251 49694 5629
rect 49654 3245 49706 3251
rect 49654 3187 49706 3193
rect 49654 3023 49706 3029
rect 49654 2965 49706 2971
rect 49666 800 49694 2965
rect 49762 2752 49790 6073
rect 49846 4355 49898 4361
rect 49846 4297 49898 4303
rect 49858 2955 49886 4297
rect 49942 4281 49994 4287
rect 49942 4223 49994 4229
rect 49846 2949 49898 2955
rect 49846 2891 49898 2897
rect 49762 2724 49886 2752
rect 49858 800 49886 2724
rect 49954 800 49982 4223
rect 50038 2875 50090 2881
rect 50038 2817 50090 2823
rect 50050 800 50078 2817
rect 50146 800 50174 6887
rect 50818 6433 50846 11771
rect 50998 9461 51050 9467
rect 50998 9403 51050 9409
rect 51010 7765 51038 9403
rect 51190 8203 51242 8209
rect 51190 8145 51242 8151
rect 51202 7913 51230 8145
rect 51190 7907 51242 7913
rect 51190 7849 51242 7855
rect 50998 7759 51050 7765
rect 50998 7701 51050 7707
rect 50806 6427 50858 6433
rect 50806 6369 50858 6375
rect 51094 6131 51146 6137
rect 51094 6073 51146 6079
rect 50348 6022 50644 6042
rect 50404 6020 50428 6022
rect 50484 6020 50508 6022
rect 50564 6020 50588 6022
rect 50426 5968 50428 6020
rect 50490 5968 50502 6020
rect 50564 5968 50566 6020
rect 50404 5966 50428 5968
rect 50484 5966 50508 5968
rect 50564 5966 50588 5968
rect 50348 5946 50644 5966
rect 50710 5687 50762 5693
rect 50710 5629 50762 5635
rect 50422 5021 50474 5027
rect 50422 4963 50474 4969
rect 50434 4824 50462 4963
rect 50242 4796 50462 4824
rect 50242 2604 50270 4796
rect 50348 4690 50644 4710
rect 50404 4688 50428 4690
rect 50484 4688 50508 4690
rect 50564 4688 50588 4690
rect 50426 4636 50428 4688
rect 50490 4636 50502 4688
rect 50564 4636 50566 4688
rect 50404 4634 50428 4636
rect 50484 4634 50508 4636
rect 50564 4634 50588 4636
rect 50348 4614 50644 4634
rect 50722 3843 50750 5629
rect 50902 5021 50954 5027
rect 50902 4963 50954 4969
rect 50710 3837 50762 3843
rect 50710 3779 50762 3785
rect 50710 3689 50762 3695
rect 50710 3631 50762 3637
rect 50806 3689 50858 3695
rect 50806 3631 50858 3637
rect 50348 3358 50644 3378
rect 50404 3356 50428 3358
rect 50484 3356 50508 3358
rect 50564 3356 50588 3358
rect 50426 3304 50428 3356
rect 50490 3304 50502 3356
rect 50564 3304 50566 3356
rect 50404 3302 50428 3304
rect 50484 3302 50508 3304
rect 50564 3302 50588 3304
rect 50348 3282 50644 3302
rect 50242 2576 50366 2604
rect 50338 800 50366 2576
rect 50722 1864 50750 3631
rect 50434 1836 50750 1864
rect 50434 800 50462 1836
rect 50710 1765 50762 1771
rect 50710 1707 50762 1713
rect 50518 1691 50570 1697
rect 50518 1633 50570 1639
rect 50530 800 50558 1633
rect 50722 800 50750 1707
rect 50818 800 50846 3631
rect 50914 1771 50942 4963
rect 50998 4281 51050 4287
rect 50998 4223 51050 4229
rect 50902 1765 50954 1771
rect 50902 1707 50954 1713
rect 50902 1617 50954 1623
rect 50902 1559 50954 1565
rect 50914 800 50942 1559
rect 51010 800 51038 4223
rect 51106 1697 51134 6073
rect 51298 3843 51326 56171
rect 51778 55717 51806 59200
rect 52258 56975 52286 59200
rect 52246 56969 52298 56975
rect 52246 56911 52298 56917
rect 52834 56531 52862 59200
rect 53314 56531 53342 59200
rect 53890 56901 53918 59200
rect 53878 56895 53930 56901
rect 53878 56837 53930 56843
rect 53878 56747 53930 56753
rect 53878 56689 53930 56695
rect 52822 56525 52874 56531
rect 52822 56467 52874 56473
rect 53302 56525 53354 56531
rect 53302 56467 53354 56473
rect 52918 56229 52970 56235
rect 52918 56171 52970 56177
rect 51766 55711 51818 55717
rect 51766 55653 51818 55659
rect 51958 55563 52010 55569
rect 51958 55505 52010 55511
rect 51478 33881 51530 33887
rect 51478 33823 51530 33829
rect 51490 7913 51518 33823
rect 51970 32185 51998 55505
rect 52246 43575 52298 43581
rect 52246 43517 52298 43523
rect 51958 32179 52010 32185
rect 51958 32121 52010 32127
rect 51862 30773 51914 30779
rect 51862 30715 51914 30721
rect 51574 30329 51626 30335
rect 51574 30271 51626 30277
rect 51478 7907 51530 7913
rect 51478 7849 51530 7855
rect 51382 6945 51434 6951
rect 51382 6887 51434 6893
rect 51286 3837 51338 3843
rect 51286 3779 51338 3785
rect 51286 3689 51338 3695
rect 51202 3649 51286 3677
rect 51094 1691 51146 1697
rect 51094 1633 51146 1639
rect 51202 800 51230 3649
rect 51286 3631 51338 3637
rect 51394 3492 51422 6887
rect 51586 6433 51614 30271
rect 51874 13833 51902 30715
rect 52150 30403 52202 30409
rect 52150 30345 52202 30351
rect 51862 13827 51914 13833
rect 51862 13769 51914 13775
rect 51862 10793 51914 10799
rect 51862 10735 51914 10741
rect 51670 7833 51722 7839
rect 51874 7784 51902 10735
rect 51722 7781 51902 7784
rect 51670 7775 51902 7781
rect 51682 7756 51902 7775
rect 51670 7463 51722 7469
rect 51670 7405 51722 7411
rect 51574 6427 51626 6433
rect 51574 6369 51626 6375
rect 51574 6205 51626 6211
rect 51574 6147 51626 6153
rect 51298 3464 51422 3492
rect 51298 800 51326 3464
rect 51478 3023 51530 3029
rect 51478 2965 51530 2971
rect 51382 2949 51434 2955
rect 51382 2891 51434 2897
rect 51394 800 51422 2891
rect 51490 800 51518 2965
rect 51586 1623 51614 6147
rect 51574 1617 51626 1623
rect 51574 1559 51626 1565
rect 51682 800 51710 7405
rect 52162 7099 52190 30345
rect 52258 7173 52286 43517
rect 52930 37217 52958 56171
rect 52918 37211 52970 37217
rect 52918 37153 52970 37159
rect 53206 34769 53258 34775
rect 53206 34711 53258 34717
rect 52534 27591 52586 27597
rect 52534 27533 52586 27539
rect 52546 8431 52574 27533
rect 53218 23749 53246 34711
rect 53398 34177 53450 34183
rect 53398 34119 53450 34125
rect 53302 32105 53354 32111
rect 53302 32047 53354 32053
rect 53206 23743 53258 23749
rect 53206 23685 53258 23691
rect 52822 12421 52874 12427
rect 52822 12363 52874 12369
rect 52630 11681 52682 11687
rect 52630 11623 52682 11629
rect 52534 8425 52586 8431
rect 52534 8367 52586 8373
rect 52534 8129 52586 8135
rect 52534 8071 52586 8077
rect 52546 7691 52574 8071
rect 52642 7765 52670 11623
rect 52630 7759 52682 7765
rect 52630 7701 52682 7707
rect 52534 7685 52586 7691
rect 52534 7627 52586 7633
rect 52342 7463 52394 7469
rect 52342 7405 52394 7411
rect 52726 7463 52778 7469
rect 52726 7405 52778 7411
rect 52246 7167 52298 7173
rect 52246 7109 52298 7115
rect 52150 7093 52202 7099
rect 52150 7035 52202 7041
rect 52150 5687 52202 5693
rect 52150 5629 52202 5635
rect 51862 5021 51914 5027
rect 51862 4963 51914 4969
rect 51766 3097 51818 3103
rect 51766 3039 51818 3045
rect 51778 800 51806 3039
rect 51874 2955 51902 4963
rect 52054 3689 52106 3695
rect 51970 3649 52054 3677
rect 51862 2949 51914 2955
rect 51862 2891 51914 2897
rect 51970 1864 51998 3649
rect 52054 3631 52106 3637
rect 52054 3245 52106 3251
rect 52054 3187 52106 3193
rect 51874 1836 51998 1864
rect 51874 800 51902 1836
rect 52066 800 52094 3187
rect 52162 800 52190 5629
rect 52246 5021 52298 5027
rect 52246 4963 52298 4969
rect 52258 3103 52286 4963
rect 52246 3097 52298 3103
rect 52246 3039 52298 3045
rect 52246 2949 52298 2955
rect 52246 2891 52298 2897
rect 52258 800 52286 2891
rect 52354 800 52382 7405
rect 52438 6945 52490 6951
rect 52438 6887 52490 6893
rect 52450 3251 52478 6887
rect 52534 5687 52586 5693
rect 52534 5629 52586 5635
rect 52438 3245 52490 3251
rect 52438 3187 52490 3193
rect 52546 800 52574 5629
rect 52630 4355 52682 4361
rect 52630 4297 52682 4303
rect 52642 800 52670 4297
rect 52738 800 52766 7405
rect 52834 7099 52862 12363
rect 53206 8943 53258 8949
rect 53206 8885 53258 8891
rect 52918 8351 52970 8357
rect 52918 8293 52970 8299
rect 52822 7093 52874 7099
rect 52822 7035 52874 7041
rect 52930 3048 52958 8293
rect 53110 8277 53162 8283
rect 53110 8219 53162 8225
rect 53014 4281 53066 4287
rect 53014 4223 53066 4229
rect 52834 3020 52958 3048
rect 52834 2881 52862 3020
rect 52918 2949 52970 2955
rect 52918 2891 52970 2897
rect 52822 2875 52874 2881
rect 52822 2817 52874 2823
rect 52930 800 52958 2891
rect 53026 800 53054 4223
rect 53122 800 53150 8219
rect 53218 3103 53246 8885
rect 53314 8431 53342 32047
rect 53302 8425 53354 8431
rect 53302 8367 53354 8373
rect 53410 7765 53438 34119
rect 53890 21455 53918 56689
rect 54370 56531 54398 59200
rect 54946 56531 54974 59200
rect 55426 56901 55454 59200
rect 55414 56895 55466 56901
rect 55414 56837 55466 56843
rect 55510 56747 55562 56753
rect 55510 56689 55562 56695
rect 54358 56525 54410 56531
rect 54358 56467 54410 56473
rect 54934 56525 54986 56531
rect 54934 56467 54986 56473
rect 53974 56229 54026 56235
rect 53974 56171 54026 56177
rect 54550 56229 54602 56235
rect 54550 56171 54602 56177
rect 54934 56229 54986 56235
rect 54934 56171 54986 56177
rect 53878 21449 53930 21455
rect 53878 21391 53930 21397
rect 53986 19901 54014 56171
rect 54562 51425 54590 56171
rect 54550 51419 54602 51425
rect 54550 51361 54602 51367
rect 54946 50463 54974 56171
rect 55030 50753 55082 50759
rect 55030 50695 55082 50701
rect 54934 50457 54986 50463
rect 54934 50399 54986 50405
rect 54070 43649 54122 43655
rect 54070 43591 54122 43597
rect 53974 19895 54026 19901
rect 53974 19837 54026 19843
rect 54082 9911 54110 43591
rect 54646 18785 54698 18791
rect 54646 18727 54698 18733
rect 54454 14789 54506 14795
rect 54454 14731 54506 14737
rect 54070 9905 54122 9911
rect 54070 9847 54122 9853
rect 54466 9763 54494 14731
rect 54658 11095 54686 18727
rect 54646 11089 54698 11095
rect 54646 11031 54698 11037
rect 55042 10429 55070 50695
rect 55318 30773 55370 30779
rect 55318 30715 55370 30721
rect 55330 30557 55358 30715
rect 55318 30551 55370 30557
rect 55318 30493 55370 30499
rect 55522 21529 55550 56689
rect 56002 56531 56030 59200
rect 55990 56525 56042 56531
rect 55990 56467 56042 56473
rect 56482 55717 56510 59200
rect 56758 56747 56810 56753
rect 56758 56689 56810 56695
rect 56770 56457 56798 56689
rect 56758 56451 56810 56457
rect 56758 56393 56810 56399
rect 57058 56309 57086 59200
rect 57046 56303 57098 56309
rect 57046 56245 57098 56251
rect 57538 55717 57566 59200
rect 56470 55711 56522 55717
rect 56470 55653 56522 55659
rect 57526 55711 57578 55717
rect 57526 55653 57578 55659
rect 55606 55415 55658 55421
rect 55606 55357 55658 55363
rect 56278 55415 56330 55421
rect 56278 55357 56330 55363
rect 57334 55415 57386 55421
rect 57334 55357 57386 55363
rect 55618 55125 55646 55357
rect 55606 55119 55658 55125
rect 55606 55061 55658 55067
rect 56290 33517 56318 55357
rect 56854 50753 56906 50759
rect 56854 50695 56906 50701
rect 56662 35435 56714 35441
rect 56662 35377 56714 35383
rect 56278 33511 56330 33517
rect 56278 33453 56330 33459
rect 56674 26857 56702 35377
rect 56662 26851 56714 26857
rect 56662 26793 56714 26799
rect 55510 21523 55562 21529
rect 55510 21465 55562 21471
rect 56866 17294 56894 50695
rect 57142 46535 57194 46541
rect 57142 46477 57194 46483
rect 57154 37454 57182 46477
rect 57238 40097 57290 40103
rect 57238 40039 57290 40045
rect 57250 39881 57278 40039
rect 57238 39875 57290 39881
rect 57238 39817 57290 39823
rect 57154 37426 57278 37454
rect 57046 34769 57098 34775
rect 57046 34711 57098 34717
rect 56950 25445 57002 25451
rect 56950 25387 57002 25393
rect 56674 17266 56894 17294
rect 56278 11459 56330 11465
rect 56278 11401 56330 11407
rect 55030 10423 55082 10429
rect 55030 10365 55082 10371
rect 55702 10127 55754 10133
rect 55702 10069 55754 10075
rect 56086 10127 56138 10133
rect 56086 10069 56138 10075
rect 54454 9757 54506 9763
rect 54454 9699 54506 9705
rect 54262 9609 54314 9615
rect 54262 9551 54314 9557
rect 55318 9609 55370 9615
rect 55318 9551 55370 9557
rect 53782 9461 53834 9467
rect 53782 9403 53834 9409
rect 53794 9245 53822 9403
rect 53782 9239 53834 9245
rect 53782 9181 53834 9187
rect 53878 8795 53930 8801
rect 53878 8737 53930 8743
rect 53494 8277 53546 8283
rect 53494 8219 53546 8225
rect 53398 7759 53450 7765
rect 53398 7701 53450 7707
rect 53302 5021 53354 5027
rect 53302 4963 53354 4969
rect 53206 3097 53258 3103
rect 53206 3039 53258 3045
rect 53314 2900 53342 4963
rect 53398 3689 53450 3695
rect 53398 3631 53450 3637
rect 53218 2872 53342 2900
rect 53218 800 53246 2872
rect 53410 800 53438 3631
rect 53506 800 53534 8219
rect 53686 5687 53738 5693
rect 53686 5629 53738 5635
rect 53590 5613 53642 5619
rect 53590 5555 53642 5561
rect 53602 800 53630 5555
rect 53698 2955 53726 5629
rect 53782 3023 53834 3029
rect 53782 2965 53834 2971
rect 53686 2949 53738 2955
rect 53686 2891 53738 2897
rect 53794 1568 53822 2965
rect 53698 1540 53822 1568
rect 53698 800 53726 1540
rect 53890 800 53918 8737
rect 53974 6353 54026 6359
rect 53974 6295 54026 6301
rect 53986 800 54014 6295
rect 54070 4355 54122 4361
rect 54070 4297 54122 4303
rect 54082 800 54110 4297
rect 54274 800 54302 9551
rect 54934 9535 54986 9541
rect 54934 9477 54986 9483
rect 54646 8795 54698 8801
rect 54646 8737 54698 8743
rect 54658 7214 54686 8737
rect 54562 7186 54686 7214
rect 54358 3837 54410 3843
rect 54358 3779 54410 3785
rect 54370 800 54398 3779
rect 54454 3541 54506 3547
rect 54454 3483 54506 3489
rect 54466 800 54494 3483
rect 54562 800 54590 7186
rect 54742 7019 54794 7025
rect 54742 6961 54794 6967
rect 54754 800 54782 6961
rect 54838 2949 54890 2955
rect 54838 2891 54890 2897
rect 54850 800 54878 2891
rect 54946 800 54974 9477
rect 55222 6353 55274 6359
rect 55222 6295 55274 6301
rect 55126 6279 55178 6285
rect 55126 6221 55178 6227
rect 55030 6205 55082 6211
rect 55030 6147 55082 6153
rect 55042 800 55070 6147
rect 55138 4287 55166 6221
rect 55126 4281 55178 4287
rect 55126 4223 55178 4229
rect 55234 3843 55262 6295
rect 55222 3837 55274 3843
rect 55222 3779 55274 3785
rect 55222 3467 55274 3473
rect 55222 3409 55274 3415
rect 55234 800 55262 3409
rect 55330 800 55358 9551
rect 55414 7019 55466 7025
rect 55414 6961 55466 6967
rect 55426 800 55454 6961
rect 55606 4355 55658 4361
rect 55606 4297 55658 4303
rect 55618 800 55646 4297
rect 55714 800 55742 10069
rect 55894 9017 55946 9023
rect 55894 8959 55946 8965
rect 55798 7685 55850 7691
rect 55798 7627 55850 7633
rect 55810 800 55838 7627
rect 55906 4139 55934 8959
rect 55894 4133 55946 4139
rect 55894 4075 55946 4081
rect 55894 3763 55946 3769
rect 55894 3705 55946 3711
rect 55906 800 55934 3705
rect 56098 800 56126 10069
rect 56182 7685 56234 7691
rect 56182 7627 56234 7633
rect 56194 800 56222 7627
rect 56290 3677 56318 11401
rect 56470 10201 56522 10207
rect 56470 10143 56522 10149
rect 56374 6945 56426 6951
rect 56374 6887 56426 6893
rect 56386 4287 56414 6887
rect 56374 4281 56426 4287
rect 56374 4223 56426 4229
rect 56290 3649 56414 3677
rect 56278 3615 56330 3621
rect 56278 3557 56330 3563
rect 56290 800 56318 3557
rect 56386 3547 56414 3649
rect 56374 3541 56426 3547
rect 56374 3483 56426 3489
rect 56482 800 56510 10143
rect 56674 8209 56702 17266
rect 56962 13759 56990 25387
rect 56950 13753 57002 13759
rect 56950 13695 57002 13701
rect 57058 13685 57086 34711
rect 57046 13679 57098 13685
rect 57046 13621 57098 13627
rect 57250 12575 57278 37426
rect 57346 16201 57374 55357
rect 57814 54897 57866 54903
rect 57814 54839 57866 54845
rect 57718 53417 57770 53423
rect 57718 53359 57770 53365
rect 57622 38765 57674 38771
rect 57622 38707 57674 38713
rect 57334 16195 57386 16201
rect 57334 16137 57386 16143
rect 57238 12569 57290 12575
rect 57238 12511 57290 12517
rect 57526 12199 57578 12205
rect 57526 12141 57578 12147
rect 56758 10941 56810 10947
rect 56758 10883 56810 10889
rect 56662 8203 56714 8209
rect 56662 8145 56714 8151
rect 56662 7685 56714 7691
rect 56662 7627 56714 7633
rect 56674 7214 56702 7627
rect 56578 7186 56702 7214
rect 56578 800 56606 7186
rect 56662 4355 56714 4361
rect 56662 4297 56714 4303
rect 56674 800 56702 4297
rect 56770 800 56798 10883
rect 56854 10867 56906 10873
rect 56854 10809 56906 10815
rect 56866 3251 56894 10809
rect 57238 9017 57290 9023
rect 57238 8959 57290 8965
rect 56950 8351 57002 8357
rect 56950 8293 57002 8299
rect 56854 3245 56906 3251
rect 56854 3187 56906 3193
rect 56962 800 56990 8293
rect 57142 7611 57194 7617
rect 57142 7553 57194 7559
rect 57046 6501 57098 6507
rect 57046 6443 57098 6449
rect 57058 5120 57086 6443
rect 57154 5249 57182 7553
rect 57142 5243 57194 5249
rect 57142 5185 57194 5191
rect 57058 5092 57182 5120
rect 57046 5021 57098 5027
rect 57046 4963 57098 4969
rect 57058 800 57086 4963
rect 57154 3843 57182 5092
rect 57142 3837 57194 3843
rect 57142 3779 57194 3785
rect 57142 3541 57194 3547
rect 57142 3483 57194 3489
rect 57154 800 57182 3483
rect 57250 800 57278 8959
rect 57334 8943 57386 8949
rect 57334 8885 57386 8891
rect 57346 3917 57374 8885
rect 57430 5687 57482 5693
rect 57430 5629 57482 5635
rect 57334 3911 57386 3917
rect 57334 3853 57386 3859
rect 57334 3763 57386 3769
rect 57334 3705 57386 3711
rect 57346 3177 57374 3705
rect 57334 3171 57386 3177
rect 57334 3113 57386 3119
rect 57442 800 57470 5629
rect 57538 800 57566 12141
rect 57634 9856 57662 38707
rect 57730 13463 57758 53359
rect 57718 13457 57770 13463
rect 57718 13399 57770 13405
rect 57634 9828 57758 9856
rect 57826 9837 57854 54839
rect 58114 54385 58142 59200
rect 58594 56901 58622 59200
rect 58582 56895 58634 56901
rect 58582 56837 58634 56843
rect 59170 55199 59198 59200
rect 59158 55193 59210 55199
rect 59158 55135 59210 55141
rect 58102 54379 58154 54385
rect 58102 54321 58154 54327
rect 58102 54083 58154 54089
rect 58102 54025 58154 54031
rect 57910 39431 57962 39437
rect 57910 39373 57962 39379
rect 57922 11095 57950 39373
rect 58114 21603 58142 54025
rect 59650 53867 59678 59200
rect 59638 53861 59690 53867
rect 59638 53803 59690 53809
rect 58102 21597 58154 21603
rect 58102 21539 58154 21545
rect 59734 11607 59786 11613
rect 59734 11549 59786 11555
rect 57910 11089 57962 11095
rect 57910 11031 57962 11037
rect 58582 10571 58634 10577
rect 58582 10513 58634 10519
rect 57622 9683 57674 9689
rect 57622 9625 57674 9631
rect 57634 800 57662 9625
rect 57730 8135 57758 9828
rect 57814 9831 57866 9837
rect 57814 9773 57866 9779
rect 58390 8277 58442 8283
rect 58390 8219 58442 8225
rect 57718 8129 57770 8135
rect 57718 8071 57770 8077
rect 58102 6353 58154 6359
rect 58102 6295 58154 6301
rect 57814 4947 57866 4953
rect 57814 4889 57866 4895
rect 57826 800 57854 4889
rect 57910 4133 57962 4139
rect 57910 4075 57962 4081
rect 57922 800 57950 4075
rect 58006 3171 58058 3177
rect 58006 3113 58058 3119
rect 58018 800 58046 3113
rect 58114 800 58142 6295
rect 58294 3245 58346 3251
rect 58294 3187 58346 3193
rect 58306 800 58334 3187
rect 58402 800 58430 8219
rect 58486 7019 58538 7025
rect 58486 6961 58538 6967
rect 58498 800 58526 6961
rect 58594 800 58622 10513
rect 58966 8573 59018 8579
rect 58966 8515 59018 8521
rect 58774 7759 58826 7765
rect 58774 7701 58826 7707
rect 58786 800 58814 7701
rect 58870 6279 58922 6285
rect 58870 6221 58922 6227
rect 58882 800 58910 6221
rect 58978 800 59006 8515
rect 59350 7537 59402 7543
rect 59350 7479 59402 7485
rect 59254 4873 59306 4879
rect 59254 4815 59306 4821
rect 59158 3911 59210 3917
rect 59158 3853 59210 3859
rect 59170 800 59198 3853
rect 59266 800 59294 4815
rect 59362 800 59390 7479
rect 59638 5613 59690 5619
rect 59638 5555 59690 5561
rect 59446 4281 59498 4287
rect 59446 4223 59498 4229
rect 59458 800 59486 4223
rect 59650 800 59678 5555
rect 59746 800 59774 11549
rect 59830 8425 59882 8431
rect 59830 8367 59882 8373
rect 59842 800 59870 8367
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1364 0 1420 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2708 0 2764 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3188 0 3244 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 4052 0 4108 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4532 0 4588 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4916 0 4972 800
rect 5012 0 5068 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5396 0 5452 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5876 0 5932 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6260 0 6316 800
rect 6356 0 6412 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6740 0 6796 800
rect 6836 0 6892 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7220 0 7276 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7604 0 7660 800
rect 7700 0 7756 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 8084 0 8140 800
rect 8180 0 8236 800
rect 8276 0 8332 800
rect 8468 0 8524 800
rect 8564 0 8620 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8948 0 9004 800
rect 9044 0 9100 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9428 0 9484 800
rect 9524 0 9580 800
rect 9620 0 9676 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10004 0 10060 800
rect 10100 0 10156 800
rect 10292 0 10348 800
rect 10388 0 10444 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10772 0 10828 800
rect 10868 0 10924 800
rect 10964 0 11020 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11348 0 11404 800
rect 11444 0 11500 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11828 0 11884 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12212 0 12268 800
rect 12308 0 12364 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12692 0 12748 800
rect 12788 0 12844 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13172 0 13228 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13652 0 13708 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14036 0 14092 800
rect 14132 0 14188 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14516 0 14572 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 14996 0 15052 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15380 0 15436 800
rect 15476 0 15532 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15860 0 15916 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16340 0 16396 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17204 0 17260 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17684 0 17740 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19028 0 19084 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20468 0 20524 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21812 0 21868 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22292 0 22348 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23156 0 23212 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23636 0 23692 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 24020 0 24076 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24500 0 24556 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24980 0 25036 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25364 0 25420 800
rect 25460 0 25516 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25844 0 25900 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26324 0 26380 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26708 0 26764 800
rect 26804 0 26860 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27188 0 27244 800
rect 27284 0 27340 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27668 0 27724 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 28052 0 28108 800
rect 28148 0 28204 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28532 0 28588 800
rect 28628 0 28684 800
rect 28724 0 28780 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29108 0 29164 800
rect 29204 0 29260 800
rect 29396 0 29452 800
rect 29492 0 29548 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29876 0 29932 800
rect 29972 0 30028 800
rect 30068 0 30124 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30452 0 30508 800
rect 30548 0 30604 800
rect 30740 0 30796 800
rect 30836 0 30892 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31220 0 31276 800
rect 31316 0 31372 800
rect 31412 0 31468 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31796 0 31852 800
rect 31892 0 31948 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32276 0 32332 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32660 0 32716 800
rect 32756 0 32812 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33140 0 33196 800
rect 33236 0 33292 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33620 0 33676 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34100 0 34156 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34484 0 34540 800
rect 34580 0 34636 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 34964 0 35020 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35444 0 35500 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36308 0 36364 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36788 0 36844 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37652 0 37708 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38132 0 38188 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39476 0 39532 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40916 0 40972 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42260 0 42316 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42740 0 42796 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43604 0 43660 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 44084 0 44140 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44468 0 44524 800
rect 44564 0 44620 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44948 0 45004 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45428 0 45484 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45812 0 45868 800
rect 45908 0 45964 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46292 0 46348 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46772 0 46828 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47156 0 47212 800
rect 47252 0 47308 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47636 0 47692 800
rect 47732 0 47788 800
rect 47828 0 47884 800
rect 48020 0 48076 800
rect 48116 0 48172 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48500 0 48556 800
rect 48596 0 48652 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48980 0 49036 800
rect 49076 0 49132 800
rect 49172 0 49228 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49556 0 49612 800
rect 49652 0 49708 800
rect 49844 0 49900 800
rect 49940 0 49996 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50324 0 50380 800
rect 50420 0 50476 800
rect 50516 0 50572 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50900 0 50956 800
rect 50996 0 51052 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51380 0 51436 800
rect 51476 0 51532 800
rect 51668 0 51724 800
rect 51764 0 51820 800
rect 51860 0 51916 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52244 0 52300 800
rect 52340 0 52396 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52724 0 52780 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53108 0 53164 800
rect 53204 0 53260 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53588 0 53644 800
rect 53684 0 53740 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54068 0 54124 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54548 0 54604 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 54932 0 54988 800
rect 55028 0 55084 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55412 0 55468 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55892 0 55948 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56756 0 56812 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57236 0 57292 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58580 0 58636 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< via2 >>
rect 4268 57302 4324 57304
rect 4348 57302 4404 57304
rect 4428 57302 4484 57304
rect 4508 57302 4564 57304
rect 4268 57250 4294 57302
rect 4294 57250 4324 57302
rect 4348 57250 4358 57302
rect 4358 57250 4404 57302
rect 4428 57250 4474 57302
rect 4474 57250 4484 57302
rect 4508 57250 4538 57302
rect 4538 57250 4564 57302
rect 4268 57248 4324 57250
rect 4348 57248 4404 57250
rect 4428 57248 4484 57250
rect 4508 57248 4564 57250
rect 4268 55970 4324 55972
rect 4348 55970 4404 55972
rect 4428 55970 4484 55972
rect 4508 55970 4564 55972
rect 4268 55918 4294 55970
rect 4294 55918 4324 55970
rect 4348 55918 4358 55970
rect 4358 55918 4404 55970
rect 4428 55918 4474 55970
rect 4474 55918 4484 55970
rect 4508 55918 4538 55970
rect 4538 55918 4564 55970
rect 4268 55916 4324 55918
rect 4348 55916 4404 55918
rect 4428 55916 4484 55918
rect 4508 55916 4564 55918
rect 4268 54638 4324 54640
rect 4348 54638 4404 54640
rect 4428 54638 4484 54640
rect 4508 54638 4564 54640
rect 4268 54586 4294 54638
rect 4294 54586 4324 54638
rect 4348 54586 4358 54638
rect 4358 54586 4404 54638
rect 4428 54586 4474 54638
rect 4474 54586 4484 54638
rect 4508 54586 4538 54638
rect 4538 54586 4564 54638
rect 4268 54584 4324 54586
rect 4348 54584 4404 54586
rect 4428 54584 4484 54586
rect 4508 54584 4564 54586
rect 4268 53306 4324 53308
rect 4348 53306 4404 53308
rect 4428 53306 4484 53308
rect 4508 53306 4564 53308
rect 4268 53254 4294 53306
rect 4294 53254 4324 53306
rect 4348 53254 4358 53306
rect 4358 53254 4404 53306
rect 4428 53254 4474 53306
rect 4474 53254 4484 53306
rect 4508 53254 4538 53306
rect 4538 53254 4564 53306
rect 4268 53252 4324 53254
rect 4348 53252 4404 53254
rect 4428 53252 4484 53254
rect 4508 53252 4564 53254
rect 4268 51974 4324 51976
rect 4348 51974 4404 51976
rect 4428 51974 4484 51976
rect 4508 51974 4564 51976
rect 4268 51922 4294 51974
rect 4294 51922 4324 51974
rect 4348 51922 4358 51974
rect 4358 51922 4404 51974
rect 4428 51922 4474 51974
rect 4474 51922 4484 51974
rect 4508 51922 4538 51974
rect 4538 51922 4564 51974
rect 4268 51920 4324 51922
rect 4348 51920 4404 51922
rect 4428 51920 4484 51922
rect 4508 51920 4564 51922
rect 4268 50642 4324 50644
rect 4348 50642 4404 50644
rect 4428 50642 4484 50644
rect 4508 50642 4564 50644
rect 4268 50590 4294 50642
rect 4294 50590 4324 50642
rect 4348 50590 4358 50642
rect 4358 50590 4404 50642
rect 4428 50590 4474 50642
rect 4474 50590 4484 50642
rect 4508 50590 4538 50642
rect 4538 50590 4564 50642
rect 4268 50588 4324 50590
rect 4348 50588 4404 50590
rect 4428 50588 4484 50590
rect 4508 50588 4564 50590
rect 4268 49310 4324 49312
rect 4348 49310 4404 49312
rect 4428 49310 4484 49312
rect 4508 49310 4564 49312
rect 4268 49258 4294 49310
rect 4294 49258 4324 49310
rect 4348 49258 4358 49310
rect 4358 49258 4404 49310
rect 4428 49258 4474 49310
rect 4474 49258 4484 49310
rect 4508 49258 4538 49310
rect 4538 49258 4564 49310
rect 4268 49256 4324 49258
rect 4348 49256 4404 49258
rect 4428 49256 4484 49258
rect 4508 49256 4564 49258
rect 4268 47978 4324 47980
rect 4348 47978 4404 47980
rect 4428 47978 4484 47980
rect 4508 47978 4564 47980
rect 4268 47926 4294 47978
rect 4294 47926 4324 47978
rect 4348 47926 4358 47978
rect 4358 47926 4404 47978
rect 4428 47926 4474 47978
rect 4474 47926 4484 47978
rect 4508 47926 4538 47978
rect 4538 47926 4564 47978
rect 4268 47924 4324 47926
rect 4348 47924 4404 47926
rect 4428 47924 4484 47926
rect 4508 47924 4564 47926
rect 4268 46646 4324 46648
rect 4348 46646 4404 46648
rect 4428 46646 4484 46648
rect 4508 46646 4564 46648
rect 4268 46594 4294 46646
rect 4294 46594 4324 46646
rect 4348 46594 4358 46646
rect 4358 46594 4404 46646
rect 4428 46594 4474 46646
rect 4474 46594 4484 46646
rect 4508 46594 4538 46646
rect 4538 46594 4564 46646
rect 4268 46592 4324 46594
rect 4348 46592 4404 46594
rect 4428 46592 4484 46594
rect 4508 46592 4564 46594
rect 4268 45314 4324 45316
rect 4348 45314 4404 45316
rect 4428 45314 4484 45316
rect 4508 45314 4564 45316
rect 4268 45262 4294 45314
rect 4294 45262 4324 45314
rect 4348 45262 4358 45314
rect 4358 45262 4404 45314
rect 4428 45262 4474 45314
rect 4474 45262 4484 45314
rect 4508 45262 4538 45314
rect 4538 45262 4564 45314
rect 4268 45260 4324 45262
rect 4348 45260 4404 45262
rect 4428 45260 4484 45262
rect 4508 45260 4564 45262
rect 4268 43982 4324 43984
rect 4348 43982 4404 43984
rect 4428 43982 4484 43984
rect 4508 43982 4564 43984
rect 4268 43930 4294 43982
rect 4294 43930 4324 43982
rect 4348 43930 4358 43982
rect 4358 43930 4404 43982
rect 4428 43930 4474 43982
rect 4474 43930 4484 43982
rect 4508 43930 4538 43982
rect 4538 43930 4564 43982
rect 4268 43928 4324 43930
rect 4348 43928 4404 43930
rect 4428 43928 4484 43930
rect 4508 43928 4564 43930
rect 4268 42650 4324 42652
rect 4348 42650 4404 42652
rect 4428 42650 4484 42652
rect 4508 42650 4564 42652
rect 4268 42598 4294 42650
rect 4294 42598 4324 42650
rect 4348 42598 4358 42650
rect 4358 42598 4404 42650
rect 4428 42598 4474 42650
rect 4474 42598 4484 42650
rect 4508 42598 4538 42650
rect 4538 42598 4564 42650
rect 4268 42596 4324 42598
rect 4348 42596 4404 42598
rect 4428 42596 4484 42598
rect 4508 42596 4564 42598
rect 4268 41318 4324 41320
rect 4348 41318 4404 41320
rect 4428 41318 4484 41320
rect 4508 41318 4564 41320
rect 4268 41266 4294 41318
rect 4294 41266 4324 41318
rect 4348 41266 4358 41318
rect 4358 41266 4404 41318
rect 4428 41266 4474 41318
rect 4474 41266 4484 41318
rect 4508 41266 4538 41318
rect 4538 41266 4564 41318
rect 4268 41264 4324 41266
rect 4348 41264 4404 41266
rect 4428 41264 4484 41266
rect 4508 41264 4564 41266
rect 4268 39986 4324 39988
rect 4348 39986 4404 39988
rect 4428 39986 4484 39988
rect 4508 39986 4564 39988
rect 4268 39934 4294 39986
rect 4294 39934 4324 39986
rect 4348 39934 4358 39986
rect 4358 39934 4404 39986
rect 4428 39934 4474 39986
rect 4474 39934 4484 39986
rect 4508 39934 4538 39986
rect 4538 39934 4564 39986
rect 4268 39932 4324 39934
rect 4348 39932 4404 39934
rect 4428 39932 4484 39934
rect 4508 39932 4564 39934
rect 4268 38654 4324 38656
rect 4348 38654 4404 38656
rect 4428 38654 4484 38656
rect 4508 38654 4564 38656
rect 4268 38602 4294 38654
rect 4294 38602 4324 38654
rect 4348 38602 4358 38654
rect 4358 38602 4404 38654
rect 4428 38602 4474 38654
rect 4474 38602 4484 38654
rect 4508 38602 4538 38654
rect 4538 38602 4564 38654
rect 4268 38600 4324 38602
rect 4348 38600 4404 38602
rect 4428 38600 4484 38602
rect 4508 38600 4564 38602
rect 4268 37322 4324 37324
rect 4348 37322 4404 37324
rect 4428 37322 4484 37324
rect 4508 37322 4564 37324
rect 4268 37270 4294 37322
rect 4294 37270 4324 37322
rect 4348 37270 4358 37322
rect 4358 37270 4404 37322
rect 4428 37270 4474 37322
rect 4474 37270 4484 37322
rect 4508 37270 4538 37322
rect 4538 37270 4564 37322
rect 4268 37268 4324 37270
rect 4348 37268 4404 37270
rect 4428 37268 4484 37270
rect 4508 37268 4564 37270
rect 4268 35990 4324 35992
rect 4348 35990 4404 35992
rect 4428 35990 4484 35992
rect 4508 35990 4564 35992
rect 4268 35938 4294 35990
rect 4294 35938 4324 35990
rect 4348 35938 4358 35990
rect 4358 35938 4404 35990
rect 4428 35938 4474 35990
rect 4474 35938 4484 35990
rect 4508 35938 4538 35990
rect 4538 35938 4564 35990
rect 4268 35936 4324 35938
rect 4348 35936 4404 35938
rect 4428 35936 4484 35938
rect 4508 35936 4564 35938
rect 4268 34658 4324 34660
rect 4348 34658 4404 34660
rect 4428 34658 4484 34660
rect 4508 34658 4564 34660
rect 4268 34606 4294 34658
rect 4294 34606 4324 34658
rect 4348 34606 4358 34658
rect 4358 34606 4404 34658
rect 4428 34606 4474 34658
rect 4474 34606 4484 34658
rect 4508 34606 4538 34658
rect 4538 34606 4564 34658
rect 4268 34604 4324 34606
rect 4348 34604 4404 34606
rect 4428 34604 4484 34606
rect 4508 34604 4564 34606
rect 4268 33326 4324 33328
rect 4348 33326 4404 33328
rect 4428 33326 4484 33328
rect 4508 33326 4564 33328
rect 4268 33274 4294 33326
rect 4294 33274 4324 33326
rect 4348 33274 4358 33326
rect 4358 33274 4404 33326
rect 4428 33274 4474 33326
rect 4474 33274 4484 33326
rect 4508 33274 4538 33326
rect 4538 33274 4564 33326
rect 4268 33272 4324 33274
rect 4348 33272 4404 33274
rect 4428 33272 4484 33274
rect 4508 33272 4564 33274
rect 4268 31994 4324 31996
rect 4348 31994 4404 31996
rect 4428 31994 4484 31996
rect 4508 31994 4564 31996
rect 4268 31942 4294 31994
rect 4294 31942 4324 31994
rect 4348 31942 4358 31994
rect 4358 31942 4404 31994
rect 4428 31942 4474 31994
rect 4474 31942 4484 31994
rect 4508 31942 4538 31994
rect 4538 31942 4564 31994
rect 4268 31940 4324 31942
rect 4348 31940 4404 31942
rect 4428 31940 4484 31942
rect 4508 31940 4564 31942
rect 4268 30662 4324 30664
rect 4348 30662 4404 30664
rect 4428 30662 4484 30664
rect 4508 30662 4564 30664
rect 4268 30610 4294 30662
rect 4294 30610 4324 30662
rect 4348 30610 4358 30662
rect 4358 30610 4404 30662
rect 4428 30610 4474 30662
rect 4474 30610 4484 30662
rect 4508 30610 4538 30662
rect 4538 30610 4564 30662
rect 4268 30608 4324 30610
rect 4348 30608 4404 30610
rect 4428 30608 4484 30610
rect 4508 30608 4564 30610
rect 4268 29330 4324 29332
rect 4348 29330 4404 29332
rect 4428 29330 4484 29332
rect 4508 29330 4564 29332
rect 4268 29278 4294 29330
rect 4294 29278 4324 29330
rect 4348 29278 4358 29330
rect 4358 29278 4404 29330
rect 4428 29278 4474 29330
rect 4474 29278 4484 29330
rect 4508 29278 4538 29330
rect 4538 29278 4564 29330
rect 4268 29276 4324 29278
rect 4348 29276 4404 29278
rect 4428 29276 4484 29278
rect 4508 29276 4564 29278
rect 4268 27998 4324 28000
rect 4348 27998 4404 28000
rect 4428 27998 4484 28000
rect 4508 27998 4564 28000
rect 4268 27946 4294 27998
rect 4294 27946 4324 27998
rect 4348 27946 4358 27998
rect 4358 27946 4404 27998
rect 4428 27946 4474 27998
rect 4474 27946 4484 27998
rect 4508 27946 4538 27998
rect 4538 27946 4564 27998
rect 4268 27944 4324 27946
rect 4348 27944 4404 27946
rect 4428 27944 4484 27946
rect 4508 27944 4564 27946
rect 4268 26666 4324 26668
rect 4348 26666 4404 26668
rect 4428 26666 4484 26668
rect 4508 26666 4564 26668
rect 4268 26614 4294 26666
rect 4294 26614 4324 26666
rect 4348 26614 4358 26666
rect 4358 26614 4404 26666
rect 4428 26614 4474 26666
rect 4474 26614 4484 26666
rect 4508 26614 4538 26666
rect 4538 26614 4564 26666
rect 4268 26612 4324 26614
rect 4348 26612 4404 26614
rect 4428 26612 4484 26614
rect 4508 26612 4564 26614
rect 4268 25334 4324 25336
rect 4348 25334 4404 25336
rect 4428 25334 4484 25336
rect 4508 25334 4564 25336
rect 4268 25282 4294 25334
rect 4294 25282 4324 25334
rect 4348 25282 4358 25334
rect 4358 25282 4404 25334
rect 4428 25282 4474 25334
rect 4474 25282 4484 25334
rect 4508 25282 4538 25334
rect 4538 25282 4564 25334
rect 4268 25280 4324 25282
rect 4348 25280 4404 25282
rect 4428 25280 4484 25282
rect 4508 25280 4564 25282
rect 4268 24002 4324 24004
rect 4348 24002 4404 24004
rect 4428 24002 4484 24004
rect 4508 24002 4564 24004
rect 4268 23950 4294 24002
rect 4294 23950 4324 24002
rect 4348 23950 4358 24002
rect 4358 23950 4404 24002
rect 4428 23950 4474 24002
rect 4474 23950 4484 24002
rect 4508 23950 4538 24002
rect 4538 23950 4564 24002
rect 4268 23948 4324 23950
rect 4348 23948 4404 23950
rect 4428 23948 4484 23950
rect 4508 23948 4564 23950
rect 4268 22670 4324 22672
rect 4348 22670 4404 22672
rect 4428 22670 4484 22672
rect 4508 22670 4564 22672
rect 4268 22618 4294 22670
rect 4294 22618 4324 22670
rect 4348 22618 4358 22670
rect 4358 22618 4404 22670
rect 4428 22618 4474 22670
rect 4474 22618 4484 22670
rect 4508 22618 4538 22670
rect 4538 22618 4564 22670
rect 4268 22616 4324 22618
rect 4348 22616 4404 22618
rect 4428 22616 4484 22618
rect 4508 22616 4564 22618
rect 4268 21338 4324 21340
rect 4348 21338 4404 21340
rect 4428 21338 4484 21340
rect 4508 21338 4564 21340
rect 4268 21286 4294 21338
rect 4294 21286 4324 21338
rect 4348 21286 4358 21338
rect 4358 21286 4404 21338
rect 4428 21286 4474 21338
rect 4474 21286 4484 21338
rect 4508 21286 4538 21338
rect 4538 21286 4564 21338
rect 4268 21284 4324 21286
rect 4348 21284 4404 21286
rect 4428 21284 4484 21286
rect 4508 21284 4564 21286
rect 4268 20006 4324 20008
rect 4348 20006 4404 20008
rect 4428 20006 4484 20008
rect 4508 20006 4564 20008
rect 4268 19954 4294 20006
rect 4294 19954 4324 20006
rect 4348 19954 4358 20006
rect 4358 19954 4404 20006
rect 4428 19954 4474 20006
rect 4474 19954 4484 20006
rect 4508 19954 4538 20006
rect 4538 19954 4564 20006
rect 4268 19952 4324 19954
rect 4348 19952 4404 19954
rect 4428 19952 4484 19954
rect 4508 19952 4564 19954
rect 4268 18674 4324 18676
rect 4348 18674 4404 18676
rect 4428 18674 4484 18676
rect 4508 18674 4564 18676
rect 4268 18622 4294 18674
rect 4294 18622 4324 18674
rect 4348 18622 4358 18674
rect 4358 18622 4404 18674
rect 4428 18622 4474 18674
rect 4474 18622 4484 18674
rect 4508 18622 4538 18674
rect 4538 18622 4564 18674
rect 4268 18620 4324 18622
rect 4348 18620 4404 18622
rect 4428 18620 4484 18622
rect 4508 18620 4564 18622
rect 4268 17342 4324 17344
rect 4348 17342 4404 17344
rect 4428 17342 4484 17344
rect 4508 17342 4564 17344
rect 4268 17290 4294 17342
rect 4294 17290 4324 17342
rect 4348 17290 4358 17342
rect 4358 17290 4404 17342
rect 4428 17290 4474 17342
rect 4474 17290 4484 17342
rect 4508 17290 4538 17342
rect 4538 17290 4564 17342
rect 4268 17288 4324 17290
rect 4348 17288 4404 17290
rect 4428 17288 4484 17290
rect 4508 17288 4564 17290
rect 4268 16010 4324 16012
rect 4348 16010 4404 16012
rect 4428 16010 4484 16012
rect 4508 16010 4564 16012
rect 4268 15958 4294 16010
rect 4294 15958 4324 16010
rect 4348 15958 4358 16010
rect 4358 15958 4404 16010
rect 4428 15958 4474 16010
rect 4474 15958 4484 16010
rect 4508 15958 4538 16010
rect 4538 15958 4564 16010
rect 4268 15956 4324 15958
rect 4348 15956 4404 15958
rect 4428 15956 4484 15958
rect 4508 15956 4564 15958
rect 4268 14678 4324 14680
rect 4348 14678 4404 14680
rect 4428 14678 4484 14680
rect 4508 14678 4564 14680
rect 4268 14626 4294 14678
rect 4294 14626 4324 14678
rect 4348 14626 4358 14678
rect 4358 14626 4404 14678
rect 4428 14626 4474 14678
rect 4474 14626 4484 14678
rect 4508 14626 4538 14678
rect 4538 14626 4564 14678
rect 4268 14624 4324 14626
rect 4348 14624 4404 14626
rect 4428 14624 4484 14626
rect 4508 14624 4564 14626
rect 4268 13346 4324 13348
rect 4348 13346 4404 13348
rect 4428 13346 4484 13348
rect 4508 13346 4564 13348
rect 4268 13294 4294 13346
rect 4294 13294 4324 13346
rect 4348 13294 4358 13346
rect 4358 13294 4404 13346
rect 4428 13294 4474 13346
rect 4474 13294 4484 13346
rect 4508 13294 4538 13346
rect 4538 13294 4564 13346
rect 4268 13292 4324 13294
rect 4348 13292 4404 13294
rect 4428 13292 4484 13294
rect 4508 13292 4564 13294
rect 4268 12014 4324 12016
rect 4348 12014 4404 12016
rect 4428 12014 4484 12016
rect 4508 12014 4564 12016
rect 4268 11962 4294 12014
rect 4294 11962 4324 12014
rect 4348 11962 4358 12014
rect 4358 11962 4404 12014
rect 4428 11962 4474 12014
rect 4474 11962 4484 12014
rect 4508 11962 4538 12014
rect 4538 11962 4564 12014
rect 4268 11960 4324 11962
rect 4348 11960 4404 11962
rect 4428 11960 4484 11962
rect 4508 11960 4564 11962
rect 4268 10682 4324 10684
rect 4348 10682 4404 10684
rect 4428 10682 4484 10684
rect 4508 10682 4564 10684
rect 4268 10630 4294 10682
rect 4294 10630 4324 10682
rect 4348 10630 4358 10682
rect 4358 10630 4404 10682
rect 4428 10630 4474 10682
rect 4474 10630 4484 10682
rect 4508 10630 4538 10682
rect 4538 10630 4564 10682
rect 4268 10628 4324 10630
rect 4348 10628 4404 10630
rect 4428 10628 4484 10630
rect 4508 10628 4564 10630
rect 4268 9350 4324 9352
rect 4348 9350 4404 9352
rect 4428 9350 4484 9352
rect 4508 9350 4564 9352
rect 4268 9298 4294 9350
rect 4294 9298 4324 9350
rect 4348 9298 4358 9350
rect 4358 9298 4404 9350
rect 4428 9298 4474 9350
rect 4474 9298 4484 9350
rect 4508 9298 4538 9350
rect 4538 9298 4564 9350
rect 4268 9296 4324 9298
rect 4348 9296 4404 9298
rect 4428 9296 4484 9298
rect 4508 9296 4564 9298
rect 4268 8018 4324 8020
rect 4348 8018 4404 8020
rect 4428 8018 4484 8020
rect 4508 8018 4564 8020
rect 4268 7966 4294 8018
rect 4294 7966 4324 8018
rect 4348 7966 4358 8018
rect 4358 7966 4404 8018
rect 4428 7966 4474 8018
rect 4474 7966 4484 8018
rect 4508 7966 4538 8018
rect 4538 7966 4564 8018
rect 4268 7964 4324 7966
rect 4348 7964 4404 7966
rect 4428 7964 4484 7966
rect 4508 7964 4564 7966
rect 4268 6686 4324 6688
rect 4348 6686 4404 6688
rect 4428 6686 4484 6688
rect 4508 6686 4564 6688
rect 4268 6634 4294 6686
rect 4294 6634 4324 6686
rect 4348 6634 4358 6686
rect 4358 6634 4404 6686
rect 4428 6634 4474 6686
rect 4474 6634 4484 6686
rect 4508 6634 4538 6686
rect 4538 6634 4564 6686
rect 4268 6632 4324 6634
rect 4348 6632 4404 6634
rect 4428 6632 4484 6634
rect 4508 6632 4564 6634
rect 4268 5354 4324 5356
rect 4348 5354 4404 5356
rect 4428 5354 4484 5356
rect 4508 5354 4564 5356
rect 4268 5302 4294 5354
rect 4294 5302 4324 5354
rect 4348 5302 4358 5354
rect 4358 5302 4404 5354
rect 4428 5302 4474 5354
rect 4474 5302 4484 5354
rect 4508 5302 4538 5354
rect 4538 5302 4564 5354
rect 4268 5300 4324 5302
rect 4348 5300 4404 5302
rect 4428 5300 4484 5302
rect 4508 5300 4564 5302
rect 4268 4022 4324 4024
rect 4348 4022 4404 4024
rect 4428 4022 4484 4024
rect 4508 4022 4564 4024
rect 4268 3970 4294 4022
rect 4294 3970 4324 4022
rect 4348 3970 4358 4022
rect 4358 3970 4404 4022
rect 4428 3970 4474 4022
rect 4474 3970 4484 4022
rect 4508 3970 4538 4022
rect 4538 3970 4564 4022
rect 4268 3968 4324 3970
rect 4348 3968 4404 3970
rect 4428 3968 4484 3970
rect 4508 3968 4564 3970
rect 4268 2690 4324 2692
rect 4348 2690 4404 2692
rect 4428 2690 4484 2692
rect 4508 2690 4564 2692
rect 4268 2638 4294 2690
rect 4294 2638 4324 2690
rect 4348 2638 4358 2690
rect 4358 2638 4404 2690
rect 4428 2638 4474 2690
rect 4474 2638 4484 2690
rect 4508 2638 4538 2690
rect 4538 2638 4564 2690
rect 4268 2636 4324 2638
rect 4348 2636 4404 2638
rect 4428 2636 4484 2638
rect 4508 2636 4564 2638
rect 4916 7759 4972 7798
rect 4916 7742 4918 7759
rect 4918 7742 4970 7759
rect 4970 7742 4972 7759
rect 7604 14419 7660 14458
rect 7604 14402 7606 14419
rect 7606 14402 7658 14419
rect 7658 14402 7660 14419
rect 7940 8778 7996 8834
rect 7940 7890 7996 7946
rect 8180 14441 8182 14458
rect 8182 14441 8234 14458
rect 8234 14441 8236 14458
rect 8180 14402 8236 14441
rect 8276 8778 8332 8834
rect 8228 7611 8284 7650
rect 8228 7594 8230 7611
rect 8230 7594 8282 7611
rect 8282 7594 8284 7611
rect 8564 7742 8620 7798
rect 9524 7594 9580 7650
rect 12212 7890 12268 7946
rect 19628 56636 19684 56638
rect 19708 56636 19764 56638
rect 19788 56636 19844 56638
rect 19868 56636 19924 56638
rect 19628 56584 19654 56636
rect 19654 56584 19684 56636
rect 19708 56584 19718 56636
rect 19718 56584 19764 56636
rect 19788 56584 19834 56636
rect 19834 56584 19844 56636
rect 19868 56584 19898 56636
rect 19898 56584 19924 56636
rect 19628 56582 19684 56584
rect 19708 56582 19764 56584
rect 19788 56582 19844 56584
rect 19868 56582 19924 56584
rect 19628 55304 19684 55306
rect 19708 55304 19764 55306
rect 19788 55304 19844 55306
rect 19868 55304 19924 55306
rect 19628 55252 19654 55304
rect 19654 55252 19684 55304
rect 19708 55252 19718 55304
rect 19718 55252 19764 55304
rect 19788 55252 19834 55304
rect 19834 55252 19844 55304
rect 19868 55252 19898 55304
rect 19898 55252 19924 55304
rect 19628 55250 19684 55252
rect 19708 55250 19764 55252
rect 19788 55250 19844 55252
rect 19868 55250 19924 55252
rect 19628 53972 19684 53974
rect 19708 53972 19764 53974
rect 19788 53972 19844 53974
rect 19868 53972 19924 53974
rect 19628 53920 19654 53972
rect 19654 53920 19684 53972
rect 19708 53920 19718 53972
rect 19718 53920 19764 53972
rect 19788 53920 19834 53972
rect 19834 53920 19844 53972
rect 19868 53920 19898 53972
rect 19898 53920 19924 53972
rect 19628 53918 19684 53920
rect 19708 53918 19764 53920
rect 19788 53918 19844 53920
rect 19868 53918 19924 53920
rect 19628 52640 19684 52642
rect 19708 52640 19764 52642
rect 19788 52640 19844 52642
rect 19868 52640 19924 52642
rect 19628 52588 19654 52640
rect 19654 52588 19684 52640
rect 19708 52588 19718 52640
rect 19718 52588 19764 52640
rect 19788 52588 19834 52640
rect 19834 52588 19844 52640
rect 19868 52588 19898 52640
rect 19898 52588 19924 52640
rect 19628 52586 19684 52588
rect 19708 52586 19764 52588
rect 19788 52586 19844 52588
rect 19868 52586 19924 52588
rect 19628 51308 19684 51310
rect 19708 51308 19764 51310
rect 19788 51308 19844 51310
rect 19868 51308 19924 51310
rect 19628 51256 19654 51308
rect 19654 51256 19684 51308
rect 19708 51256 19718 51308
rect 19718 51256 19764 51308
rect 19788 51256 19834 51308
rect 19834 51256 19844 51308
rect 19868 51256 19898 51308
rect 19898 51256 19924 51308
rect 19628 51254 19684 51256
rect 19708 51254 19764 51256
rect 19788 51254 19844 51256
rect 19868 51254 19924 51256
rect 19628 49976 19684 49978
rect 19708 49976 19764 49978
rect 19788 49976 19844 49978
rect 19868 49976 19924 49978
rect 19628 49924 19654 49976
rect 19654 49924 19684 49976
rect 19708 49924 19718 49976
rect 19718 49924 19764 49976
rect 19788 49924 19834 49976
rect 19834 49924 19844 49976
rect 19868 49924 19898 49976
rect 19898 49924 19924 49976
rect 19628 49922 19684 49924
rect 19708 49922 19764 49924
rect 19788 49922 19844 49924
rect 19868 49922 19924 49924
rect 19628 48644 19684 48646
rect 19708 48644 19764 48646
rect 19788 48644 19844 48646
rect 19868 48644 19924 48646
rect 19628 48592 19654 48644
rect 19654 48592 19684 48644
rect 19708 48592 19718 48644
rect 19718 48592 19764 48644
rect 19788 48592 19834 48644
rect 19834 48592 19844 48644
rect 19868 48592 19898 48644
rect 19898 48592 19924 48644
rect 19628 48590 19684 48592
rect 19708 48590 19764 48592
rect 19788 48590 19844 48592
rect 19868 48590 19924 48592
rect 19628 47312 19684 47314
rect 19708 47312 19764 47314
rect 19788 47312 19844 47314
rect 19868 47312 19924 47314
rect 19628 47260 19654 47312
rect 19654 47260 19684 47312
rect 19708 47260 19718 47312
rect 19718 47260 19764 47312
rect 19788 47260 19834 47312
rect 19834 47260 19844 47312
rect 19868 47260 19898 47312
rect 19898 47260 19924 47312
rect 19628 47258 19684 47260
rect 19708 47258 19764 47260
rect 19788 47258 19844 47260
rect 19868 47258 19924 47260
rect 19628 45980 19684 45982
rect 19708 45980 19764 45982
rect 19788 45980 19844 45982
rect 19868 45980 19924 45982
rect 19628 45928 19654 45980
rect 19654 45928 19684 45980
rect 19708 45928 19718 45980
rect 19718 45928 19764 45980
rect 19788 45928 19834 45980
rect 19834 45928 19844 45980
rect 19868 45928 19898 45980
rect 19898 45928 19924 45980
rect 19628 45926 19684 45928
rect 19708 45926 19764 45928
rect 19788 45926 19844 45928
rect 19868 45926 19924 45928
rect 19628 44648 19684 44650
rect 19708 44648 19764 44650
rect 19788 44648 19844 44650
rect 19868 44648 19924 44650
rect 19628 44596 19654 44648
rect 19654 44596 19684 44648
rect 19708 44596 19718 44648
rect 19718 44596 19764 44648
rect 19788 44596 19834 44648
rect 19834 44596 19844 44648
rect 19868 44596 19898 44648
rect 19898 44596 19924 44648
rect 19628 44594 19684 44596
rect 19708 44594 19764 44596
rect 19788 44594 19844 44596
rect 19868 44594 19924 44596
rect 19628 43316 19684 43318
rect 19708 43316 19764 43318
rect 19788 43316 19844 43318
rect 19868 43316 19924 43318
rect 19628 43264 19654 43316
rect 19654 43264 19684 43316
rect 19708 43264 19718 43316
rect 19718 43264 19764 43316
rect 19788 43264 19834 43316
rect 19834 43264 19844 43316
rect 19868 43264 19898 43316
rect 19898 43264 19924 43316
rect 19628 43262 19684 43264
rect 19708 43262 19764 43264
rect 19788 43262 19844 43264
rect 19868 43262 19924 43264
rect 19628 41984 19684 41986
rect 19708 41984 19764 41986
rect 19788 41984 19844 41986
rect 19868 41984 19924 41986
rect 19628 41932 19654 41984
rect 19654 41932 19684 41984
rect 19708 41932 19718 41984
rect 19718 41932 19764 41984
rect 19788 41932 19834 41984
rect 19834 41932 19844 41984
rect 19868 41932 19898 41984
rect 19898 41932 19924 41984
rect 19628 41930 19684 41932
rect 19708 41930 19764 41932
rect 19788 41930 19844 41932
rect 19868 41930 19924 41932
rect 19628 40652 19684 40654
rect 19708 40652 19764 40654
rect 19788 40652 19844 40654
rect 19868 40652 19924 40654
rect 19628 40600 19654 40652
rect 19654 40600 19684 40652
rect 19708 40600 19718 40652
rect 19718 40600 19764 40652
rect 19788 40600 19834 40652
rect 19834 40600 19844 40652
rect 19868 40600 19898 40652
rect 19898 40600 19924 40652
rect 19628 40598 19684 40600
rect 19708 40598 19764 40600
rect 19788 40598 19844 40600
rect 19868 40598 19924 40600
rect 19628 39320 19684 39322
rect 19708 39320 19764 39322
rect 19788 39320 19844 39322
rect 19868 39320 19924 39322
rect 19628 39268 19654 39320
rect 19654 39268 19684 39320
rect 19708 39268 19718 39320
rect 19718 39268 19764 39320
rect 19788 39268 19834 39320
rect 19834 39268 19844 39320
rect 19868 39268 19898 39320
rect 19898 39268 19924 39320
rect 19628 39266 19684 39268
rect 19708 39266 19764 39268
rect 19788 39266 19844 39268
rect 19868 39266 19924 39268
rect 19628 37988 19684 37990
rect 19708 37988 19764 37990
rect 19788 37988 19844 37990
rect 19868 37988 19924 37990
rect 19628 37936 19654 37988
rect 19654 37936 19684 37988
rect 19708 37936 19718 37988
rect 19718 37936 19764 37988
rect 19788 37936 19834 37988
rect 19834 37936 19844 37988
rect 19868 37936 19898 37988
rect 19898 37936 19924 37988
rect 19628 37934 19684 37936
rect 19708 37934 19764 37936
rect 19788 37934 19844 37936
rect 19868 37934 19924 37936
rect 19628 36656 19684 36658
rect 19708 36656 19764 36658
rect 19788 36656 19844 36658
rect 19868 36656 19924 36658
rect 19628 36604 19654 36656
rect 19654 36604 19684 36656
rect 19708 36604 19718 36656
rect 19718 36604 19764 36656
rect 19788 36604 19834 36656
rect 19834 36604 19844 36656
rect 19868 36604 19898 36656
rect 19898 36604 19924 36656
rect 19628 36602 19684 36604
rect 19708 36602 19764 36604
rect 19788 36602 19844 36604
rect 19868 36602 19924 36604
rect 19628 35324 19684 35326
rect 19708 35324 19764 35326
rect 19788 35324 19844 35326
rect 19868 35324 19924 35326
rect 19628 35272 19654 35324
rect 19654 35272 19684 35324
rect 19708 35272 19718 35324
rect 19718 35272 19764 35324
rect 19788 35272 19834 35324
rect 19834 35272 19844 35324
rect 19868 35272 19898 35324
rect 19898 35272 19924 35324
rect 19628 35270 19684 35272
rect 19708 35270 19764 35272
rect 19788 35270 19844 35272
rect 19868 35270 19924 35272
rect 19628 33992 19684 33994
rect 19708 33992 19764 33994
rect 19788 33992 19844 33994
rect 19868 33992 19924 33994
rect 19628 33940 19654 33992
rect 19654 33940 19684 33992
rect 19708 33940 19718 33992
rect 19718 33940 19764 33992
rect 19788 33940 19834 33992
rect 19834 33940 19844 33992
rect 19868 33940 19898 33992
rect 19898 33940 19924 33992
rect 19628 33938 19684 33940
rect 19708 33938 19764 33940
rect 19788 33938 19844 33940
rect 19868 33938 19924 33940
rect 19628 32660 19684 32662
rect 19708 32660 19764 32662
rect 19788 32660 19844 32662
rect 19868 32660 19924 32662
rect 19628 32608 19654 32660
rect 19654 32608 19684 32660
rect 19708 32608 19718 32660
rect 19718 32608 19764 32660
rect 19788 32608 19834 32660
rect 19834 32608 19844 32660
rect 19868 32608 19898 32660
rect 19898 32608 19924 32660
rect 19628 32606 19684 32608
rect 19708 32606 19764 32608
rect 19788 32606 19844 32608
rect 19868 32606 19924 32608
rect 19628 31328 19684 31330
rect 19708 31328 19764 31330
rect 19788 31328 19844 31330
rect 19868 31328 19924 31330
rect 19628 31276 19654 31328
rect 19654 31276 19684 31328
rect 19708 31276 19718 31328
rect 19718 31276 19764 31328
rect 19788 31276 19834 31328
rect 19834 31276 19844 31328
rect 19868 31276 19898 31328
rect 19898 31276 19924 31328
rect 19628 31274 19684 31276
rect 19708 31274 19764 31276
rect 19788 31274 19844 31276
rect 19868 31274 19924 31276
rect 19628 29996 19684 29998
rect 19708 29996 19764 29998
rect 19788 29996 19844 29998
rect 19868 29996 19924 29998
rect 19628 29944 19654 29996
rect 19654 29944 19684 29996
rect 19708 29944 19718 29996
rect 19718 29944 19764 29996
rect 19788 29944 19834 29996
rect 19834 29944 19844 29996
rect 19868 29944 19898 29996
rect 19898 29944 19924 29996
rect 19628 29942 19684 29944
rect 19708 29942 19764 29944
rect 19788 29942 19844 29944
rect 19868 29942 19924 29944
rect 19628 28664 19684 28666
rect 19708 28664 19764 28666
rect 19788 28664 19844 28666
rect 19868 28664 19924 28666
rect 19628 28612 19654 28664
rect 19654 28612 19684 28664
rect 19708 28612 19718 28664
rect 19718 28612 19764 28664
rect 19788 28612 19834 28664
rect 19834 28612 19844 28664
rect 19868 28612 19898 28664
rect 19898 28612 19924 28664
rect 19628 28610 19684 28612
rect 19708 28610 19764 28612
rect 19788 28610 19844 28612
rect 19868 28610 19924 28612
rect 19628 27332 19684 27334
rect 19708 27332 19764 27334
rect 19788 27332 19844 27334
rect 19868 27332 19924 27334
rect 19628 27280 19654 27332
rect 19654 27280 19684 27332
rect 19708 27280 19718 27332
rect 19718 27280 19764 27332
rect 19788 27280 19834 27332
rect 19834 27280 19844 27332
rect 19868 27280 19898 27332
rect 19898 27280 19924 27332
rect 19628 27278 19684 27280
rect 19708 27278 19764 27280
rect 19788 27278 19844 27280
rect 19868 27278 19924 27280
rect 19628 26000 19684 26002
rect 19708 26000 19764 26002
rect 19788 26000 19844 26002
rect 19868 26000 19924 26002
rect 19628 25948 19654 26000
rect 19654 25948 19684 26000
rect 19708 25948 19718 26000
rect 19718 25948 19764 26000
rect 19788 25948 19834 26000
rect 19834 25948 19844 26000
rect 19868 25948 19898 26000
rect 19898 25948 19924 26000
rect 19628 25946 19684 25948
rect 19708 25946 19764 25948
rect 19788 25946 19844 25948
rect 19868 25946 19924 25948
rect 19628 24668 19684 24670
rect 19708 24668 19764 24670
rect 19788 24668 19844 24670
rect 19868 24668 19924 24670
rect 19628 24616 19654 24668
rect 19654 24616 19684 24668
rect 19708 24616 19718 24668
rect 19718 24616 19764 24668
rect 19788 24616 19834 24668
rect 19834 24616 19844 24668
rect 19868 24616 19898 24668
rect 19898 24616 19924 24668
rect 19628 24614 19684 24616
rect 19708 24614 19764 24616
rect 19788 24614 19844 24616
rect 19868 24614 19924 24616
rect 19628 23336 19684 23338
rect 19708 23336 19764 23338
rect 19788 23336 19844 23338
rect 19868 23336 19924 23338
rect 19628 23284 19654 23336
rect 19654 23284 19684 23336
rect 19708 23284 19718 23336
rect 19718 23284 19764 23336
rect 19788 23284 19834 23336
rect 19834 23284 19844 23336
rect 19868 23284 19898 23336
rect 19898 23284 19924 23336
rect 19628 23282 19684 23284
rect 19708 23282 19764 23284
rect 19788 23282 19844 23284
rect 19868 23282 19924 23284
rect 19628 22004 19684 22006
rect 19708 22004 19764 22006
rect 19788 22004 19844 22006
rect 19868 22004 19924 22006
rect 19628 21952 19654 22004
rect 19654 21952 19684 22004
rect 19708 21952 19718 22004
rect 19718 21952 19764 22004
rect 19788 21952 19834 22004
rect 19834 21952 19844 22004
rect 19868 21952 19898 22004
rect 19898 21952 19924 22004
rect 19628 21950 19684 21952
rect 19708 21950 19764 21952
rect 19788 21950 19844 21952
rect 19868 21950 19924 21952
rect 19628 20672 19684 20674
rect 19708 20672 19764 20674
rect 19788 20672 19844 20674
rect 19868 20672 19924 20674
rect 19628 20620 19654 20672
rect 19654 20620 19684 20672
rect 19708 20620 19718 20672
rect 19718 20620 19764 20672
rect 19788 20620 19834 20672
rect 19834 20620 19844 20672
rect 19868 20620 19898 20672
rect 19898 20620 19924 20672
rect 19628 20618 19684 20620
rect 19708 20618 19764 20620
rect 19788 20618 19844 20620
rect 19868 20618 19924 20620
rect 19628 19340 19684 19342
rect 19708 19340 19764 19342
rect 19788 19340 19844 19342
rect 19868 19340 19924 19342
rect 19628 19288 19654 19340
rect 19654 19288 19684 19340
rect 19708 19288 19718 19340
rect 19718 19288 19764 19340
rect 19788 19288 19834 19340
rect 19834 19288 19844 19340
rect 19868 19288 19898 19340
rect 19898 19288 19924 19340
rect 19628 19286 19684 19288
rect 19708 19286 19764 19288
rect 19788 19286 19844 19288
rect 19868 19286 19924 19288
rect 19628 18008 19684 18010
rect 19708 18008 19764 18010
rect 19788 18008 19844 18010
rect 19868 18008 19924 18010
rect 19628 17956 19654 18008
rect 19654 17956 19684 18008
rect 19708 17956 19718 18008
rect 19718 17956 19764 18008
rect 19788 17956 19834 18008
rect 19834 17956 19844 18008
rect 19868 17956 19898 18008
rect 19898 17956 19924 18008
rect 19628 17954 19684 17956
rect 19708 17954 19764 17956
rect 19788 17954 19844 17956
rect 19868 17954 19924 17956
rect 19628 16676 19684 16678
rect 19708 16676 19764 16678
rect 19788 16676 19844 16678
rect 19868 16676 19924 16678
rect 19628 16624 19654 16676
rect 19654 16624 19684 16676
rect 19708 16624 19718 16676
rect 19718 16624 19764 16676
rect 19788 16624 19834 16676
rect 19834 16624 19844 16676
rect 19868 16624 19898 16676
rect 19898 16624 19924 16676
rect 19628 16622 19684 16624
rect 19708 16622 19764 16624
rect 19788 16622 19844 16624
rect 19868 16622 19924 16624
rect 19628 15344 19684 15346
rect 19708 15344 19764 15346
rect 19788 15344 19844 15346
rect 19868 15344 19924 15346
rect 19628 15292 19654 15344
rect 19654 15292 19684 15344
rect 19708 15292 19718 15344
rect 19718 15292 19764 15344
rect 19788 15292 19834 15344
rect 19834 15292 19844 15344
rect 19868 15292 19898 15344
rect 19898 15292 19924 15344
rect 19628 15290 19684 15292
rect 19708 15290 19764 15292
rect 19788 15290 19844 15292
rect 19868 15290 19924 15292
rect 19628 14012 19684 14014
rect 19708 14012 19764 14014
rect 19788 14012 19844 14014
rect 19868 14012 19924 14014
rect 19628 13960 19654 14012
rect 19654 13960 19684 14012
rect 19708 13960 19718 14012
rect 19718 13960 19764 14012
rect 19788 13960 19834 14012
rect 19834 13960 19844 14012
rect 19868 13960 19898 14012
rect 19898 13960 19924 14012
rect 19628 13958 19684 13960
rect 19708 13958 19764 13960
rect 19788 13958 19844 13960
rect 19868 13958 19924 13960
rect 19628 12680 19684 12682
rect 19708 12680 19764 12682
rect 19788 12680 19844 12682
rect 19868 12680 19924 12682
rect 19628 12628 19654 12680
rect 19654 12628 19684 12680
rect 19708 12628 19718 12680
rect 19718 12628 19764 12680
rect 19788 12628 19834 12680
rect 19834 12628 19844 12680
rect 19868 12628 19898 12680
rect 19898 12628 19924 12680
rect 19628 12626 19684 12628
rect 19708 12626 19764 12628
rect 19788 12626 19844 12628
rect 19868 12626 19924 12628
rect 19628 11348 19684 11350
rect 19708 11348 19764 11350
rect 19788 11348 19844 11350
rect 19868 11348 19924 11350
rect 19628 11296 19654 11348
rect 19654 11296 19684 11348
rect 19708 11296 19718 11348
rect 19718 11296 19764 11348
rect 19788 11296 19834 11348
rect 19834 11296 19844 11348
rect 19868 11296 19898 11348
rect 19898 11296 19924 11348
rect 19628 11294 19684 11296
rect 19708 11294 19764 11296
rect 19788 11294 19844 11296
rect 19868 11294 19924 11296
rect 19628 10016 19684 10018
rect 19708 10016 19764 10018
rect 19788 10016 19844 10018
rect 19868 10016 19924 10018
rect 19628 9964 19654 10016
rect 19654 9964 19684 10016
rect 19708 9964 19718 10016
rect 19718 9964 19764 10016
rect 19788 9964 19834 10016
rect 19834 9964 19844 10016
rect 19868 9964 19898 10016
rect 19898 9964 19924 10016
rect 19628 9962 19684 9964
rect 19708 9962 19764 9964
rect 19788 9962 19844 9964
rect 19868 9962 19924 9964
rect 19628 8684 19684 8686
rect 19708 8684 19764 8686
rect 19788 8684 19844 8686
rect 19868 8684 19924 8686
rect 19628 8632 19654 8684
rect 19654 8632 19684 8684
rect 19708 8632 19718 8684
rect 19718 8632 19764 8684
rect 19788 8632 19834 8684
rect 19834 8632 19844 8684
rect 19868 8632 19898 8684
rect 19898 8632 19924 8684
rect 19628 8630 19684 8632
rect 19708 8630 19764 8632
rect 19788 8630 19844 8632
rect 19868 8630 19924 8632
rect 19628 7352 19684 7354
rect 19708 7352 19764 7354
rect 19788 7352 19844 7354
rect 19868 7352 19924 7354
rect 19628 7300 19654 7352
rect 19654 7300 19684 7352
rect 19708 7300 19718 7352
rect 19718 7300 19764 7352
rect 19788 7300 19834 7352
rect 19834 7300 19844 7352
rect 19868 7300 19898 7352
rect 19898 7300 19924 7352
rect 19628 7298 19684 7300
rect 19708 7298 19764 7300
rect 19788 7298 19844 7300
rect 19868 7298 19924 7300
rect 19628 6020 19684 6022
rect 19708 6020 19764 6022
rect 19788 6020 19844 6022
rect 19868 6020 19924 6022
rect 19628 5968 19654 6020
rect 19654 5968 19684 6020
rect 19708 5968 19718 6020
rect 19718 5968 19764 6020
rect 19788 5968 19834 6020
rect 19834 5968 19844 6020
rect 19868 5968 19898 6020
rect 19898 5968 19924 6020
rect 19628 5966 19684 5968
rect 19708 5966 19764 5968
rect 19788 5966 19844 5968
rect 19868 5966 19924 5968
rect 19628 4688 19684 4690
rect 19708 4688 19764 4690
rect 19788 4688 19844 4690
rect 19868 4688 19924 4690
rect 19628 4636 19654 4688
rect 19654 4636 19684 4688
rect 19708 4636 19718 4688
rect 19718 4636 19764 4688
rect 19788 4636 19834 4688
rect 19834 4636 19844 4688
rect 19868 4636 19898 4688
rect 19898 4636 19924 4688
rect 19628 4634 19684 4636
rect 19708 4634 19764 4636
rect 19788 4634 19844 4636
rect 19868 4634 19924 4636
rect 19628 3356 19684 3358
rect 19708 3356 19764 3358
rect 19788 3356 19844 3358
rect 19868 3356 19924 3358
rect 19628 3304 19654 3356
rect 19654 3304 19684 3356
rect 19708 3304 19718 3356
rect 19718 3304 19764 3356
rect 19788 3304 19834 3356
rect 19834 3304 19844 3356
rect 19868 3304 19898 3356
rect 19898 3304 19924 3356
rect 19628 3302 19684 3304
rect 19708 3302 19764 3304
rect 19788 3302 19844 3304
rect 19868 3302 19924 3304
rect 34988 57302 35044 57304
rect 35068 57302 35124 57304
rect 35148 57302 35204 57304
rect 35228 57302 35284 57304
rect 34988 57250 35014 57302
rect 35014 57250 35044 57302
rect 35068 57250 35078 57302
rect 35078 57250 35124 57302
rect 35148 57250 35194 57302
rect 35194 57250 35204 57302
rect 35228 57250 35258 57302
rect 35258 57250 35284 57302
rect 34988 57248 35044 57250
rect 35068 57248 35124 57250
rect 35148 57248 35204 57250
rect 35228 57248 35284 57250
rect 34988 55970 35044 55972
rect 35068 55970 35124 55972
rect 35148 55970 35204 55972
rect 35228 55970 35284 55972
rect 34988 55918 35014 55970
rect 35014 55918 35044 55970
rect 35068 55918 35078 55970
rect 35078 55918 35124 55970
rect 35148 55918 35194 55970
rect 35194 55918 35204 55970
rect 35228 55918 35258 55970
rect 35258 55918 35284 55970
rect 34988 55916 35044 55918
rect 35068 55916 35124 55918
rect 35148 55916 35204 55918
rect 35228 55916 35284 55918
rect 34988 54638 35044 54640
rect 35068 54638 35124 54640
rect 35148 54638 35204 54640
rect 35228 54638 35284 54640
rect 34988 54586 35014 54638
rect 35014 54586 35044 54638
rect 35068 54586 35078 54638
rect 35078 54586 35124 54638
rect 35148 54586 35194 54638
rect 35194 54586 35204 54638
rect 35228 54586 35258 54638
rect 35258 54586 35284 54638
rect 34988 54584 35044 54586
rect 35068 54584 35124 54586
rect 35148 54584 35204 54586
rect 35228 54584 35284 54586
rect 34988 53306 35044 53308
rect 35068 53306 35124 53308
rect 35148 53306 35204 53308
rect 35228 53306 35284 53308
rect 34988 53254 35014 53306
rect 35014 53254 35044 53306
rect 35068 53254 35078 53306
rect 35078 53254 35124 53306
rect 35148 53254 35194 53306
rect 35194 53254 35204 53306
rect 35228 53254 35258 53306
rect 35258 53254 35284 53306
rect 34988 53252 35044 53254
rect 35068 53252 35124 53254
rect 35148 53252 35204 53254
rect 35228 53252 35284 53254
rect 34988 51974 35044 51976
rect 35068 51974 35124 51976
rect 35148 51974 35204 51976
rect 35228 51974 35284 51976
rect 34988 51922 35014 51974
rect 35014 51922 35044 51974
rect 35068 51922 35078 51974
rect 35078 51922 35124 51974
rect 35148 51922 35194 51974
rect 35194 51922 35204 51974
rect 35228 51922 35258 51974
rect 35258 51922 35284 51974
rect 34988 51920 35044 51922
rect 35068 51920 35124 51922
rect 35148 51920 35204 51922
rect 35228 51920 35284 51922
rect 34988 50642 35044 50644
rect 35068 50642 35124 50644
rect 35148 50642 35204 50644
rect 35228 50642 35284 50644
rect 34988 50590 35014 50642
rect 35014 50590 35044 50642
rect 35068 50590 35078 50642
rect 35078 50590 35124 50642
rect 35148 50590 35194 50642
rect 35194 50590 35204 50642
rect 35228 50590 35258 50642
rect 35258 50590 35284 50642
rect 34988 50588 35044 50590
rect 35068 50588 35124 50590
rect 35148 50588 35204 50590
rect 35228 50588 35284 50590
rect 34988 49310 35044 49312
rect 35068 49310 35124 49312
rect 35148 49310 35204 49312
rect 35228 49310 35284 49312
rect 34988 49258 35014 49310
rect 35014 49258 35044 49310
rect 35068 49258 35078 49310
rect 35078 49258 35124 49310
rect 35148 49258 35194 49310
rect 35194 49258 35204 49310
rect 35228 49258 35258 49310
rect 35258 49258 35284 49310
rect 34988 49256 35044 49258
rect 35068 49256 35124 49258
rect 35148 49256 35204 49258
rect 35228 49256 35284 49258
rect 34988 47978 35044 47980
rect 35068 47978 35124 47980
rect 35148 47978 35204 47980
rect 35228 47978 35284 47980
rect 34988 47926 35014 47978
rect 35014 47926 35044 47978
rect 35068 47926 35078 47978
rect 35078 47926 35124 47978
rect 35148 47926 35194 47978
rect 35194 47926 35204 47978
rect 35228 47926 35258 47978
rect 35258 47926 35284 47978
rect 34988 47924 35044 47926
rect 35068 47924 35124 47926
rect 35148 47924 35204 47926
rect 35228 47924 35284 47926
rect 34988 46646 35044 46648
rect 35068 46646 35124 46648
rect 35148 46646 35204 46648
rect 35228 46646 35284 46648
rect 34988 46594 35014 46646
rect 35014 46594 35044 46646
rect 35068 46594 35078 46646
rect 35078 46594 35124 46646
rect 35148 46594 35194 46646
rect 35194 46594 35204 46646
rect 35228 46594 35258 46646
rect 35258 46594 35284 46646
rect 34988 46592 35044 46594
rect 35068 46592 35124 46594
rect 35148 46592 35204 46594
rect 35228 46592 35284 46594
rect 34988 45314 35044 45316
rect 35068 45314 35124 45316
rect 35148 45314 35204 45316
rect 35228 45314 35284 45316
rect 34988 45262 35014 45314
rect 35014 45262 35044 45314
rect 35068 45262 35078 45314
rect 35078 45262 35124 45314
rect 35148 45262 35194 45314
rect 35194 45262 35204 45314
rect 35228 45262 35258 45314
rect 35258 45262 35284 45314
rect 34988 45260 35044 45262
rect 35068 45260 35124 45262
rect 35148 45260 35204 45262
rect 35228 45260 35284 45262
rect 34988 43982 35044 43984
rect 35068 43982 35124 43984
rect 35148 43982 35204 43984
rect 35228 43982 35284 43984
rect 34988 43930 35014 43982
rect 35014 43930 35044 43982
rect 35068 43930 35078 43982
rect 35078 43930 35124 43982
rect 35148 43930 35194 43982
rect 35194 43930 35204 43982
rect 35228 43930 35258 43982
rect 35258 43930 35284 43982
rect 34988 43928 35044 43930
rect 35068 43928 35124 43930
rect 35148 43928 35204 43930
rect 35228 43928 35284 43930
rect 34988 42650 35044 42652
rect 35068 42650 35124 42652
rect 35148 42650 35204 42652
rect 35228 42650 35284 42652
rect 34988 42598 35014 42650
rect 35014 42598 35044 42650
rect 35068 42598 35078 42650
rect 35078 42598 35124 42650
rect 35148 42598 35194 42650
rect 35194 42598 35204 42650
rect 35228 42598 35258 42650
rect 35258 42598 35284 42650
rect 34988 42596 35044 42598
rect 35068 42596 35124 42598
rect 35148 42596 35204 42598
rect 35228 42596 35284 42598
rect 34988 41318 35044 41320
rect 35068 41318 35124 41320
rect 35148 41318 35204 41320
rect 35228 41318 35284 41320
rect 34988 41266 35014 41318
rect 35014 41266 35044 41318
rect 35068 41266 35078 41318
rect 35078 41266 35124 41318
rect 35148 41266 35194 41318
rect 35194 41266 35204 41318
rect 35228 41266 35258 41318
rect 35258 41266 35284 41318
rect 34988 41264 35044 41266
rect 35068 41264 35124 41266
rect 35148 41264 35204 41266
rect 35228 41264 35284 41266
rect 34988 39986 35044 39988
rect 35068 39986 35124 39988
rect 35148 39986 35204 39988
rect 35228 39986 35284 39988
rect 34988 39934 35014 39986
rect 35014 39934 35044 39986
rect 35068 39934 35078 39986
rect 35078 39934 35124 39986
rect 35148 39934 35194 39986
rect 35194 39934 35204 39986
rect 35228 39934 35258 39986
rect 35258 39934 35284 39986
rect 34988 39932 35044 39934
rect 35068 39932 35124 39934
rect 35148 39932 35204 39934
rect 35228 39932 35284 39934
rect 34988 38654 35044 38656
rect 35068 38654 35124 38656
rect 35148 38654 35204 38656
rect 35228 38654 35284 38656
rect 34988 38602 35014 38654
rect 35014 38602 35044 38654
rect 35068 38602 35078 38654
rect 35078 38602 35124 38654
rect 35148 38602 35194 38654
rect 35194 38602 35204 38654
rect 35228 38602 35258 38654
rect 35258 38602 35284 38654
rect 34988 38600 35044 38602
rect 35068 38600 35124 38602
rect 35148 38600 35204 38602
rect 35228 38600 35284 38602
rect 34988 37322 35044 37324
rect 35068 37322 35124 37324
rect 35148 37322 35204 37324
rect 35228 37322 35284 37324
rect 34988 37270 35014 37322
rect 35014 37270 35044 37322
rect 35068 37270 35078 37322
rect 35078 37270 35124 37322
rect 35148 37270 35194 37322
rect 35194 37270 35204 37322
rect 35228 37270 35258 37322
rect 35258 37270 35284 37322
rect 34988 37268 35044 37270
rect 35068 37268 35124 37270
rect 35148 37268 35204 37270
rect 35228 37268 35284 37270
rect 34988 35990 35044 35992
rect 35068 35990 35124 35992
rect 35148 35990 35204 35992
rect 35228 35990 35284 35992
rect 34988 35938 35014 35990
rect 35014 35938 35044 35990
rect 35068 35938 35078 35990
rect 35078 35938 35124 35990
rect 35148 35938 35194 35990
rect 35194 35938 35204 35990
rect 35228 35938 35258 35990
rect 35258 35938 35284 35990
rect 34988 35936 35044 35938
rect 35068 35936 35124 35938
rect 35148 35936 35204 35938
rect 35228 35936 35284 35938
rect 34988 34658 35044 34660
rect 35068 34658 35124 34660
rect 35148 34658 35204 34660
rect 35228 34658 35284 34660
rect 34988 34606 35014 34658
rect 35014 34606 35044 34658
rect 35068 34606 35078 34658
rect 35078 34606 35124 34658
rect 35148 34606 35194 34658
rect 35194 34606 35204 34658
rect 35228 34606 35258 34658
rect 35258 34606 35284 34658
rect 34988 34604 35044 34606
rect 35068 34604 35124 34606
rect 35148 34604 35204 34606
rect 35228 34604 35284 34606
rect 34988 33326 35044 33328
rect 35068 33326 35124 33328
rect 35148 33326 35204 33328
rect 35228 33326 35284 33328
rect 34988 33274 35014 33326
rect 35014 33274 35044 33326
rect 35068 33274 35078 33326
rect 35078 33274 35124 33326
rect 35148 33274 35194 33326
rect 35194 33274 35204 33326
rect 35228 33274 35258 33326
rect 35258 33274 35284 33326
rect 34988 33272 35044 33274
rect 35068 33272 35124 33274
rect 35148 33272 35204 33274
rect 35228 33272 35284 33274
rect 34988 31994 35044 31996
rect 35068 31994 35124 31996
rect 35148 31994 35204 31996
rect 35228 31994 35284 31996
rect 34988 31942 35014 31994
rect 35014 31942 35044 31994
rect 35068 31942 35078 31994
rect 35078 31942 35124 31994
rect 35148 31942 35194 31994
rect 35194 31942 35204 31994
rect 35228 31942 35258 31994
rect 35258 31942 35284 31994
rect 34988 31940 35044 31942
rect 35068 31940 35124 31942
rect 35148 31940 35204 31942
rect 35228 31940 35284 31942
rect 34988 30662 35044 30664
rect 35068 30662 35124 30664
rect 35148 30662 35204 30664
rect 35228 30662 35284 30664
rect 34988 30610 35014 30662
rect 35014 30610 35044 30662
rect 35068 30610 35078 30662
rect 35078 30610 35124 30662
rect 35148 30610 35194 30662
rect 35194 30610 35204 30662
rect 35228 30610 35258 30662
rect 35258 30610 35284 30662
rect 34988 30608 35044 30610
rect 35068 30608 35124 30610
rect 35148 30608 35204 30610
rect 35228 30608 35284 30610
rect 34988 29330 35044 29332
rect 35068 29330 35124 29332
rect 35148 29330 35204 29332
rect 35228 29330 35284 29332
rect 34988 29278 35014 29330
rect 35014 29278 35044 29330
rect 35068 29278 35078 29330
rect 35078 29278 35124 29330
rect 35148 29278 35194 29330
rect 35194 29278 35204 29330
rect 35228 29278 35258 29330
rect 35258 29278 35284 29330
rect 34988 29276 35044 29278
rect 35068 29276 35124 29278
rect 35148 29276 35204 29278
rect 35228 29276 35284 29278
rect 34988 27998 35044 28000
rect 35068 27998 35124 28000
rect 35148 27998 35204 28000
rect 35228 27998 35284 28000
rect 34988 27946 35014 27998
rect 35014 27946 35044 27998
rect 35068 27946 35078 27998
rect 35078 27946 35124 27998
rect 35148 27946 35194 27998
rect 35194 27946 35204 27998
rect 35228 27946 35258 27998
rect 35258 27946 35284 27998
rect 34988 27944 35044 27946
rect 35068 27944 35124 27946
rect 35148 27944 35204 27946
rect 35228 27944 35284 27946
rect 34988 26666 35044 26668
rect 35068 26666 35124 26668
rect 35148 26666 35204 26668
rect 35228 26666 35284 26668
rect 34988 26614 35014 26666
rect 35014 26614 35044 26666
rect 35068 26614 35078 26666
rect 35078 26614 35124 26666
rect 35148 26614 35194 26666
rect 35194 26614 35204 26666
rect 35228 26614 35258 26666
rect 35258 26614 35284 26666
rect 34988 26612 35044 26614
rect 35068 26612 35124 26614
rect 35148 26612 35204 26614
rect 35228 26612 35284 26614
rect 34988 25334 35044 25336
rect 35068 25334 35124 25336
rect 35148 25334 35204 25336
rect 35228 25334 35284 25336
rect 34988 25282 35014 25334
rect 35014 25282 35044 25334
rect 35068 25282 35078 25334
rect 35078 25282 35124 25334
rect 35148 25282 35194 25334
rect 35194 25282 35204 25334
rect 35228 25282 35258 25334
rect 35258 25282 35284 25334
rect 34988 25280 35044 25282
rect 35068 25280 35124 25282
rect 35148 25280 35204 25282
rect 35228 25280 35284 25282
rect 34988 24002 35044 24004
rect 35068 24002 35124 24004
rect 35148 24002 35204 24004
rect 35228 24002 35284 24004
rect 34988 23950 35014 24002
rect 35014 23950 35044 24002
rect 35068 23950 35078 24002
rect 35078 23950 35124 24002
rect 35148 23950 35194 24002
rect 35194 23950 35204 24002
rect 35228 23950 35258 24002
rect 35258 23950 35284 24002
rect 34988 23948 35044 23950
rect 35068 23948 35124 23950
rect 35148 23948 35204 23950
rect 35228 23948 35284 23950
rect 34988 22670 35044 22672
rect 35068 22670 35124 22672
rect 35148 22670 35204 22672
rect 35228 22670 35284 22672
rect 34988 22618 35014 22670
rect 35014 22618 35044 22670
rect 35068 22618 35078 22670
rect 35078 22618 35124 22670
rect 35148 22618 35194 22670
rect 35194 22618 35204 22670
rect 35228 22618 35258 22670
rect 35258 22618 35284 22670
rect 34988 22616 35044 22618
rect 35068 22616 35124 22618
rect 35148 22616 35204 22618
rect 35228 22616 35284 22618
rect 34988 21338 35044 21340
rect 35068 21338 35124 21340
rect 35148 21338 35204 21340
rect 35228 21338 35284 21340
rect 34988 21286 35014 21338
rect 35014 21286 35044 21338
rect 35068 21286 35078 21338
rect 35078 21286 35124 21338
rect 35148 21286 35194 21338
rect 35194 21286 35204 21338
rect 35228 21286 35258 21338
rect 35258 21286 35284 21338
rect 34988 21284 35044 21286
rect 35068 21284 35124 21286
rect 35148 21284 35204 21286
rect 35228 21284 35284 21286
rect 34988 20006 35044 20008
rect 35068 20006 35124 20008
rect 35148 20006 35204 20008
rect 35228 20006 35284 20008
rect 34988 19954 35014 20006
rect 35014 19954 35044 20006
rect 35068 19954 35078 20006
rect 35078 19954 35124 20006
rect 35148 19954 35194 20006
rect 35194 19954 35204 20006
rect 35228 19954 35258 20006
rect 35258 19954 35284 20006
rect 34988 19952 35044 19954
rect 35068 19952 35124 19954
rect 35148 19952 35204 19954
rect 35228 19952 35284 19954
rect 34988 18674 35044 18676
rect 35068 18674 35124 18676
rect 35148 18674 35204 18676
rect 35228 18674 35284 18676
rect 34988 18622 35014 18674
rect 35014 18622 35044 18674
rect 35068 18622 35078 18674
rect 35078 18622 35124 18674
rect 35148 18622 35194 18674
rect 35194 18622 35204 18674
rect 35228 18622 35258 18674
rect 35258 18622 35284 18674
rect 34988 18620 35044 18622
rect 35068 18620 35124 18622
rect 35148 18620 35204 18622
rect 35228 18620 35284 18622
rect 34988 17342 35044 17344
rect 35068 17342 35124 17344
rect 35148 17342 35204 17344
rect 35228 17342 35284 17344
rect 34988 17290 35014 17342
rect 35014 17290 35044 17342
rect 35068 17290 35078 17342
rect 35078 17290 35124 17342
rect 35148 17290 35194 17342
rect 35194 17290 35204 17342
rect 35228 17290 35258 17342
rect 35258 17290 35284 17342
rect 34988 17288 35044 17290
rect 35068 17288 35124 17290
rect 35148 17288 35204 17290
rect 35228 17288 35284 17290
rect 34988 16010 35044 16012
rect 35068 16010 35124 16012
rect 35148 16010 35204 16012
rect 35228 16010 35284 16012
rect 34988 15958 35014 16010
rect 35014 15958 35044 16010
rect 35068 15958 35078 16010
rect 35078 15958 35124 16010
rect 35148 15958 35194 16010
rect 35194 15958 35204 16010
rect 35228 15958 35258 16010
rect 35258 15958 35284 16010
rect 34988 15956 35044 15958
rect 35068 15956 35124 15958
rect 35148 15956 35204 15958
rect 35228 15956 35284 15958
rect 34988 14678 35044 14680
rect 35068 14678 35124 14680
rect 35148 14678 35204 14680
rect 35228 14678 35284 14680
rect 34988 14626 35014 14678
rect 35014 14626 35044 14678
rect 35068 14626 35078 14678
rect 35078 14626 35124 14678
rect 35148 14626 35194 14678
rect 35194 14626 35204 14678
rect 35228 14626 35258 14678
rect 35258 14626 35284 14678
rect 34988 14624 35044 14626
rect 35068 14624 35124 14626
rect 35148 14624 35204 14626
rect 35228 14624 35284 14626
rect 34988 13346 35044 13348
rect 35068 13346 35124 13348
rect 35148 13346 35204 13348
rect 35228 13346 35284 13348
rect 34988 13294 35014 13346
rect 35014 13294 35044 13346
rect 35068 13294 35078 13346
rect 35078 13294 35124 13346
rect 35148 13294 35194 13346
rect 35194 13294 35204 13346
rect 35228 13294 35258 13346
rect 35258 13294 35284 13346
rect 34988 13292 35044 13294
rect 35068 13292 35124 13294
rect 35148 13292 35204 13294
rect 35228 13292 35284 13294
rect 34988 12014 35044 12016
rect 35068 12014 35124 12016
rect 35148 12014 35204 12016
rect 35228 12014 35284 12016
rect 34988 11962 35014 12014
rect 35014 11962 35044 12014
rect 35068 11962 35078 12014
rect 35078 11962 35124 12014
rect 35148 11962 35194 12014
rect 35194 11962 35204 12014
rect 35228 11962 35258 12014
rect 35258 11962 35284 12014
rect 34988 11960 35044 11962
rect 35068 11960 35124 11962
rect 35148 11960 35204 11962
rect 35228 11960 35284 11962
rect 34988 10682 35044 10684
rect 35068 10682 35124 10684
rect 35148 10682 35204 10684
rect 35228 10682 35284 10684
rect 34988 10630 35014 10682
rect 35014 10630 35044 10682
rect 35068 10630 35078 10682
rect 35078 10630 35124 10682
rect 35148 10630 35194 10682
rect 35194 10630 35204 10682
rect 35228 10630 35258 10682
rect 35258 10630 35284 10682
rect 34988 10628 35044 10630
rect 35068 10628 35124 10630
rect 35148 10628 35204 10630
rect 35228 10628 35284 10630
rect 34988 9350 35044 9352
rect 35068 9350 35124 9352
rect 35148 9350 35204 9352
rect 35228 9350 35284 9352
rect 34988 9298 35014 9350
rect 35014 9298 35044 9350
rect 35068 9298 35078 9350
rect 35078 9298 35124 9350
rect 35148 9298 35194 9350
rect 35194 9298 35204 9350
rect 35228 9298 35258 9350
rect 35258 9298 35284 9350
rect 34988 9296 35044 9298
rect 35068 9296 35124 9298
rect 35148 9296 35204 9298
rect 35228 9296 35284 9298
rect 34988 8018 35044 8020
rect 35068 8018 35124 8020
rect 35148 8018 35204 8020
rect 35228 8018 35284 8020
rect 34988 7966 35014 8018
rect 35014 7966 35044 8018
rect 35068 7966 35078 8018
rect 35078 7966 35124 8018
rect 35148 7966 35194 8018
rect 35194 7966 35204 8018
rect 35228 7966 35258 8018
rect 35258 7966 35284 8018
rect 34988 7964 35044 7966
rect 35068 7964 35124 7966
rect 35148 7964 35204 7966
rect 35228 7964 35284 7966
rect 34484 2858 34540 2914
rect 34988 6686 35044 6688
rect 35068 6686 35124 6688
rect 35148 6686 35204 6688
rect 35228 6686 35284 6688
rect 34988 6634 35014 6686
rect 35014 6634 35044 6686
rect 35068 6634 35078 6686
rect 35078 6634 35124 6686
rect 35148 6634 35194 6686
rect 35194 6634 35204 6686
rect 35228 6634 35258 6686
rect 35258 6634 35284 6686
rect 34988 6632 35044 6634
rect 35068 6632 35124 6634
rect 35148 6632 35204 6634
rect 35228 6632 35284 6634
rect 34988 5354 35044 5356
rect 35068 5354 35124 5356
rect 35148 5354 35204 5356
rect 35228 5354 35284 5356
rect 34988 5302 35014 5354
rect 35014 5302 35044 5354
rect 35068 5302 35078 5354
rect 35078 5302 35124 5354
rect 35148 5302 35194 5354
rect 35194 5302 35204 5354
rect 35228 5302 35258 5354
rect 35258 5302 35284 5354
rect 34988 5300 35044 5302
rect 35068 5300 35124 5302
rect 35148 5300 35204 5302
rect 35228 5300 35284 5302
rect 34988 4022 35044 4024
rect 35068 4022 35124 4024
rect 35148 4022 35204 4024
rect 35228 4022 35284 4024
rect 34988 3970 35014 4022
rect 35014 3970 35044 4022
rect 35068 3970 35078 4022
rect 35078 3970 35124 4022
rect 35148 3970 35194 4022
rect 35194 3970 35204 4022
rect 35228 3970 35258 4022
rect 35258 3970 35284 4022
rect 34988 3968 35044 3970
rect 35068 3968 35124 3970
rect 35148 3968 35204 3970
rect 35228 3968 35284 3970
rect 35252 2858 35308 2914
rect 34988 2690 35044 2692
rect 35068 2690 35124 2692
rect 35148 2690 35204 2692
rect 35228 2690 35284 2692
rect 34988 2638 35014 2690
rect 35014 2638 35044 2690
rect 35068 2638 35078 2690
rect 35078 2638 35124 2690
rect 35148 2638 35194 2690
rect 35194 2638 35204 2690
rect 35228 2638 35258 2690
rect 35258 2638 35284 2690
rect 34988 2636 35044 2638
rect 35068 2636 35124 2638
rect 35148 2636 35204 2638
rect 35228 2636 35284 2638
rect 35156 2414 35212 2470
rect 35924 3154 35980 3210
rect 50348 56636 50404 56638
rect 50428 56636 50484 56638
rect 50508 56636 50564 56638
rect 50588 56636 50644 56638
rect 50348 56584 50374 56636
rect 50374 56584 50404 56636
rect 50428 56584 50438 56636
rect 50438 56584 50484 56636
rect 50508 56584 50554 56636
rect 50554 56584 50564 56636
rect 50588 56584 50618 56636
rect 50618 56584 50644 56636
rect 50348 56582 50404 56584
rect 50428 56582 50484 56584
rect 50508 56582 50564 56584
rect 50588 56582 50644 56584
rect 50348 55304 50404 55306
rect 50428 55304 50484 55306
rect 50508 55304 50564 55306
rect 50588 55304 50644 55306
rect 50348 55252 50374 55304
rect 50374 55252 50404 55304
rect 50428 55252 50438 55304
rect 50438 55252 50484 55304
rect 50508 55252 50554 55304
rect 50554 55252 50564 55304
rect 50588 55252 50618 55304
rect 50618 55252 50644 55304
rect 50348 55250 50404 55252
rect 50428 55250 50484 55252
rect 50508 55250 50564 55252
rect 50588 55250 50644 55252
rect 50348 53972 50404 53974
rect 50428 53972 50484 53974
rect 50508 53972 50564 53974
rect 50588 53972 50644 53974
rect 50348 53920 50374 53972
rect 50374 53920 50404 53972
rect 50428 53920 50438 53972
rect 50438 53920 50484 53972
rect 50508 53920 50554 53972
rect 50554 53920 50564 53972
rect 50588 53920 50618 53972
rect 50618 53920 50644 53972
rect 50348 53918 50404 53920
rect 50428 53918 50484 53920
rect 50508 53918 50564 53920
rect 50588 53918 50644 53920
rect 50348 52640 50404 52642
rect 50428 52640 50484 52642
rect 50508 52640 50564 52642
rect 50588 52640 50644 52642
rect 50348 52588 50374 52640
rect 50374 52588 50404 52640
rect 50428 52588 50438 52640
rect 50438 52588 50484 52640
rect 50508 52588 50554 52640
rect 50554 52588 50564 52640
rect 50588 52588 50618 52640
rect 50618 52588 50644 52640
rect 50348 52586 50404 52588
rect 50428 52586 50484 52588
rect 50508 52586 50564 52588
rect 50588 52586 50644 52588
rect 50348 51308 50404 51310
rect 50428 51308 50484 51310
rect 50508 51308 50564 51310
rect 50588 51308 50644 51310
rect 50348 51256 50374 51308
rect 50374 51256 50404 51308
rect 50428 51256 50438 51308
rect 50438 51256 50484 51308
rect 50508 51256 50554 51308
rect 50554 51256 50564 51308
rect 50588 51256 50618 51308
rect 50618 51256 50644 51308
rect 50348 51254 50404 51256
rect 50428 51254 50484 51256
rect 50508 51254 50564 51256
rect 50588 51254 50644 51256
rect 50348 49976 50404 49978
rect 50428 49976 50484 49978
rect 50508 49976 50564 49978
rect 50588 49976 50644 49978
rect 50348 49924 50374 49976
rect 50374 49924 50404 49976
rect 50428 49924 50438 49976
rect 50438 49924 50484 49976
rect 50508 49924 50554 49976
rect 50554 49924 50564 49976
rect 50588 49924 50618 49976
rect 50618 49924 50644 49976
rect 50348 49922 50404 49924
rect 50428 49922 50484 49924
rect 50508 49922 50564 49924
rect 50588 49922 50644 49924
rect 50348 48644 50404 48646
rect 50428 48644 50484 48646
rect 50508 48644 50564 48646
rect 50588 48644 50644 48646
rect 50348 48592 50374 48644
rect 50374 48592 50404 48644
rect 50428 48592 50438 48644
rect 50438 48592 50484 48644
rect 50508 48592 50554 48644
rect 50554 48592 50564 48644
rect 50588 48592 50618 48644
rect 50618 48592 50644 48644
rect 50348 48590 50404 48592
rect 50428 48590 50484 48592
rect 50508 48590 50564 48592
rect 50588 48590 50644 48592
rect 50348 47312 50404 47314
rect 50428 47312 50484 47314
rect 50508 47312 50564 47314
rect 50588 47312 50644 47314
rect 50348 47260 50374 47312
rect 50374 47260 50404 47312
rect 50428 47260 50438 47312
rect 50438 47260 50484 47312
rect 50508 47260 50554 47312
rect 50554 47260 50564 47312
rect 50588 47260 50618 47312
rect 50618 47260 50644 47312
rect 50348 47258 50404 47260
rect 50428 47258 50484 47260
rect 50508 47258 50564 47260
rect 50588 47258 50644 47260
rect 50348 45980 50404 45982
rect 50428 45980 50484 45982
rect 50508 45980 50564 45982
rect 50588 45980 50644 45982
rect 50348 45928 50374 45980
rect 50374 45928 50404 45980
rect 50428 45928 50438 45980
rect 50438 45928 50484 45980
rect 50508 45928 50554 45980
rect 50554 45928 50564 45980
rect 50588 45928 50618 45980
rect 50618 45928 50644 45980
rect 50348 45926 50404 45928
rect 50428 45926 50484 45928
rect 50508 45926 50564 45928
rect 50588 45926 50644 45928
rect 50348 44648 50404 44650
rect 50428 44648 50484 44650
rect 50508 44648 50564 44650
rect 50588 44648 50644 44650
rect 50348 44596 50374 44648
rect 50374 44596 50404 44648
rect 50428 44596 50438 44648
rect 50438 44596 50484 44648
rect 50508 44596 50554 44648
rect 50554 44596 50564 44648
rect 50588 44596 50618 44648
rect 50618 44596 50644 44648
rect 50348 44594 50404 44596
rect 50428 44594 50484 44596
rect 50508 44594 50564 44596
rect 50588 44594 50644 44596
rect 50348 43316 50404 43318
rect 50428 43316 50484 43318
rect 50508 43316 50564 43318
rect 50588 43316 50644 43318
rect 50348 43264 50374 43316
rect 50374 43264 50404 43316
rect 50428 43264 50438 43316
rect 50438 43264 50484 43316
rect 50508 43264 50554 43316
rect 50554 43264 50564 43316
rect 50588 43264 50618 43316
rect 50618 43264 50644 43316
rect 50348 43262 50404 43264
rect 50428 43262 50484 43264
rect 50508 43262 50564 43264
rect 50588 43262 50644 43264
rect 50348 41984 50404 41986
rect 50428 41984 50484 41986
rect 50508 41984 50564 41986
rect 50588 41984 50644 41986
rect 50348 41932 50374 41984
rect 50374 41932 50404 41984
rect 50428 41932 50438 41984
rect 50438 41932 50484 41984
rect 50508 41932 50554 41984
rect 50554 41932 50564 41984
rect 50588 41932 50618 41984
rect 50618 41932 50644 41984
rect 50348 41930 50404 41932
rect 50428 41930 50484 41932
rect 50508 41930 50564 41932
rect 50588 41930 50644 41932
rect 50348 40652 50404 40654
rect 50428 40652 50484 40654
rect 50508 40652 50564 40654
rect 50588 40652 50644 40654
rect 50348 40600 50374 40652
rect 50374 40600 50404 40652
rect 50428 40600 50438 40652
rect 50438 40600 50484 40652
rect 50508 40600 50554 40652
rect 50554 40600 50564 40652
rect 50588 40600 50618 40652
rect 50618 40600 50644 40652
rect 50348 40598 50404 40600
rect 50428 40598 50484 40600
rect 50508 40598 50564 40600
rect 50588 40598 50644 40600
rect 50348 39320 50404 39322
rect 50428 39320 50484 39322
rect 50508 39320 50564 39322
rect 50588 39320 50644 39322
rect 50348 39268 50374 39320
rect 50374 39268 50404 39320
rect 50428 39268 50438 39320
rect 50438 39268 50484 39320
rect 50508 39268 50554 39320
rect 50554 39268 50564 39320
rect 50588 39268 50618 39320
rect 50618 39268 50644 39320
rect 50348 39266 50404 39268
rect 50428 39266 50484 39268
rect 50508 39266 50564 39268
rect 50588 39266 50644 39268
rect 50348 37988 50404 37990
rect 50428 37988 50484 37990
rect 50508 37988 50564 37990
rect 50588 37988 50644 37990
rect 50348 37936 50374 37988
rect 50374 37936 50404 37988
rect 50428 37936 50438 37988
rect 50438 37936 50484 37988
rect 50508 37936 50554 37988
rect 50554 37936 50564 37988
rect 50588 37936 50618 37988
rect 50618 37936 50644 37988
rect 50348 37934 50404 37936
rect 50428 37934 50484 37936
rect 50508 37934 50564 37936
rect 50588 37934 50644 37936
rect 50348 36656 50404 36658
rect 50428 36656 50484 36658
rect 50508 36656 50564 36658
rect 50588 36656 50644 36658
rect 50348 36604 50374 36656
rect 50374 36604 50404 36656
rect 50428 36604 50438 36656
rect 50438 36604 50484 36656
rect 50508 36604 50554 36656
rect 50554 36604 50564 36656
rect 50588 36604 50618 36656
rect 50618 36604 50644 36656
rect 50348 36602 50404 36604
rect 50428 36602 50484 36604
rect 50508 36602 50564 36604
rect 50588 36602 50644 36604
rect 50348 35324 50404 35326
rect 50428 35324 50484 35326
rect 50508 35324 50564 35326
rect 50588 35324 50644 35326
rect 50348 35272 50374 35324
rect 50374 35272 50404 35324
rect 50428 35272 50438 35324
rect 50438 35272 50484 35324
rect 50508 35272 50554 35324
rect 50554 35272 50564 35324
rect 50588 35272 50618 35324
rect 50618 35272 50644 35324
rect 50348 35270 50404 35272
rect 50428 35270 50484 35272
rect 50508 35270 50564 35272
rect 50588 35270 50644 35272
rect 50348 33992 50404 33994
rect 50428 33992 50484 33994
rect 50508 33992 50564 33994
rect 50588 33992 50644 33994
rect 50348 33940 50374 33992
rect 50374 33940 50404 33992
rect 50428 33940 50438 33992
rect 50438 33940 50484 33992
rect 50508 33940 50554 33992
rect 50554 33940 50564 33992
rect 50588 33940 50618 33992
rect 50618 33940 50644 33992
rect 50348 33938 50404 33940
rect 50428 33938 50484 33940
rect 50508 33938 50564 33940
rect 50588 33938 50644 33940
rect 50348 32660 50404 32662
rect 50428 32660 50484 32662
rect 50508 32660 50564 32662
rect 50588 32660 50644 32662
rect 50348 32608 50374 32660
rect 50374 32608 50404 32660
rect 50428 32608 50438 32660
rect 50438 32608 50484 32660
rect 50508 32608 50554 32660
rect 50554 32608 50564 32660
rect 50588 32608 50618 32660
rect 50618 32608 50644 32660
rect 50348 32606 50404 32608
rect 50428 32606 50484 32608
rect 50508 32606 50564 32608
rect 50588 32606 50644 32608
rect 50348 31328 50404 31330
rect 50428 31328 50484 31330
rect 50508 31328 50564 31330
rect 50588 31328 50644 31330
rect 50348 31276 50374 31328
rect 50374 31276 50404 31328
rect 50428 31276 50438 31328
rect 50438 31276 50484 31328
rect 50508 31276 50554 31328
rect 50554 31276 50564 31328
rect 50588 31276 50618 31328
rect 50618 31276 50644 31328
rect 50348 31274 50404 31276
rect 50428 31274 50484 31276
rect 50508 31274 50564 31276
rect 50588 31274 50644 31276
rect 50348 29996 50404 29998
rect 50428 29996 50484 29998
rect 50508 29996 50564 29998
rect 50588 29996 50644 29998
rect 50348 29944 50374 29996
rect 50374 29944 50404 29996
rect 50428 29944 50438 29996
rect 50438 29944 50484 29996
rect 50508 29944 50554 29996
rect 50554 29944 50564 29996
rect 50588 29944 50618 29996
rect 50618 29944 50644 29996
rect 50348 29942 50404 29944
rect 50428 29942 50484 29944
rect 50508 29942 50564 29944
rect 50588 29942 50644 29944
rect 50348 28664 50404 28666
rect 50428 28664 50484 28666
rect 50508 28664 50564 28666
rect 50588 28664 50644 28666
rect 50348 28612 50374 28664
rect 50374 28612 50404 28664
rect 50428 28612 50438 28664
rect 50438 28612 50484 28664
rect 50508 28612 50554 28664
rect 50554 28612 50564 28664
rect 50588 28612 50618 28664
rect 50618 28612 50644 28664
rect 50348 28610 50404 28612
rect 50428 28610 50484 28612
rect 50508 28610 50564 28612
rect 50588 28610 50644 28612
rect 50348 27332 50404 27334
rect 50428 27332 50484 27334
rect 50508 27332 50564 27334
rect 50588 27332 50644 27334
rect 50348 27280 50374 27332
rect 50374 27280 50404 27332
rect 50428 27280 50438 27332
rect 50438 27280 50484 27332
rect 50508 27280 50554 27332
rect 50554 27280 50564 27332
rect 50588 27280 50618 27332
rect 50618 27280 50644 27332
rect 50348 27278 50404 27280
rect 50428 27278 50484 27280
rect 50508 27278 50564 27280
rect 50588 27278 50644 27280
rect 50348 26000 50404 26002
rect 50428 26000 50484 26002
rect 50508 26000 50564 26002
rect 50588 26000 50644 26002
rect 50348 25948 50374 26000
rect 50374 25948 50404 26000
rect 50428 25948 50438 26000
rect 50438 25948 50484 26000
rect 50508 25948 50554 26000
rect 50554 25948 50564 26000
rect 50588 25948 50618 26000
rect 50618 25948 50644 26000
rect 50348 25946 50404 25948
rect 50428 25946 50484 25948
rect 50508 25946 50564 25948
rect 50588 25946 50644 25948
rect 50348 24668 50404 24670
rect 50428 24668 50484 24670
rect 50508 24668 50564 24670
rect 50588 24668 50644 24670
rect 50348 24616 50374 24668
rect 50374 24616 50404 24668
rect 50428 24616 50438 24668
rect 50438 24616 50484 24668
rect 50508 24616 50554 24668
rect 50554 24616 50564 24668
rect 50588 24616 50618 24668
rect 50618 24616 50644 24668
rect 50348 24614 50404 24616
rect 50428 24614 50484 24616
rect 50508 24614 50564 24616
rect 50588 24614 50644 24616
rect 50348 23336 50404 23338
rect 50428 23336 50484 23338
rect 50508 23336 50564 23338
rect 50588 23336 50644 23338
rect 50348 23284 50374 23336
rect 50374 23284 50404 23336
rect 50428 23284 50438 23336
rect 50438 23284 50484 23336
rect 50508 23284 50554 23336
rect 50554 23284 50564 23336
rect 50588 23284 50618 23336
rect 50618 23284 50644 23336
rect 50348 23282 50404 23284
rect 50428 23282 50484 23284
rect 50508 23282 50564 23284
rect 50588 23282 50644 23284
rect 50348 22004 50404 22006
rect 50428 22004 50484 22006
rect 50508 22004 50564 22006
rect 50588 22004 50644 22006
rect 50348 21952 50374 22004
rect 50374 21952 50404 22004
rect 50428 21952 50438 22004
rect 50438 21952 50484 22004
rect 50508 21952 50554 22004
rect 50554 21952 50564 22004
rect 50588 21952 50618 22004
rect 50618 21952 50644 22004
rect 50348 21950 50404 21952
rect 50428 21950 50484 21952
rect 50508 21950 50564 21952
rect 50588 21950 50644 21952
rect 50348 20672 50404 20674
rect 50428 20672 50484 20674
rect 50508 20672 50564 20674
rect 50588 20672 50644 20674
rect 50348 20620 50374 20672
rect 50374 20620 50404 20672
rect 50428 20620 50438 20672
rect 50438 20620 50484 20672
rect 50508 20620 50554 20672
rect 50554 20620 50564 20672
rect 50588 20620 50618 20672
rect 50618 20620 50644 20672
rect 50348 20618 50404 20620
rect 50428 20618 50484 20620
rect 50508 20618 50564 20620
rect 50588 20618 50644 20620
rect 50348 19340 50404 19342
rect 50428 19340 50484 19342
rect 50508 19340 50564 19342
rect 50588 19340 50644 19342
rect 50348 19288 50374 19340
rect 50374 19288 50404 19340
rect 50428 19288 50438 19340
rect 50438 19288 50484 19340
rect 50508 19288 50554 19340
rect 50554 19288 50564 19340
rect 50588 19288 50618 19340
rect 50618 19288 50644 19340
rect 50348 19286 50404 19288
rect 50428 19286 50484 19288
rect 50508 19286 50564 19288
rect 50588 19286 50644 19288
rect 50348 18008 50404 18010
rect 50428 18008 50484 18010
rect 50508 18008 50564 18010
rect 50588 18008 50644 18010
rect 50348 17956 50374 18008
rect 50374 17956 50404 18008
rect 50428 17956 50438 18008
rect 50438 17956 50484 18008
rect 50508 17956 50554 18008
rect 50554 17956 50564 18008
rect 50588 17956 50618 18008
rect 50618 17956 50644 18008
rect 50348 17954 50404 17956
rect 50428 17954 50484 17956
rect 50508 17954 50564 17956
rect 50588 17954 50644 17956
rect 50348 16676 50404 16678
rect 50428 16676 50484 16678
rect 50508 16676 50564 16678
rect 50588 16676 50644 16678
rect 50348 16624 50374 16676
rect 50374 16624 50404 16676
rect 50428 16624 50438 16676
rect 50438 16624 50484 16676
rect 50508 16624 50554 16676
rect 50554 16624 50564 16676
rect 50588 16624 50618 16676
rect 50618 16624 50644 16676
rect 50348 16622 50404 16624
rect 50428 16622 50484 16624
rect 50508 16622 50564 16624
rect 50588 16622 50644 16624
rect 50348 15344 50404 15346
rect 50428 15344 50484 15346
rect 50508 15344 50564 15346
rect 50588 15344 50644 15346
rect 50348 15292 50374 15344
rect 50374 15292 50404 15344
rect 50428 15292 50438 15344
rect 50438 15292 50484 15344
rect 50508 15292 50554 15344
rect 50554 15292 50564 15344
rect 50588 15292 50618 15344
rect 50618 15292 50644 15344
rect 50348 15290 50404 15292
rect 50428 15290 50484 15292
rect 50508 15290 50564 15292
rect 50588 15290 50644 15292
rect 50348 14012 50404 14014
rect 50428 14012 50484 14014
rect 50508 14012 50564 14014
rect 50588 14012 50644 14014
rect 50348 13960 50374 14012
rect 50374 13960 50404 14012
rect 50428 13960 50438 14012
rect 50438 13960 50484 14012
rect 50508 13960 50554 14012
rect 50554 13960 50564 14012
rect 50588 13960 50618 14012
rect 50618 13960 50644 14012
rect 50348 13958 50404 13960
rect 50428 13958 50484 13960
rect 50508 13958 50564 13960
rect 50588 13958 50644 13960
rect 50348 12680 50404 12682
rect 50428 12680 50484 12682
rect 50508 12680 50564 12682
rect 50588 12680 50644 12682
rect 50348 12628 50374 12680
rect 50374 12628 50404 12680
rect 50428 12628 50438 12680
rect 50438 12628 50484 12680
rect 50508 12628 50554 12680
rect 50554 12628 50564 12680
rect 50588 12628 50618 12680
rect 50618 12628 50644 12680
rect 50348 12626 50404 12628
rect 50428 12626 50484 12628
rect 50508 12626 50564 12628
rect 50588 12626 50644 12628
rect 50348 11348 50404 11350
rect 50428 11348 50484 11350
rect 50508 11348 50564 11350
rect 50588 11348 50644 11350
rect 50348 11296 50374 11348
rect 50374 11296 50404 11348
rect 50428 11296 50438 11348
rect 50438 11296 50484 11348
rect 50508 11296 50554 11348
rect 50554 11296 50564 11348
rect 50588 11296 50618 11348
rect 50618 11296 50644 11348
rect 50348 11294 50404 11296
rect 50428 11294 50484 11296
rect 50508 11294 50564 11296
rect 50588 11294 50644 11296
rect 50348 10016 50404 10018
rect 50428 10016 50484 10018
rect 50508 10016 50564 10018
rect 50588 10016 50644 10018
rect 50348 9964 50374 10016
rect 50374 9964 50404 10016
rect 50428 9964 50438 10016
rect 50438 9964 50484 10016
rect 50508 9964 50554 10016
rect 50554 9964 50564 10016
rect 50588 9964 50618 10016
rect 50618 9964 50644 10016
rect 50348 9962 50404 9964
rect 50428 9962 50484 9964
rect 50508 9962 50564 9964
rect 50588 9962 50644 9964
rect 50348 8684 50404 8686
rect 50428 8684 50484 8686
rect 50508 8684 50564 8686
rect 50588 8684 50644 8686
rect 50348 8632 50374 8684
rect 50374 8632 50404 8684
rect 50428 8632 50438 8684
rect 50438 8632 50484 8684
rect 50508 8632 50554 8684
rect 50554 8632 50564 8684
rect 50588 8632 50618 8684
rect 50618 8632 50644 8684
rect 50348 8630 50404 8632
rect 50428 8630 50484 8632
rect 50508 8630 50564 8632
rect 50588 8630 50644 8632
rect 50348 7352 50404 7354
rect 50428 7352 50484 7354
rect 50508 7352 50564 7354
rect 50588 7352 50644 7354
rect 50348 7300 50374 7352
rect 50374 7300 50404 7352
rect 50428 7300 50438 7352
rect 50438 7300 50484 7352
rect 50508 7300 50554 7352
rect 50554 7300 50564 7352
rect 50588 7300 50618 7352
rect 50618 7300 50644 7352
rect 50348 7298 50404 7300
rect 50428 7298 50484 7300
rect 50508 7298 50564 7300
rect 50588 7298 50644 7300
rect 50348 6020 50404 6022
rect 50428 6020 50484 6022
rect 50508 6020 50564 6022
rect 50588 6020 50644 6022
rect 50348 5968 50374 6020
rect 50374 5968 50404 6020
rect 50428 5968 50438 6020
rect 50438 5968 50484 6020
rect 50508 5968 50554 6020
rect 50554 5968 50564 6020
rect 50588 5968 50618 6020
rect 50618 5968 50644 6020
rect 50348 5966 50404 5968
rect 50428 5966 50484 5968
rect 50508 5966 50564 5968
rect 50588 5966 50644 5968
rect 50348 4688 50404 4690
rect 50428 4688 50484 4690
rect 50508 4688 50564 4690
rect 50588 4688 50644 4690
rect 50348 4636 50374 4688
rect 50374 4636 50404 4688
rect 50428 4636 50438 4688
rect 50438 4636 50484 4688
rect 50508 4636 50554 4688
rect 50554 4636 50564 4688
rect 50588 4636 50618 4688
rect 50618 4636 50644 4688
rect 50348 4634 50404 4636
rect 50428 4634 50484 4636
rect 50508 4634 50564 4636
rect 50588 4634 50644 4636
rect 50348 3356 50404 3358
rect 50428 3356 50484 3358
rect 50508 3356 50564 3358
rect 50588 3356 50644 3358
rect 50348 3304 50374 3356
rect 50374 3304 50404 3356
rect 50428 3304 50438 3356
rect 50438 3304 50484 3356
rect 50508 3304 50554 3356
rect 50554 3304 50564 3356
rect 50588 3304 50618 3356
rect 50618 3304 50644 3356
rect 50348 3302 50404 3304
rect 50428 3302 50484 3304
rect 50508 3302 50564 3304
rect 50588 3302 50644 3304
<< metal3 >>
rect 4256 57308 4576 57309
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 57243 4576 57244
rect 34976 57308 35296 57309
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 57243 35296 57244
rect 19616 56642 19936 56643
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 56577 19936 56578
rect 50336 56642 50656 56643
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 56577 50656 56578
rect 4256 55976 4576 55977
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 55911 4576 55912
rect 34976 55976 35296 55977
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 55911 35296 55912
rect 19616 55310 19936 55311
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 55245 19936 55246
rect 50336 55310 50656 55311
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 55245 50656 55246
rect 4256 54644 4576 54645
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 54579 4576 54580
rect 34976 54644 35296 54645
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 54579 35296 54580
rect 19616 53978 19936 53979
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 53913 19936 53914
rect 50336 53978 50656 53979
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 53913 50656 53914
rect 4256 53312 4576 53313
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 53247 4576 53248
rect 34976 53312 35296 53313
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 53247 35296 53248
rect 19616 52646 19936 52647
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 52581 19936 52582
rect 50336 52646 50656 52647
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 52581 50656 52582
rect 4256 51980 4576 51981
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 51915 4576 51916
rect 34976 51980 35296 51981
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 51915 35296 51916
rect 19616 51314 19936 51315
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 51249 19936 51250
rect 50336 51314 50656 51315
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 51249 50656 51250
rect 4256 50648 4576 50649
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 50583 4576 50584
rect 34976 50648 35296 50649
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 50583 35296 50584
rect 19616 49982 19936 49983
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 49917 19936 49918
rect 50336 49982 50656 49983
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 49917 50656 49918
rect 4256 49316 4576 49317
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 49251 4576 49252
rect 34976 49316 35296 49317
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 49251 35296 49252
rect 19616 48650 19936 48651
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 48585 19936 48586
rect 50336 48650 50656 48651
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 48585 50656 48586
rect 4256 47984 4576 47985
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 47919 4576 47920
rect 34976 47984 35296 47985
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 47919 35296 47920
rect 19616 47318 19936 47319
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 47253 19936 47254
rect 50336 47318 50656 47319
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 47253 50656 47254
rect 4256 46652 4576 46653
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 46587 4576 46588
rect 34976 46652 35296 46653
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 46587 35296 46588
rect 19616 45986 19936 45987
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 45921 19936 45922
rect 50336 45986 50656 45987
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 45921 50656 45922
rect 4256 45320 4576 45321
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 45255 4576 45256
rect 34976 45320 35296 45321
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 45255 35296 45256
rect 19616 44654 19936 44655
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 44589 19936 44590
rect 50336 44654 50656 44655
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 44589 50656 44590
rect 4256 43988 4576 43989
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 43923 4576 43924
rect 34976 43988 35296 43989
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 43923 35296 43924
rect 19616 43322 19936 43323
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 43257 19936 43258
rect 50336 43322 50656 43323
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 43257 50656 43258
rect 4256 42656 4576 42657
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 42591 4576 42592
rect 34976 42656 35296 42657
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 42591 35296 42592
rect 19616 41990 19936 41991
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 41925 19936 41926
rect 50336 41990 50656 41991
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 41925 50656 41926
rect 4256 41324 4576 41325
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 41259 4576 41260
rect 34976 41324 35296 41325
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 41259 35296 41260
rect 19616 40658 19936 40659
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 40593 19936 40594
rect 50336 40658 50656 40659
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 40593 50656 40594
rect 4256 39992 4576 39993
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 39927 4576 39928
rect 34976 39992 35296 39993
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 39927 35296 39928
rect 19616 39326 19936 39327
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 39261 19936 39262
rect 50336 39326 50656 39327
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 39261 50656 39262
rect 4256 38660 4576 38661
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 38595 4576 38596
rect 34976 38660 35296 38661
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 38595 35296 38596
rect 19616 37994 19936 37995
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 37929 19936 37930
rect 50336 37994 50656 37995
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 37929 50656 37930
rect 4256 37328 4576 37329
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 37263 4576 37264
rect 34976 37328 35296 37329
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 37263 35296 37264
rect 19616 36662 19936 36663
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 36597 19936 36598
rect 50336 36662 50656 36663
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 36597 50656 36598
rect 4256 35996 4576 35997
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 35931 4576 35932
rect 34976 35996 35296 35997
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 35931 35296 35932
rect 19616 35330 19936 35331
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 35265 19936 35266
rect 50336 35330 50656 35331
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 35265 50656 35266
rect 4256 34664 4576 34665
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 34599 4576 34600
rect 34976 34664 35296 34665
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 34599 35296 34600
rect 19616 33998 19936 33999
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 33933 19936 33934
rect 50336 33998 50656 33999
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 33933 50656 33934
rect 4256 33332 4576 33333
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 33267 4576 33268
rect 34976 33332 35296 33333
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 33267 35296 33268
rect 19616 32666 19936 32667
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 32601 19936 32602
rect 50336 32666 50656 32667
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 32601 50656 32602
rect 4256 32000 4576 32001
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 31935 4576 31936
rect 34976 32000 35296 32001
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 31935 35296 31936
rect 19616 31334 19936 31335
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 31269 19936 31270
rect 50336 31334 50656 31335
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 31269 50656 31270
rect 4256 30668 4576 30669
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 30603 4576 30604
rect 34976 30668 35296 30669
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 30603 35296 30604
rect 19616 30002 19936 30003
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 29937 19936 29938
rect 50336 30002 50656 30003
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 29937 50656 29938
rect 4256 29336 4576 29337
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 29271 4576 29272
rect 34976 29336 35296 29337
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 29271 35296 29272
rect 19616 28670 19936 28671
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 28605 19936 28606
rect 50336 28670 50656 28671
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 28605 50656 28606
rect 4256 28004 4576 28005
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 27939 4576 27940
rect 34976 28004 35296 28005
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 27939 35296 27940
rect 19616 27338 19936 27339
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 27273 19936 27274
rect 50336 27338 50656 27339
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 27273 50656 27274
rect 4256 26672 4576 26673
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 26607 4576 26608
rect 34976 26672 35296 26673
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 26607 35296 26608
rect 19616 26006 19936 26007
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 25941 19936 25942
rect 50336 26006 50656 26007
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 25941 50656 25942
rect 4256 25340 4576 25341
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 25275 4576 25276
rect 34976 25340 35296 25341
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 25275 35296 25276
rect 19616 24674 19936 24675
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 24609 19936 24610
rect 50336 24674 50656 24675
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 24609 50656 24610
rect 4256 24008 4576 24009
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 23943 4576 23944
rect 34976 24008 35296 24009
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 23943 35296 23944
rect 19616 23342 19936 23343
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 23277 19936 23278
rect 50336 23342 50656 23343
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 23277 50656 23278
rect 4256 22676 4576 22677
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 22611 4576 22612
rect 34976 22676 35296 22677
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 22611 35296 22612
rect 19616 22010 19936 22011
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 21945 19936 21946
rect 50336 22010 50656 22011
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 21945 50656 21946
rect 4256 21344 4576 21345
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 21279 4576 21280
rect 34976 21344 35296 21345
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 21279 35296 21280
rect 19616 20678 19936 20679
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 20613 19936 20614
rect 50336 20678 50656 20679
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 20613 50656 20614
rect 4256 20012 4576 20013
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 19947 4576 19948
rect 34976 20012 35296 20013
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 19947 35296 19948
rect 19616 19346 19936 19347
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 19281 19936 19282
rect 50336 19346 50656 19347
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 19281 50656 19282
rect 4256 18680 4576 18681
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 18615 4576 18616
rect 34976 18680 35296 18681
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 18615 35296 18616
rect 19616 18014 19936 18015
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 17949 19936 17950
rect 50336 18014 50656 18015
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 17949 50656 17950
rect 4256 17348 4576 17349
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 17283 4576 17284
rect 34976 17348 35296 17349
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 17283 35296 17284
rect 19616 16682 19936 16683
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 16617 19936 16618
rect 50336 16682 50656 16683
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 16617 50656 16618
rect 4256 16016 4576 16017
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 15951 4576 15952
rect 34976 16016 35296 16017
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 15951 35296 15952
rect 19616 15350 19936 15351
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 15285 19936 15286
rect 50336 15350 50656 15351
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 15285 50656 15286
rect 4256 14684 4576 14685
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 14619 4576 14620
rect 34976 14684 35296 14685
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 14619 35296 14620
rect 7599 14460 7665 14463
rect 8175 14460 8241 14463
rect 7599 14458 8241 14460
rect 7599 14402 7604 14458
rect 7660 14402 8180 14458
rect 8236 14402 8241 14458
rect 7599 14400 8241 14402
rect 7599 14397 7665 14400
rect 8175 14397 8241 14400
rect 19616 14018 19936 14019
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 13953 19936 13954
rect 50336 14018 50656 14019
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 13953 50656 13954
rect 4256 13352 4576 13353
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 13287 4576 13288
rect 34976 13352 35296 13353
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 13287 35296 13288
rect 19616 12686 19936 12687
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 12621 19936 12622
rect 50336 12686 50656 12687
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 12621 50656 12622
rect 4256 12020 4576 12021
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 11955 4576 11956
rect 34976 12020 35296 12021
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 11955 35296 11956
rect 19616 11354 19936 11355
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 11289 19936 11290
rect 50336 11354 50656 11355
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 11289 50656 11290
rect 4256 10688 4576 10689
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 10623 4576 10624
rect 34976 10688 35296 10689
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 10623 35296 10624
rect 19616 10022 19936 10023
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 9957 19936 9958
rect 50336 10022 50656 10023
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 9957 50656 9958
rect 4256 9356 4576 9357
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 9291 4576 9292
rect 34976 9356 35296 9357
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 9291 35296 9292
rect 7935 8836 8001 8839
rect 8271 8836 8337 8839
rect 7935 8834 8337 8836
rect 7935 8778 7940 8834
rect 7996 8778 8276 8834
rect 8332 8778 8337 8834
rect 7935 8776 8337 8778
rect 7935 8773 8001 8776
rect 8271 8773 8337 8776
rect 19616 8690 19936 8691
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 8625 19936 8626
rect 50336 8690 50656 8691
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 8625 50656 8626
rect 4256 8024 4576 8025
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 7959 4576 7960
rect 34976 8024 35296 8025
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 7959 35296 7960
rect 7935 7948 8001 7951
rect 12207 7948 12273 7951
rect 7935 7946 12273 7948
rect 7935 7890 7940 7946
rect 7996 7890 12212 7946
rect 12268 7890 12273 7946
rect 7935 7888 12273 7890
rect 7935 7885 8001 7888
rect 12207 7885 12273 7888
rect 4911 7800 4977 7803
rect 8559 7800 8625 7803
rect 4911 7798 8625 7800
rect 4911 7742 4916 7798
rect 4972 7742 8564 7798
rect 8620 7742 8625 7798
rect 4911 7740 8625 7742
rect 4911 7737 4977 7740
rect 8559 7737 8625 7740
rect 8223 7652 8289 7655
rect 9519 7652 9585 7655
rect 8223 7650 9585 7652
rect 8223 7594 8228 7650
rect 8284 7594 9524 7650
rect 9580 7594 9585 7650
rect 8223 7592 9585 7594
rect 8223 7589 8289 7592
rect 9519 7589 9585 7592
rect 19616 7358 19936 7359
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 7293 19936 7294
rect 50336 7358 50656 7359
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 7293 50656 7294
rect 4256 6692 4576 6693
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 6627 4576 6628
rect 34976 6692 35296 6693
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 6627 35296 6628
rect 19616 6026 19936 6027
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 5961 19936 5962
rect 50336 6026 50656 6027
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 5961 50656 5962
rect 4256 5360 4576 5361
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 5295 4576 5296
rect 34976 5360 35296 5361
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 5295 35296 5296
rect 19616 4694 19936 4695
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 4629 19936 4630
rect 50336 4694 50656 4695
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 4629 50656 4630
rect 4256 4028 4576 4029
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 3963 4576 3964
rect 34976 4028 35296 4029
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 3963 35296 3964
rect 19616 3362 19936 3363
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 19616 3297 19936 3298
rect 50336 3362 50656 3363
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 50336 3297 50656 3298
rect 35919 3212 35985 3215
rect 35394 3210 35985 3212
rect 35394 3154 35924 3210
rect 35980 3154 35985 3210
rect 35394 3152 35985 3154
rect 34479 2916 34545 2919
rect 35247 2916 35313 2919
rect 34479 2914 35313 2916
rect 34479 2858 34484 2914
rect 34540 2858 35252 2914
rect 35308 2858 35313 2914
rect 34479 2856 35313 2858
rect 34479 2853 34545 2856
rect 35247 2853 35313 2856
rect 4256 2696 4576 2697
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4256 2631 4576 2632
rect 34976 2696 35296 2697
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 34976 2631 35296 2632
rect 35151 2472 35217 2475
rect 35394 2472 35454 3152
rect 35919 3149 35985 3152
rect 35151 2470 35454 2472
rect 35151 2414 35156 2470
rect 35212 2414 35454 2470
rect 35151 2412 35454 2414
rect 35151 2409 35217 2412
<< via3 >>
rect 4264 57304 4328 57308
rect 4264 57248 4268 57304
rect 4268 57248 4324 57304
rect 4324 57248 4328 57304
rect 4264 57244 4328 57248
rect 4344 57304 4408 57308
rect 4344 57248 4348 57304
rect 4348 57248 4404 57304
rect 4404 57248 4408 57304
rect 4344 57244 4408 57248
rect 4424 57304 4488 57308
rect 4424 57248 4428 57304
rect 4428 57248 4484 57304
rect 4484 57248 4488 57304
rect 4424 57244 4488 57248
rect 4504 57304 4568 57308
rect 4504 57248 4508 57304
rect 4508 57248 4564 57304
rect 4564 57248 4568 57304
rect 4504 57244 4568 57248
rect 34984 57304 35048 57308
rect 34984 57248 34988 57304
rect 34988 57248 35044 57304
rect 35044 57248 35048 57304
rect 34984 57244 35048 57248
rect 35064 57304 35128 57308
rect 35064 57248 35068 57304
rect 35068 57248 35124 57304
rect 35124 57248 35128 57304
rect 35064 57244 35128 57248
rect 35144 57304 35208 57308
rect 35144 57248 35148 57304
rect 35148 57248 35204 57304
rect 35204 57248 35208 57304
rect 35144 57244 35208 57248
rect 35224 57304 35288 57308
rect 35224 57248 35228 57304
rect 35228 57248 35284 57304
rect 35284 57248 35288 57304
rect 35224 57244 35288 57248
rect 19624 56638 19688 56642
rect 19624 56582 19628 56638
rect 19628 56582 19684 56638
rect 19684 56582 19688 56638
rect 19624 56578 19688 56582
rect 19704 56638 19768 56642
rect 19704 56582 19708 56638
rect 19708 56582 19764 56638
rect 19764 56582 19768 56638
rect 19704 56578 19768 56582
rect 19784 56638 19848 56642
rect 19784 56582 19788 56638
rect 19788 56582 19844 56638
rect 19844 56582 19848 56638
rect 19784 56578 19848 56582
rect 19864 56638 19928 56642
rect 19864 56582 19868 56638
rect 19868 56582 19924 56638
rect 19924 56582 19928 56638
rect 19864 56578 19928 56582
rect 50344 56638 50408 56642
rect 50344 56582 50348 56638
rect 50348 56582 50404 56638
rect 50404 56582 50408 56638
rect 50344 56578 50408 56582
rect 50424 56638 50488 56642
rect 50424 56582 50428 56638
rect 50428 56582 50484 56638
rect 50484 56582 50488 56638
rect 50424 56578 50488 56582
rect 50504 56638 50568 56642
rect 50504 56582 50508 56638
rect 50508 56582 50564 56638
rect 50564 56582 50568 56638
rect 50504 56578 50568 56582
rect 50584 56638 50648 56642
rect 50584 56582 50588 56638
rect 50588 56582 50644 56638
rect 50644 56582 50648 56638
rect 50584 56578 50648 56582
rect 4264 55972 4328 55976
rect 4264 55916 4268 55972
rect 4268 55916 4324 55972
rect 4324 55916 4328 55972
rect 4264 55912 4328 55916
rect 4344 55972 4408 55976
rect 4344 55916 4348 55972
rect 4348 55916 4404 55972
rect 4404 55916 4408 55972
rect 4344 55912 4408 55916
rect 4424 55972 4488 55976
rect 4424 55916 4428 55972
rect 4428 55916 4484 55972
rect 4484 55916 4488 55972
rect 4424 55912 4488 55916
rect 4504 55972 4568 55976
rect 4504 55916 4508 55972
rect 4508 55916 4564 55972
rect 4564 55916 4568 55972
rect 4504 55912 4568 55916
rect 34984 55972 35048 55976
rect 34984 55916 34988 55972
rect 34988 55916 35044 55972
rect 35044 55916 35048 55972
rect 34984 55912 35048 55916
rect 35064 55972 35128 55976
rect 35064 55916 35068 55972
rect 35068 55916 35124 55972
rect 35124 55916 35128 55972
rect 35064 55912 35128 55916
rect 35144 55972 35208 55976
rect 35144 55916 35148 55972
rect 35148 55916 35204 55972
rect 35204 55916 35208 55972
rect 35144 55912 35208 55916
rect 35224 55972 35288 55976
rect 35224 55916 35228 55972
rect 35228 55916 35284 55972
rect 35284 55916 35288 55972
rect 35224 55912 35288 55916
rect 19624 55306 19688 55310
rect 19624 55250 19628 55306
rect 19628 55250 19684 55306
rect 19684 55250 19688 55306
rect 19624 55246 19688 55250
rect 19704 55306 19768 55310
rect 19704 55250 19708 55306
rect 19708 55250 19764 55306
rect 19764 55250 19768 55306
rect 19704 55246 19768 55250
rect 19784 55306 19848 55310
rect 19784 55250 19788 55306
rect 19788 55250 19844 55306
rect 19844 55250 19848 55306
rect 19784 55246 19848 55250
rect 19864 55306 19928 55310
rect 19864 55250 19868 55306
rect 19868 55250 19924 55306
rect 19924 55250 19928 55306
rect 19864 55246 19928 55250
rect 50344 55306 50408 55310
rect 50344 55250 50348 55306
rect 50348 55250 50404 55306
rect 50404 55250 50408 55306
rect 50344 55246 50408 55250
rect 50424 55306 50488 55310
rect 50424 55250 50428 55306
rect 50428 55250 50484 55306
rect 50484 55250 50488 55306
rect 50424 55246 50488 55250
rect 50504 55306 50568 55310
rect 50504 55250 50508 55306
rect 50508 55250 50564 55306
rect 50564 55250 50568 55306
rect 50504 55246 50568 55250
rect 50584 55306 50648 55310
rect 50584 55250 50588 55306
rect 50588 55250 50644 55306
rect 50644 55250 50648 55306
rect 50584 55246 50648 55250
rect 4264 54640 4328 54644
rect 4264 54584 4268 54640
rect 4268 54584 4324 54640
rect 4324 54584 4328 54640
rect 4264 54580 4328 54584
rect 4344 54640 4408 54644
rect 4344 54584 4348 54640
rect 4348 54584 4404 54640
rect 4404 54584 4408 54640
rect 4344 54580 4408 54584
rect 4424 54640 4488 54644
rect 4424 54584 4428 54640
rect 4428 54584 4484 54640
rect 4484 54584 4488 54640
rect 4424 54580 4488 54584
rect 4504 54640 4568 54644
rect 4504 54584 4508 54640
rect 4508 54584 4564 54640
rect 4564 54584 4568 54640
rect 4504 54580 4568 54584
rect 34984 54640 35048 54644
rect 34984 54584 34988 54640
rect 34988 54584 35044 54640
rect 35044 54584 35048 54640
rect 34984 54580 35048 54584
rect 35064 54640 35128 54644
rect 35064 54584 35068 54640
rect 35068 54584 35124 54640
rect 35124 54584 35128 54640
rect 35064 54580 35128 54584
rect 35144 54640 35208 54644
rect 35144 54584 35148 54640
rect 35148 54584 35204 54640
rect 35204 54584 35208 54640
rect 35144 54580 35208 54584
rect 35224 54640 35288 54644
rect 35224 54584 35228 54640
rect 35228 54584 35284 54640
rect 35284 54584 35288 54640
rect 35224 54580 35288 54584
rect 19624 53974 19688 53978
rect 19624 53918 19628 53974
rect 19628 53918 19684 53974
rect 19684 53918 19688 53974
rect 19624 53914 19688 53918
rect 19704 53974 19768 53978
rect 19704 53918 19708 53974
rect 19708 53918 19764 53974
rect 19764 53918 19768 53974
rect 19704 53914 19768 53918
rect 19784 53974 19848 53978
rect 19784 53918 19788 53974
rect 19788 53918 19844 53974
rect 19844 53918 19848 53974
rect 19784 53914 19848 53918
rect 19864 53974 19928 53978
rect 19864 53918 19868 53974
rect 19868 53918 19924 53974
rect 19924 53918 19928 53974
rect 19864 53914 19928 53918
rect 50344 53974 50408 53978
rect 50344 53918 50348 53974
rect 50348 53918 50404 53974
rect 50404 53918 50408 53974
rect 50344 53914 50408 53918
rect 50424 53974 50488 53978
rect 50424 53918 50428 53974
rect 50428 53918 50484 53974
rect 50484 53918 50488 53974
rect 50424 53914 50488 53918
rect 50504 53974 50568 53978
rect 50504 53918 50508 53974
rect 50508 53918 50564 53974
rect 50564 53918 50568 53974
rect 50504 53914 50568 53918
rect 50584 53974 50648 53978
rect 50584 53918 50588 53974
rect 50588 53918 50644 53974
rect 50644 53918 50648 53974
rect 50584 53914 50648 53918
rect 4264 53308 4328 53312
rect 4264 53252 4268 53308
rect 4268 53252 4324 53308
rect 4324 53252 4328 53308
rect 4264 53248 4328 53252
rect 4344 53308 4408 53312
rect 4344 53252 4348 53308
rect 4348 53252 4404 53308
rect 4404 53252 4408 53308
rect 4344 53248 4408 53252
rect 4424 53308 4488 53312
rect 4424 53252 4428 53308
rect 4428 53252 4484 53308
rect 4484 53252 4488 53308
rect 4424 53248 4488 53252
rect 4504 53308 4568 53312
rect 4504 53252 4508 53308
rect 4508 53252 4564 53308
rect 4564 53252 4568 53308
rect 4504 53248 4568 53252
rect 34984 53308 35048 53312
rect 34984 53252 34988 53308
rect 34988 53252 35044 53308
rect 35044 53252 35048 53308
rect 34984 53248 35048 53252
rect 35064 53308 35128 53312
rect 35064 53252 35068 53308
rect 35068 53252 35124 53308
rect 35124 53252 35128 53308
rect 35064 53248 35128 53252
rect 35144 53308 35208 53312
rect 35144 53252 35148 53308
rect 35148 53252 35204 53308
rect 35204 53252 35208 53308
rect 35144 53248 35208 53252
rect 35224 53308 35288 53312
rect 35224 53252 35228 53308
rect 35228 53252 35284 53308
rect 35284 53252 35288 53308
rect 35224 53248 35288 53252
rect 19624 52642 19688 52646
rect 19624 52586 19628 52642
rect 19628 52586 19684 52642
rect 19684 52586 19688 52642
rect 19624 52582 19688 52586
rect 19704 52642 19768 52646
rect 19704 52586 19708 52642
rect 19708 52586 19764 52642
rect 19764 52586 19768 52642
rect 19704 52582 19768 52586
rect 19784 52642 19848 52646
rect 19784 52586 19788 52642
rect 19788 52586 19844 52642
rect 19844 52586 19848 52642
rect 19784 52582 19848 52586
rect 19864 52642 19928 52646
rect 19864 52586 19868 52642
rect 19868 52586 19924 52642
rect 19924 52586 19928 52642
rect 19864 52582 19928 52586
rect 50344 52642 50408 52646
rect 50344 52586 50348 52642
rect 50348 52586 50404 52642
rect 50404 52586 50408 52642
rect 50344 52582 50408 52586
rect 50424 52642 50488 52646
rect 50424 52586 50428 52642
rect 50428 52586 50484 52642
rect 50484 52586 50488 52642
rect 50424 52582 50488 52586
rect 50504 52642 50568 52646
rect 50504 52586 50508 52642
rect 50508 52586 50564 52642
rect 50564 52586 50568 52642
rect 50504 52582 50568 52586
rect 50584 52642 50648 52646
rect 50584 52586 50588 52642
rect 50588 52586 50644 52642
rect 50644 52586 50648 52642
rect 50584 52582 50648 52586
rect 4264 51976 4328 51980
rect 4264 51920 4268 51976
rect 4268 51920 4324 51976
rect 4324 51920 4328 51976
rect 4264 51916 4328 51920
rect 4344 51976 4408 51980
rect 4344 51920 4348 51976
rect 4348 51920 4404 51976
rect 4404 51920 4408 51976
rect 4344 51916 4408 51920
rect 4424 51976 4488 51980
rect 4424 51920 4428 51976
rect 4428 51920 4484 51976
rect 4484 51920 4488 51976
rect 4424 51916 4488 51920
rect 4504 51976 4568 51980
rect 4504 51920 4508 51976
rect 4508 51920 4564 51976
rect 4564 51920 4568 51976
rect 4504 51916 4568 51920
rect 34984 51976 35048 51980
rect 34984 51920 34988 51976
rect 34988 51920 35044 51976
rect 35044 51920 35048 51976
rect 34984 51916 35048 51920
rect 35064 51976 35128 51980
rect 35064 51920 35068 51976
rect 35068 51920 35124 51976
rect 35124 51920 35128 51976
rect 35064 51916 35128 51920
rect 35144 51976 35208 51980
rect 35144 51920 35148 51976
rect 35148 51920 35204 51976
rect 35204 51920 35208 51976
rect 35144 51916 35208 51920
rect 35224 51976 35288 51980
rect 35224 51920 35228 51976
rect 35228 51920 35284 51976
rect 35284 51920 35288 51976
rect 35224 51916 35288 51920
rect 19624 51310 19688 51314
rect 19624 51254 19628 51310
rect 19628 51254 19684 51310
rect 19684 51254 19688 51310
rect 19624 51250 19688 51254
rect 19704 51310 19768 51314
rect 19704 51254 19708 51310
rect 19708 51254 19764 51310
rect 19764 51254 19768 51310
rect 19704 51250 19768 51254
rect 19784 51310 19848 51314
rect 19784 51254 19788 51310
rect 19788 51254 19844 51310
rect 19844 51254 19848 51310
rect 19784 51250 19848 51254
rect 19864 51310 19928 51314
rect 19864 51254 19868 51310
rect 19868 51254 19924 51310
rect 19924 51254 19928 51310
rect 19864 51250 19928 51254
rect 50344 51310 50408 51314
rect 50344 51254 50348 51310
rect 50348 51254 50404 51310
rect 50404 51254 50408 51310
rect 50344 51250 50408 51254
rect 50424 51310 50488 51314
rect 50424 51254 50428 51310
rect 50428 51254 50484 51310
rect 50484 51254 50488 51310
rect 50424 51250 50488 51254
rect 50504 51310 50568 51314
rect 50504 51254 50508 51310
rect 50508 51254 50564 51310
rect 50564 51254 50568 51310
rect 50504 51250 50568 51254
rect 50584 51310 50648 51314
rect 50584 51254 50588 51310
rect 50588 51254 50644 51310
rect 50644 51254 50648 51310
rect 50584 51250 50648 51254
rect 4264 50644 4328 50648
rect 4264 50588 4268 50644
rect 4268 50588 4324 50644
rect 4324 50588 4328 50644
rect 4264 50584 4328 50588
rect 4344 50644 4408 50648
rect 4344 50588 4348 50644
rect 4348 50588 4404 50644
rect 4404 50588 4408 50644
rect 4344 50584 4408 50588
rect 4424 50644 4488 50648
rect 4424 50588 4428 50644
rect 4428 50588 4484 50644
rect 4484 50588 4488 50644
rect 4424 50584 4488 50588
rect 4504 50644 4568 50648
rect 4504 50588 4508 50644
rect 4508 50588 4564 50644
rect 4564 50588 4568 50644
rect 4504 50584 4568 50588
rect 34984 50644 35048 50648
rect 34984 50588 34988 50644
rect 34988 50588 35044 50644
rect 35044 50588 35048 50644
rect 34984 50584 35048 50588
rect 35064 50644 35128 50648
rect 35064 50588 35068 50644
rect 35068 50588 35124 50644
rect 35124 50588 35128 50644
rect 35064 50584 35128 50588
rect 35144 50644 35208 50648
rect 35144 50588 35148 50644
rect 35148 50588 35204 50644
rect 35204 50588 35208 50644
rect 35144 50584 35208 50588
rect 35224 50644 35288 50648
rect 35224 50588 35228 50644
rect 35228 50588 35284 50644
rect 35284 50588 35288 50644
rect 35224 50584 35288 50588
rect 19624 49978 19688 49982
rect 19624 49922 19628 49978
rect 19628 49922 19684 49978
rect 19684 49922 19688 49978
rect 19624 49918 19688 49922
rect 19704 49978 19768 49982
rect 19704 49922 19708 49978
rect 19708 49922 19764 49978
rect 19764 49922 19768 49978
rect 19704 49918 19768 49922
rect 19784 49978 19848 49982
rect 19784 49922 19788 49978
rect 19788 49922 19844 49978
rect 19844 49922 19848 49978
rect 19784 49918 19848 49922
rect 19864 49978 19928 49982
rect 19864 49922 19868 49978
rect 19868 49922 19924 49978
rect 19924 49922 19928 49978
rect 19864 49918 19928 49922
rect 50344 49978 50408 49982
rect 50344 49922 50348 49978
rect 50348 49922 50404 49978
rect 50404 49922 50408 49978
rect 50344 49918 50408 49922
rect 50424 49978 50488 49982
rect 50424 49922 50428 49978
rect 50428 49922 50484 49978
rect 50484 49922 50488 49978
rect 50424 49918 50488 49922
rect 50504 49978 50568 49982
rect 50504 49922 50508 49978
rect 50508 49922 50564 49978
rect 50564 49922 50568 49978
rect 50504 49918 50568 49922
rect 50584 49978 50648 49982
rect 50584 49922 50588 49978
rect 50588 49922 50644 49978
rect 50644 49922 50648 49978
rect 50584 49918 50648 49922
rect 4264 49312 4328 49316
rect 4264 49256 4268 49312
rect 4268 49256 4324 49312
rect 4324 49256 4328 49312
rect 4264 49252 4328 49256
rect 4344 49312 4408 49316
rect 4344 49256 4348 49312
rect 4348 49256 4404 49312
rect 4404 49256 4408 49312
rect 4344 49252 4408 49256
rect 4424 49312 4488 49316
rect 4424 49256 4428 49312
rect 4428 49256 4484 49312
rect 4484 49256 4488 49312
rect 4424 49252 4488 49256
rect 4504 49312 4568 49316
rect 4504 49256 4508 49312
rect 4508 49256 4564 49312
rect 4564 49256 4568 49312
rect 4504 49252 4568 49256
rect 34984 49312 35048 49316
rect 34984 49256 34988 49312
rect 34988 49256 35044 49312
rect 35044 49256 35048 49312
rect 34984 49252 35048 49256
rect 35064 49312 35128 49316
rect 35064 49256 35068 49312
rect 35068 49256 35124 49312
rect 35124 49256 35128 49312
rect 35064 49252 35128 49256
rect 35144 49312 35208 49316
rect 35144 49256 35148 49312
rect 35148 49256 35204 49312
rect 35204 49256 35208 49312
rect 35144 49252 35208 49256
rect 35224 49312 35288 49316
rect 35224 49256 35228 49312
rect 35228 49256 35284 49312
rect 35284 49256 35288 49312
rect 35224 49252 35288 49256
rect 19624 48646 19688 48650
rect 19624 48590 19628 48646
rect 19628 48590 19684 48646
rect 19684 48590 19688 48646
rect 19624 48586 19688 48590
rect 19704 48646 19768 48650
rect 19704 48590 19708 48646
rect 19708 48590 19764 48646
rect 19764 48590 19768 48646
rect 19704 48586 19768 48590
rect 19784 48646 19848 48650
rect 19784 48590 19788 48646
rect 19788 48590 19844 48646
rect 19844 48590 19848 48646
rect 19784 48586 19848 48590
rect 19864 48646 19928 48650
rect 19864 48590 19868 48646
rect 19868 48590 19924 48646
rect 19924 48590 19928 48646
rect 19864 48586 19928 48590
rect 50344 48646 50408 48650
rect 50344 48590 50348 48646
rect 50348 48590 50404 48646
rect 50404 48590 50408 48646
rect 50344 48586 50408 48590
rect 50424 48646 50488 48650
rect 50424 48590 50428 48646
rect 50428 48590 50484 48646
rect 50484 48590 50488 48646
rect 50424 48586 50488 48590
rect 50504 48646 50568 48650
rect 50504 48590 50508 48646
rect 50508 48590 50564 48646
rect 50564 48590 50568 48646
rect 50504 48586 50568 48590
rect 50584 48646 50648 48650
rect 50584 48590 50588 48646
rect 50588 48590 50644 48646
rect 50644 48590 50648 48646
rect 50584 48586 50648 48590
rect 4264 47980 4328 47984
rect 4264 47924 4268 47980
rect 4268 47924 4324 47980
rect 4324 47924 4328 47980
rect 4264 47920 4328 47924
rect 4344 47980 4408 47984
rect 4344 47924 4348 47980
rect 4348 47924 4404 47980
rect 4404 47924 4408 47980
rect 4344 47920 4408 47924
rect 4424 47980 4488 47984
rect 4424 47924 4428 47980
rect 4428 47924 4484 47980
rect 4484 47924 4488 47980
rect 4424 47920 4488 47924
rect 4504 47980 4568 47984
rect 4504 47924 4508 47980
rect 4508 47924 4564 47980
rect 4564 47924 4568 47980
rect 4504 47920 4568 47924
rect 34984 47980 35048 47984
rect 34984 47924 34988 47980
rect 34988 47924 35044 47980
rect 35044 47924 35048 47980
rect 34984 47920 35048 47924
rect 35064 47980 35128 47984
rect 35064 47924 35068 47980
rect 35068 47924 35124 47980
rect 35124 47924 35128 47980
rect 35064 47920 35128 47924
rect 35144 47980 35208 47984
rect 35144 47924 35148 47980
rect 35148 47924 35204 47980
rect 35204 47924 35208 47980
rect 35144 47920 35208 47924
rect 35224 47980 35288 47984
rect 35224 47924 35228 47980
rect 35228 47924 35284 47980
rect 35284 47924 35288 47980
rect 35224 47920 35288 47924
rect 19624 47314 19688 47318
rect 19624 47258 19628 47314
rect 19628 47258 19684 47314
rect 19684 47258 19688 47314
rect 19624 47254 19688 47258
rect 19704 47314 19768 47318
rect 19704 47258 19708 47314
rect 19708 47258 19764 47314
rect 19764 47258 19768 47314
rect 19704 47254 19768 47258
rect 19784 47314 19848 47318
rect 19784 47258 19788 47314
rect 19788 47258 19844 47314
rect 19844 47258 19848 47314
rect 19784 47254 19848 47258
rect 19864 47314 19928 47318
rect 19864 47258 19868 47314
rect 19868 47258 19924 47314
rect 19924 47258 19928 47314
rect 19864 47254 19928 47258
rect 50344 47314 50408 47318
rect 50344 47258 50348 47314
rect 50348 47258 50404 47314
rect 50404 47258 50408 47314
rect 50344 47254 50408 47258
rect 50424 47314 50488 47318
rect 50424 47258 50428 47314
rect 50428 47258 50484 47314
rect 50484 47258 50488 47314
rect 50424 47254 50488 47258
rect 50504 47314 50568 47318
rect 50504 47258 50508 47314
rect 50508 47258 50564 47314
rect 50564 47258 50568 47314
rect 50504 47254 50568 47258
rect 50584 47314 50648 47318
rect 50584 47258 50588 47314
rect 50588 47258 50644 47314
rect 50644 47258 50648 47314
rect 50584 47254 50648 47258
rect 4264 46648 4328 46652
rect 4264 46592 4268 46648
rect 4268 46592 4324 46648
rect 4324 46592 4328 46648
rect 4264 46588 4328 46592
rect 4344 46648 4408 46652
rect 4344 46592 4348 46648
rect 4348 46592 4404 46648
rect 4404 46592 4408 46648
rect 4344 46588 4408 46592
rect 4424 46648 4488 46652
rect 4424 46592 4428 46648
rect 4428 46592 4484 46648
rect 4484 46592 4488 46648
rect 4424 46588 4488 46592
rect 4504 46648 4568 46652
rect 4504 46592 4508 46648
rect 4508 46592 4564 46648
rect 4564 46592 4568 46648
rect 4504 46588 4568 46592
rect 34984 46648 35048 46652
rect 34984 46592 34988 46648
rect 34988 46592 35044 46648
rect 35044 46592 35048 46648
rect 34984 46588 35048 46592
rect 35064 46648 35128 46652
rect 35064 46592 35068 46648
rect 35068 46592 35124 46648
rect 35124 46592 35128 46648
rect 35064 46588 35128 46592
rect 35144 46648 35208 46652
rect 35144 46592 35148 46648
rect 35148 46592 35204 46648
rect 35204 46592 35208 46648
rect 35144 46588 35208 46592
rect 35224 46648 35288 46652
rect 35224 46592 35228 46648
rect 35228 46592 35284 46648
rect 35284 46592 35288 46648
rect 35224 46588 35288 46592
rect 19624 45982 19688 45986
rect 19624 45926 19628 45982
rect 19628 45926 19684 45982
rect 19684 45926 19688 45982
rect 19624 45922 19688 45926
rect 19704 45982 19768 45986
rect 19704 45926 19708 45982
rect 19708 45926 19764 45982
rect 19764 45926 19768 45982
rect 19704 45922 19768 45926
rect 19784 45982 19848 45986
rect 19784 45926 19788 45982
rect 19788 45926 19844 45982
rect 19844 45926 19848 45982
rect 19784 45922 19848 45926
rect 19864 45982 19928 45986
rect 19864 45926 19868 45982
rect 19868 45926 19924 45982
rect 19924 45926 19928 45982
rect 19864 45922 19928 45926
rect 50344 45982 50408 45986
rect 50344 45926 50348 45982
rect 50348 45926 50404 45982
rect 50404 45926 50408 45982
rect 50344 45922 50408 45926
rect 50424 45982 50488 45986
rect 50424 45926 50428 45982
rect 50428 45926 50484 45982
rect 50484 45926 50488 45982
rect 50424 45922 50488 45926
rect 50504 45982 50568 45986
rect 50504 45926 50508 45982
rect 50508 45926 50564 45982
rect 50564 45926 50568 45982
rect 50504 45922 50568 45926
rect 50584 45982 50648 45986
rect 50584 45926 50588 45982
rect 50588 45926 50644 45982
rect 50644 45926 50648 45982
rect 50584 45922 50648 45926
rect 4264 45316 4328 45320
rect 4264 45260 4268 45316
rect 4268 45260 4324 45316
rect 4324 45260 4328 45316
rect 4264 45256 4328 45260
rect 4344 45316 4408 45320
rect 4344 45260 4348 45316
rect 4348 45260 4404 45316
rect 4404 45260 4408 45316
rect 4344 45256 4408 45260
rect 4424 45316 4488 45320
rect 4424 45260 4428 45316
rect 4428 45260 4484 45316
rect 4484 45260 4488 45316
rect 4424 45256 4488 45260
rect 4504 45316 4568 45320
rect 4504 45260 4508 45316
rect 4508 45260 4564 45316
rect 4564 45260 4568 45316
rect 4504 45256 4568 45260
rect 34984 45316 35048 45320
rect 34984 45260 34988 45316
rect 34988 45260 35044 45316
rect 35044 45260 35048 45316
rect 34984 45256 35048 45260
rect 35064 45316 35128 45320
rect 35064 45260 35068 45316
rect 35068 45260 35124 45316
rect 35124 45260 35128 45316
rect 35064 45256 35128 45260
rect 35144 45316 35208 45320
rect 35144 45260 35148 45316
rect 35148 45260 35204 45316
rect 35204 45260 35208 45316
rect 35144 45256 35208 45260
rect 35224 45316 35288 45320
rect 35224 45260 35228 45316
rect 35228 45260 35284 45316
rect 35284 45260 35288 45316
rect 35224 45256 35288 45260
rect 19624 44650 19688 44654
rect 19624 44594 19628 44650
rect 19628 44594 19684 44650
rect 19684 44594 19688 44650
rect 19624 44590 19688 44594
rect 19704 44650 19768 44654
rect 19704 44594 19708 44650
rect 19708 44594 19764 44650
rect 19764 44594 19768 44650
rect 19704 44590 19768 44594
rect 19784 44650 19848 44654
rect 19784 44594 19788 44650
rect 19788 44594 19844 44650
rect 19844 44594 19848 44650
rect 19784 44590 19848 44594
rect 19864 44650 19928 44654
rect 19864 44594 19868 44650
rect 19868 44594 19924 44650
rect 19924 44594 19928 44650
rect 19864 44590 19928 44594
rect 50344 44650 50408 44654
rect 50344 44594 50348 44650
rect 50348 44594 50404 44650
rect 50404 44594 50408 44650
rect 50344 44590 50408 44594
rect 50424 44650 50488 44654
rect 50424 44594 50428 44650
rect 50428 44594 50484 44650
rect 50484 44594 50488 44650
rect 50424 44590 50488 44594
rect 50504 44650 50568 44654
rect 50504 44594 50508 44650
rect 50508 44594 50564 44650
rect 50564 44594 50568 44650
rect 50504 44590 50568 44594
rect 50584 44650 50648 44654
rect 50584 44594 50588 44650
rect 50588 44594 50644 44650
rect 50644 44594 50648 44650
rect 50584 44590 50648 44594
rect 4264 43984 4328 43988
rect 4264 43928 4268 43984
rect 4268 43928 4324 43984
rect 4324 43928 4328 43984
rect 4264 43924 4328 43928
rect 4344 43984 4408 43988
rect 4344 43928 4348 43984
rect 4348 43928 4404 43984
rect 4404 43928 4408 43984
rect 4344 43924 4408 43928
rect 4424 43984 4488 43988
rect 4424 43928 4428 43984
rect 4428 43928 4484 43984
rect 4484 43928 4488 43984
rect 4424 43924 4488 43928
rect 4504 43984 4568 43988
rect 4504 43928 4508 43984
rect 4508 43928 4564 43984
rect 4564 43928 4568 43984
rect 4504 43924 4568 43928
rect 34984 43984 35048 43988
rect 34984 43928 34988 43984
rect 34988 43928 35044 43984
rect 35044 43928 35048 43984
rect 34984 43924 35048 43928
rect 35064 43984 35128 43988
rect 35064 43928 35068 43984
rect 35068 43928 35124 43984
rect 35124 43928 35128 43984
rect 35064 43924 35128 43928
rect 35144 43984 35208 43988
rect 35144 43928 35148 43984
rect 35148 43928 35204 43984
rect 35204 43928 35208 43984
rect 35144 43924 35208 43928
rect 35224 43984 35288 43988
rect 35224 43928 35228 43984
rect 35228 43928 35284 43984
rect 35284 43928 35288 43984
rect 35224 43924 35288 43928
rect 19624 43318 19688 43322
rect 19624 43262 19628 43318
rect 19628 43262 19684 43318
rect 19684 43262 19688 43318
rect 19624 43258 19688 43262
rect 19704 43318 19768 43322
rect 19704 43262 19708 43318
rect 19708 43262 19764 43318
rect 19764 43262 19768 43318
rect 19704 43258 19768 43262
rect 19784 43318 19848 43322
rect 19784 43262 19788 43318
rect 19788 43262 19844 43318
rect 19844 43262 19848 43318
rect 19784 43258 19848 43262
rect 19864 43318 19928 43322
rect 19864 43262 19868 43318
rect 19868 43262 19924 43318
rect 19924 43262 19928 43318
rect 19864 43258 19928 43262
rect 50344 43318 50408 43322
rect 50344 43262 50348 43318
rect 50348 43262 50404 43318
rect 50404 43262 50408 43318
rect 50344 43258 50408 43262
rect 50424 43318 50488 43322
rect 50424 43262 50428 43318
rect 50428 43262 50484 43318
rect 50484 43262 50488 43318
rect 50424 43258 50488 43262
rect 50504 43318 50568 43322
rect 50504 43262 50508 43318
rect 50508 43262 50564 43318
rect 50564 43262 50568 43318
rect 50504 43258 50568 43262
rect 50584 43318 50648 43322
rect 50584 43262 50588 43318
rect 50588 43262 50644 43318
rect 50644 43262 50648 43318
rect 50584 43258 50648 43262
rect 4264 42652 4328 42656
rect 4264 42596 4268 42652
rect 4268 42596 4324 42652
rect 4324 42596 4328 42652
rect 4264 42592 4328 42596
rect 4344 42652 4408 42656
rect 4344 42596 4348 42652
rect 4348 42596 4404 42652
rect 4404 42596 4408 42652
rect 4344 42592 4408 42596
rect 4424 42652 4488 42656
rect 4424 42596 4428 42652
rect 4428 42596 4484 42652
rect 4484 42596 4488 42652
rect 4424 42592 4488 42596
rect 4504 42652 4568 42656
rect 4504 42596 4508 42652
rect 4508 42596 4564 42652
rect 4564 42596 4568 42652
rect 4504 42592 4568 42596
rect 34984 42652 35048 42656
rect 34984 42596 34988 42652
rect 34988 42596 35044 42652
rect 35044 42596 35048 42652
rect 34984 42592 35048 42596
rect 35064 42652 35128 42656
rect 35064 42596 35068 42652
rect 35068 42596 35124 42652
rect 35124 42596 35128 42652
rect 35064 42592 35128 42596
rect 35144 42652 35208 42656
rect 35144 42596 35148 42652
rect 35148 42596 35204 42652
rect 35204 42596 35208 42652
rect 35144 42592 35208 42596
rect 35224 42652 35288 42656
rect 35224 42596 35228 42652
rect 35228 42596 35284 42652
rect 35284 42596 35288 42652
rect 35224 42592 35288 42596
rect 19624 41986 19688 41990
rect 19624 41930 19628 41986
rect 19628 41930 19684 41986
rect 19684 41930 19688 41986
rect 19624 41926 19688 41930
rect 19704 41986 19768 41990
rect 19704 41930 19708 41986
rect 19708 41930 19764 41986
rect 19764 41930 19768 41986
rect 19704 41926 19768 41930
rect 19784 41986 19848 41990
rect 19784 41930 19788 41986
rect 19788 41930 19844 41986
rect 19844 41930 19848 41986
rect 19784 41926 19848 41930
rect 19864 41986 19928 41990
rect 19864 41930 19868 41986
rect 19868 41930 19924 41986
rect 19924 41930 19928 41986
rect 19864 41926 19928 41930
rect 50344 41986 50408 41990
rect 50344 41930 50348 41986
rect 50348 41930 50404 41986
rect 50404 41930 50408 41986
rect 50344 41926 50408 41930
rect 50424 41986 50488 41990
rect 50424 41930 50428 41986
rect 50428 41930 50484 41986
rect 50484 41930 50488 41986
rect 50424 41926 50488 41930
rect 50504 41986 50568 41990
rect 50504 41930 50508 41986
rect 50508 41930 50564 41986
rect 50564 41930 50568 41986
rect 50504 41926 50568 41930
rect 50584 41986 50648 41990
rect 50584 41930 50588 41986
rect 50588 41930 50644 41986
rect 50644 41930 50648 41986
rect 50584 41926 50648 41930
rect 4264 41320 4328 41324
rect 4264 41264 4268 41320
rect 4268 41264 4324 41320
rect 4324 41264 4328 41320
rect 4264 41260 4328 41264
rect 4344 41320 4408 41324
rect 4344 41264 4348 41320
rect 4348 41264 4404 41320
rect 4404 41264 4408 41320
rect 4344 41260 4408 41264
rect 4424 41320 4488 41324
rect 4424 41264 4428 41320
rect 4428 41264 4484 41320
rect 4484 41264 4488 41320
rect 4424 41260 4488 41264
rect 4504 41320 4568 41324
rect 4504 41264 4508 41320
rect 4508 41264 4564 41320
rect 4564 41264 4568 41320
rect 4504 41260 4568 41264
rect 34984 41320 35048 41324
rect 34984 41264 34988 41320
rect 34988 41264 35044 41320
rect 35044 41264 35048 41320
rect 34984 41260 35048 41264
rect 35064 41320 35128 41324
rect 35064 41264 35068 41320
rect 35068 41264 35124 41320
rect 35124 41264 35128 41320
rect 35064 41260 35128 41264
rect 35144 41320 35208 41324
rect 35144 41264 35148 41320
rect 35148 41264 35204 41320
rect 35204 41264 35208 41320
rect 35144 41260 35208 41264
rect 35224 41320 35288 41324
rect 35224 41264 35228 41320
rect 35228 41264 35284 41320
rect 35284 41264 35288 41320
rect 35224 41260 35288 41264
rect 19624 40654 19688 40658
rect 19624 40598 19628 40654
rect 19628 40598 19684 40654
rect 19684 40598 19688 40654
rect 19624 40594 19688 40598
rect 19704 40654 19768 40658
rect 19704 40598 19708 40654
rect 19708 40598 19764 40654
rect 19764 40598 19768 40654
rect 19704 40594 19768 40598
rect 19784 40654 19848 40658
rect 19784 40598 19788 40654
rect 19788 40598 19844 40654
rect 19844 40598 19848 40654
rect 19784 40594 19848 40598
rect 19864 40654 19928 40658
rect 19864 40598 19868 40654
rect 19868 40598 19924 40654
rect 19924 40598 19928 40654
rect 19864 40594 19928 40598
rect 50344 40654 50408 40658
rect 50344 40598 50348 40654
rect 50348 40598 50404 40654
rect 50404 40598 50408 40654
rect 50344 40594 50408 40598
rect 50424 40654 50488 40658
rect 50424 40598 50428 40654
rect 50428 40598 50484 40654
rect 50484 40598 50488 40654
rect 50424 40594 50488 40598
rect 50504 40654 50568 40658
rect 50504 40598 50508 40654
rect 50508 40598 50564 40654
rect 50564 40598 50568 40654
rect 50504 40594 50568 40598
rect 50584 40654 50648 40658
rect 50584 40598 50588 40654
rect 50588 40598 50644 40654
rect 50644 40598 50648 40654
rect 50584 40594 50648 40598
rect 4264 39988 4328 39992
rect 4264 39932 4268 39988
rect 4268 39932 4324 39988
rect 4324 39932 4328 39988
rect 4264 39928 4328 39932
rect 4344 39988 4408 39992
rect 4344 39932 4348 39988
rect 4348 39932 4404 39988
rect 4404 39932 4408 39988
rect 4344 39928 4408 39932
rect 4424 39988 4488 39992
rect 4424 39932 4428 39988
rect 4428 39932 4484 39988
rect 4484 39932 4488 39988
rect 4424 39928 4488 39932
rect 4504 39988 4568 39992
rect 4504 39932 4508 39988
rect 4508 39932 4564 39988
rect 4564 39932 4568 39988
rect 4504 39928 4568 39932
rect 34984 39988 35048 39992
rect 34984 39932 34988 39988
rect 34988 39932 35044 39988
rect 35044 39932 35048 39988
rect 34984 39928 35048 39932
rect 35064 39988 35128 39992
rect 35064 39932 35068 39988
rect 35068 39932 35124 39988
rect 35124 39932 35128 39988
rect 35064 39928 35128 39932
rect 35144 39988 35208 39992
rect 35144 39932 35148 39988
rect 35148 39932 35204 39988
rect 35204 39932 35208 39988
rect 35144 39928 35208 39932
rect 35224 39988 35288 39992
rect 35224 39932 35228 39988
rect 35228 39932 35284 39988
rect 35284 39932 35288 39988
rect 35224 39928 35288 39932
rect 19624 39322 19688 39326
rect 19624 39266 19628 39322
rect 19628 39266 19684 39322
rect 19684 39266 19688 39322
rect 19624 39262 19688 39266
rect 19704 39322 19768 39326
rect 19704 39266 19708 39322
rect 19708 39266 19764 39322
rect 19764 39266 19768 39322
rect 19704 39262 19768 39266
rect 19784 39322 19848 39326
rect 19784 39266 19788 39322
rect 19788 39266 19844 39322
rect 19844 39266 19848 39322
rect 19784 39262 19848 39266
rect 19864 39322 19928 39326
rect 19864 39266 19868 39322
rect 19868 39266 19924 39322
rect 19924 39266 19928 39322
rect 19864 39262 19928 39266
rect 50344 39322 50408 39326
rect 50344 39266 50348 39322
rect 50348 39266 50404 39322
rect 50404 39266 50408 39322
rect 50344 39262 50408 39266
rect 50424 39322 50488 39326
rect 50424 39266 50428 39322
rect 50428 39266 50484 39322
rect 50484 39266 50488 39322
rect 50424 39262 50488 39266
rect 50504 39322 50568 39326
rect 50504 39266 50508 39322
rect 50508 39266 50564 39322
rect 50564 39266 50568 39322
rect 50504 39262 50568 39266
rect 50584 39322 50648 39326
rect 50584 39266 50588 39322
rect 50588 39266 50644 39322
rect 50644 39266 50648 39322
rect 50584 39262 50648 39266
rect 4264 38656 4328 38660
rect 4264 38600 4268 38656
rect 4268 38600 4324 38656
rect 4324 38600 4328 38656
rect 4264 38596 4328 38600
rect 4344 38656 4408 38660
rect 4344 38600 4348 38656
rect 4348 38600 4404 38656
rect 4404 38600 4408 38656
rect 4344 38596 4408 38600
rect 4424 38656 4488 38660
rect 4424 38600 4428 38656
rect 4428 38600 4484 38656
rect 4484 38600 4488 38656
rect 4424 38596 4488 38600
rect 4504 38656 4568 38660
rect 4504 38600 4508 38656
rect 4508 38600 4564 38656
rect 4564 38600 4568 38656
rect 4504 38596 4568 38600
rect 34984 38656 35048 38660
rect 34984 38600 34988 38656
rect 34988 38600 35044 38656
rect 35044 38600 35048 38656
rect 34984 38596 35048 38600
rect 35064 38656 35128 38660
rect 35064 38600 35068 38656
rect 35068 38600 35124 38656
rect 35124 38600 35128 38656
rect 35064 38596 35128 38600
rect 35144 38656 35208 38660
rect 35144 38600 35148 38656
rect 35148 38600 35204 38656
rect 35204 38600 35208 38656
rect 35144 38596 35208 38600
rect 35224 38656 35288 38660
rect 35224 38600 35228 38656
rect 35228 38600 35284 38656
rect 35284 38600 35288 38656
rect 35224 38596 35288 38600
rect 19624 37990 19688 37994
rect 19624 37934 19628 37990
rect 19628 37934 19684 37990
rect 19684 37934 19688 37990
rect 19624 37930 19688 37934
rect 19704 37990 19768 37994
rect 19704 37934 19708 37990
rect 19708 37934 19764 37990
rect 19764 37934 19768 37990
rect 19704 37930 19768 37934
rect 19784 37990 19848 37994
rect 19784 37934 19788 37990
rect 19788 37934 19844 37990
rect 19844 37934 19848 37990
rect 19784 37930 19848 37934
rect 19864 37990 19928 37994
rect 19864 37934 19868 37990
rect 19868 37934 19924 37990
rect 19924 37934 19928 37990
rect 19864 37930 19928 37934
rect 50344 37990 50408 37994
rect 50344 37934 50348 37990
rect 50348 37934 50404 37990
rect 50404 37934 50408 37990
rect 50344 37930 50408 37934
rect 50424 37990 50488 37994
rect 50424 37934 50428 37990
rect 50428 37934 50484 37990
rect 50484 37934 50488 37990
rect 50424 37930 50488 37934
rect 50504 37990 50568 37994
rect 50504 37934 50508 37990
rect 50508 37934 50564 37990
rect 50564 37934 50568 37990
rect 50504 37930 50568 37934
rect 50584 37990 50648 37994
rect 50584 37934 50588 37990
rect 50588 37934 50644 37990
rect 50644 37934 50648 37990
rect 50584 37930 50648 37934
rect 4264 37324 4328 37328
rect 4264 37268 4268 37324
rect 4268 37268 4324 37324
rect 4324 37268 4328 37324
rect 4264 37264 4328 37268
rect 4344 37324 4408 37328
rect 4344 37268 4348 37324
rect 4348 37268 4404 37324
rect 4404 37268 4408 37324
rect 4344 37264 4408 37268
rect 4424 37324 4488 37328
rect 4424 37268 4428 37324
rect 4428 37268 4484 37324
rect 4484 37268 4488 37324
rect 4424 37264 4488 37268
rect 4504 37324 4568 37328
rect 4504 37268 4508 37324
rect 4508 37268 4564 37324
rect 4564 37268 4568 37324
rect 4504 37264 4568 37268
rect 34984 37324 35048 37328
rect 34984 37268 34988 37324
rect 34988 37268 35044 37324
rect 35044 37268 35048 37324
rect 34984 37264 35048 37268
rect 35064 37324 35128 37328
rect 35064 37268 35068 37324
rect 35068 37268 35124 37324
rect 35124 37268 35128 37324
rect 35064 37264 35128 37268
rect 35144 37324 35208 37328
rect 35144 37268 35148 37324
rect 35148 37268 35204 37324
rect 35204 37268 35208 37324
rect 35144 37264 35208 37268
rect 35224 37324 35288 37328
rect 35224 37268 35228 37324
rect 35228 37268 35284 37324
rect 35284 37268 35288 37324
rect 35224 37264 35288 37268
rect 19624 36658 19688 36662
rect 19624 36602 19628 36658
rect 19628 36602 19684 36658
rect 19684 36602 19688 36658
rect 19624 36598 19688 36602
rect 19704 36658 19768 36662
rect 19704 36602 19708 36658
rect 19708 36602 19764 36658
rect 19764 36602 19768 36658
rect 19704 36598 19768 36602
rect 19784 36658 19848 36662
rect 19784 36602 19788 36658
rect 19788 36602 19844 36658
rect 19844 36602 19848 36658
rect 19784 36598 19848 36602
rect 19864 36658 19928 36662
rect 19864 36602 19868 36658
rect 19868 36602 19924 36658
rect 19924 36602 19928 36658
rect 19864 36598 19928 36602
rect 50344 36658 50408 36662
rect 50344 36602 50348 36658
rect 50348 36602 50404 36658
rect 50404 36602 50408 36658
rect 50344 36598 50408 36602
rect 50424 36658 50488 36662
rect 50424 36602 50428 36658
rect 50428 36602 50484 36658
rect 50484 36602 50488 36658
rect 50424 36598 50488 36602
rect 50504 36658 50568 36662
rect 50504 36602 50508 36658
rect 50508 36602 50564 36658
rect 50564 36602 50568 36658
rect 50504 36598 50568 36602
rect 50584 36658 50648 36662
rect 50584 36602 50588 36658
rect 50588 36602 50644 36658
rect 50644 36602 50648 36658
rect 50584 36598 50648 36602
rect 4264 35992 4328 35996
rect 4264 35936 4268 35992
rect 4268 35936 4324 35992
rect 4324 35936 4328 35992
rect 4264 35932 4328 35936
rect 4344 35992 4408 35996
rect 4344 35936 4348 35992
rect 4348 35936 4404 35992
rect 4404 35936 4408 35992
rect 4344 35932 4408 35936
rect 4424 35992 4488 35996
rect 4424 35936 4428 35992
rect 4428 35936 4484 35992
rect 4484 35936 4488 35992
rect 4424 35932 4488 35936
rect 4504 35992 4568 35996
rect 4504 35936 4508 35992
rect 4508 35936 4564 35992
rect 4564 35936 4568 35992
rect 4504 35932 4568 35936
rect 34984 35992 35048 35996
rect 34984 35936 34988 35992
rect 34988 35936 35044 35992
rect 35044 35936 35048 35992
rect 34984 35932 35048 35936
rect 35064 35992 35128 35996
rect 35064 35936 35068 35992
rect 35068 35936 35124 35992
rect 35124 35936 35128 35992
rect 35064 35932 35128 35936
rect 35144 35992 35208 35996
rect 35144 35936 35148 35992
rect 35148 35936 35204 35992
rect 35204 35936 35208 35992
rect 35144 35932 35208 35936
rect 35224 35992 35288 35996
rect 35224 35936 35228 35992
rect 35228 35936 35284 35992
rect 35284 35936 35288 35992
rect 35224 35932 35288 35936
rect 19624 35326 19688 35330
rect 19624 35270 19628 35326
rect 19628 35270 19684 35326
rect 19684 35270 19688 35326
rect 19624 35266 19688 35270
rect 19704 35326 19768 35330
rect 19704 35270 19708 35326
rect 19708 35270 19764 35326
rect 19764 35270 19768 35326
rect 19704 35266 19768 35270
rect 19784 35326 19848 35330
rect 19784 35270 19788 35326
rect 19788 35270 19844 35326
rect 19844 35270 19848 35326
rect 19784 35266 19848 35270
rect 19864 35326 19928 35330
rect 19864 35270 19868 35326
rect 19868 35270 19924 35326
rect 19924 35270 19928 35326
rect 19864 35266 19928 35270
rect 50344 35326 50408 35330
rect 50344 35270 50348 35326
rect 50348 35270 50404 35326
rect 50404 35270 50408 35326
rect 50344 35266 50408 35270
rect 50424 35326 50488 35330
rect 50424 35270 50428 35326
rect 50428 35270 50484 35326
rect 50484 35270 50488 35326
rect 50424 35266 50488 35270
rect 50504 35326 50568 35330
rect 50504 35270 50508 35326
rect 50508 35270 50564 35326
rect 50564 35270 50568 35326
rect 50504 35266 50568 35270
rect 50584 35326 50648 35330
rect 50584 35270 50588 35326
rect 50588 35270 50644 35326
rect 50644 35270 50648 35326
rect 50584 35266 50648 35270
rect 4264 34660 4328 34664
rect 4264 34604 4268 34660
rect 4268 34604 4324 34660
rect 4324 34604 4328 34660
rect 4264 34600 4328 34604
rect 4344 34660 4408 34664
rect 4344 34604 4348 34660
rect 4348 34604 4404 34660
rect 4404 34604 4408 34660
rect 4344 34600 4408 34604
rect 4424 34660 4488 34664
rect 4424 34604 4428 34660
rect 4428 34604 4484 34660
rect 4484 34604 4488 34660
rect 4424 34600 4488 34604
rect 4504 34660 4568 34664
rect 4504 34604 4508 34660
rect 4508 34604 4564 34660
rect 4564 34604 4568 34660
rect 4504 34600 4568 34604
rect 34984 34660 35048 34664
rect 34984 34604 34988 34660
rect 34988 34604 35044 34660
rect 35044 34604 35048 34660
rect 34984 34600 35048 34604
rect 35064 34660 35128 34664
rect 35064 34604 35068 34660
rect 35068 34604 35124 34660
rect 35124 34604 35128 34660
rect 35064 34600 35128 34604
rect 35144 34660 35208 34664
rect 35144 34604 35148 34660
rect 35148 34604 35204 34660
rect 35204 34604 35208 34660
rect 35144 34600 35208 34604
rect 35224 34660 35288 34664
rect 35224 34604 35228 34660
rect 35228 34604 35284 34660
rect 35284 34604 35288 34660
rect 35224 34600 35288 34604
rect 19624 33994 19688 33998
rect 19624 33938 19628 33994
rect 19628 33938 19684 33994
rect 19684 33938 19688 33994
rect 19624 33934 19688 33938
rect 19704 33994 19768 33998
rect 19704 33938 19708 33994
rect 19708 33938 19764 33994
rect 19764 33938 19768 33994
rect 19704 33934 19768 33938
rect 19784 33994 19848 33998
rect 19784 33938 19788 33994
rect 19788 33938 19844 33994
rect 19844 33938 19848 33994
rect 19784 33934 19848 33938
rect 19864 33994 19928 33998
rect 19864 33938 19868 33994
rect 19868 33938 19924 33994
rect 19924 33938 19928 33994
rect 19864 33934 19928 33938
rect 50344 33994 50408 33998
rect 50344 33938 50348 33994
rect 50348 33938 50404 33994
rect 50404 33938 50408 33994
rect 50344 33934 50408 33938
rect 50424 33994 50488 33998
rect 50424 33938 50428 33994
rect 50428 33938 50484 33994
rect 50484 33938 50488 33994
rect 50424 33934 50488 33938
rect 50504 33994 50568 33998
rect 50504 33938 50508 33994
rect 50508 33938 50564 33994
rect 50564 33938 50568 33994
rect 50504 33934 50568 33938
rect 50584 33994 50648 33998
rect 50584 33938 50588 33994
rect 50588 33938 50644 33994
rect 50644 33938 50648 33994
rect 50584 33934 50648 33938
rect 4264 33328 4328 33332
rect 4264 33272 4268 33328
rect 4268 33272 4324 33328
rect 4324 33272 4328 33328
rect 4264 33268 4328 33272
rect 4344 33328 4408 33332
rect 4344 33272 4348 33328
rect 4348 33272 4404 33328
rect 4404 33272 4408 33328
rect 4344 33268 4408 33272
rect 4424 33328 4488 33332
rect 4424 33272 4428 33328
rect 4428 33272 4484 33328
rect 4484 33272 4488 33328
rect 4424 33268 4488 33272
rect 4504 33328 4568 33332
rect 4504 33272 4508 33328
rect 4508 33272 4564 33328
rect 4564 33272 4568 33328
rect 4504 33268 4568 33272
rect 34984 33328 35048 33332
rect 34984 33272 34988 33328
rect 34988 33272 35044 33328
rect 35044 33272 35048 33328
rect 34984 33268 35048 33272
rect 35064 33328 35128 33332
rect 35064 33272 35068 33328
rect 35068 33272 35124 33328
rect 35124 33272 35128 33328
rect 35064 33268 35128 33272
rect 35144 33328 35208 33332
rect 35144 33272 35148 33328
rect 35148 33272 35204 33328
rect 35204 33272 35208 33328
rect 35144 33268 35208 33272
rect 35224 33328 35288 33332
rect 35224 33272 35228 33328
rect 35228 33272 35284 33328
rect 35284 33272 35288 33328
rect 35224 33268 35288 33272
rect 19624 32662 19688 32666
rect 19624 32606 19628 32662
rect 19628 32606 19684 32662
rect 19684 32606 19688 32662
rect 19624 32602 19688 32606
rect 19704 32662 19768 32666
rect 19704 32606 19708 32662
rect 19708 32606 19764 32662
rect 19764 32606 19768 32662
rect 19704 32602 19768 32606
rect 19784 32662 19848 32666
rect 19784 32606 19788 32662
rect 19788 32606 19844 32662
rect 19844 32606 19848 32662
rect 19784 32602 19848 32606
rect 19864 32662 19928 32666
rect 19864 32606 19868 32662
rect 19868 32606 19924 32662
rect 19924 32606 19928 32662
rect 19864 32602 19928 32606
rect 50344 32662 50408 32666
rect 50344 32606 50348 32662
rect 50348 32606 50404 32662
rect 50404 32606 50408 32662
rect 50344 32602 50408 32606
rect 50424 32662 50488 32666
rect 50424 32606 50428 32662
rect 50428 32606 50484 32662
rect 50484 32606 50488 32662
rect 50424 32602 50488 32606
rect 50504 32662 50568 32666
rect 50504 32606 50508 32662
rect 50508 32606 50564 32662
rect 50564 32606 50568 32662
rect 50504 32602 50568 32606
rect 50584 32662 50648 32666
rect 50584 32606 50588 32662
rect 50588 32606 50644 32662
rect 50644 32606 50648 32662
rect 50584 32602 50648 32606
rect 4264 31996 4328 32000
rect 4264 31940 4268 31996
rect 4268 31940 4324 31996
rect 4324 31940 4328 31996
rect 4264 31936 4328 31940
rect 4344 31996 4408 32000
rect 4344 31940 4348 31996
rect 4348 31940 4404 31996
rect 4404 31940 4408 31996
rect 4344 31936 4408 31940
rect 4424 31996 4488 32000
rect 4424 31940 4428 31996
rect 4428 31940 4484 31996
rect 4484 31940 4488 31996
rect 4424 31936 4488 31940
rect 4504 31996 4568 32000
rect 4504 31940 4508 31996
rect 4508 31940 4564 31996
rect 4564 31940 4568 31996
rect 4504 31936 4568 31940
rect 34984 31996 35048 32000
rect 34984 31940 34988 31996
rect 34988 31940 35044 31996
rect 35044 31940 35048 31996
rect 34984 31936 35048 31940
rect 35064 31996 35128 32000
rect 35064 31940 35068 31996
rect 35068 31940 35124 31996
rect 35124 31940 35128 31996
rect 35064 31936 35128 31940
rect 35144 31996 35208 32000
rect 35144 31940 35148 31996
rect 35148 31940 35204 31996
rect 35204 31940 35208 31996
rect 35144 31936 35208 31940
rect 35224 31996 35288 32000
rect 35224 31940 35228 31996
rect 35228 31940 35284 31996
rect 35284 31940 35288 31996
rect 35224 31936 35288 31940
rect 19624 31330 19688 31334
rect 19624 31274 19628 31330
rect 19628 31274 19684 31330
rect 19684 31274 19688 31330
rect 19624 31270 19688 31274
rect 19704 31330 19768 31334
rect 19704 31274 19708 31330
rect 19708 31274 19764 31330
rect 19764 31274 19768 31330
rect 19704 31270 19768 31274
rect 19784 31330 19848 31334
rect 19784 31274 19788 31330
rect 19788 31274 19844 31330
rect 19844 31274 19848 31330
rect 19784 31270 19848 31274
rect 19864 31330 19928 31334
rect 19864 31274 19868 31330
rect 19868 31274 19924 31330
rect 19924 31274 19928 31330
rect 19864 31270 19928 31274
rect 50344 31330 50408 31334
rect 50344 31274 50348 31330
rect 50348 31274 50404 31330
rect 50404 31274 50408 31330
rect 50344 31270 50408 31274
rect 50424 31330 50488 31334
rect 50424 31274 50428 31330
rect 50428 31274 50484 31330
rect 50484 31274 50488 31330
rect 50424 31270 50488 31274
rect 50504 31330 50568 31334
rect 50504 31274 50508 31330
rect 50508 31274 50564 31330
rect 50564 31274 50568 31330
rect 50504 31270 50568 31274
rect 50584 31330 50648 31334
rect 50584 31274 50588 31330
rect 50588 31274 50644 31330
rect 50644 31274 50648 31330
rect 50584 31270 50648 31274
rect 4264 30664 4328 30668
rect 4264 30608 4268 30664
rect 4268 30608 4324 30664
rect 4324 30608 4328 30664
rect 4264 30604 4328 30608
rect 4344 30664 4408 30668
rect 4344 30608 4348 30664
rect 4348 30608 4404 30664
rect 4404 30608 4408 30664
rect 4344 30604 4408 30608
rect 4424 30664 4488 30668
rect 4424 30608 4428 30664
rect 4428 30608 4484 30664
rect 4484 30608 4488 30664
rect 4424 30604 4488 30608
rect 4504 30664 4568 30668
rect 4504 30608 4508 30664
rect 4508 30608 4564 30664
rect 4564 30608 4568 30664
rect 4504 30604 4568 30608
rect 34984 30664 35048 30668
rect 34984 30608 34988 30664
rect 34988 30608 35044 30664
rect 35044 30608 35048 30664
rect 34984 30604 35048 30608
rect 35064 30664 35128 30668
rect 35064 30608 35068 30664
rect 35068 30608 35124 30664
rect 35124 30608 35128 30664
rect 35064 30604 35128 30608
rect 35144 30664 35208 30668
rect 35144 30608 35148 30664
rect 35148 30608 35204 30664
rect 35204 30608 35208 30664
rect 35144 30604 35208 30608
rect 35224 30664 35288 30668
rect 35224 30608 35228 30664
rect 35228 30608 35284 30664
rect 35284 30608 35288 30664
rect 35224 30604 35288 30608
rect 19624 29998 19688 30002
rect 19624 29942 19628 29998
rect 19628 29942 19684 29998
rect 19684 29942 19688 29998
rect 19624 29938 19688 29942
rect 19704 29998 19768 30002
rect 19704 29942 19708 29998
rect 19708 29942 19764 29998
rect 19764 29942 19768 29998
rect 19704 29938 19768 29942
rect 19784 29998 19848 30002
rect 19784 29942 19788 29998
rect 19788 29942 19844 29998
rect 19844 29942 19848 29998
rect 19784 29938 19848 29942
rect 19864 29998 19928 30002
rect 19864 29942 19868 29998
rect 19868 29942 19924 29998
rect 19924 29942 19928 29998
rect 19864 29938 19928 29942
rect 50344 29998 50408 30002
rect 50344 29942 50348 29998
rect 50348 29942 50404 29998
rect 50404 29942 50408 29998
rect 50344 29938 50408 29942
rect 50424 29998 50488 30002
rect 50424 29942 50428 29998
rect 50428 29942 50484 29998
rect 50484 29942 50488 29998
rect 50424 29938 50488 29942
rect 50504 29998 50568 30002
rect 50504 29942 50508 29998
rect 50508 29942 50564 29998
rect 50564 29942 50568 29998
rect 50504 29938 50568 29942
rect 50584 29998 50648 30002
rect 50584 29942 50588 29998
rect 50588 29942 50644 29998
rect 50644 29942 50648 29998
rect 50584 29938 50648 29942
rect 4264 29332 4328 29336
rect 4264 29276 4268 29332
rect 4268 29276 4324 29332
rect 4324 29276 4328 29332
rect 4264 29272 4328 29276
rect 4344 29332 4408 29336
rect 4344 29276 4348 29332
rect 4348 29276 4404 29332
rect 4404 29276 4408 29332
rect 4344 29272 4408 29276
rect 4424 29332 4488 29336
rect 4424 29276 4428 29332
rect 4428 29276 4484 29332
rect 4484 29276 4488 29332
rect 4424 29272 4488 29276
rect 4504 29332 4568 29336
rect 4504 29276 4508 29332
rect 4508 29276 4564 29332
rect 4564 29276 4568 29332
rect 4504 29272 4568 29276
rect 34984 29332 35048 29336
rect 34984 29276 34988 29332
rect 34988 29276 35044 29332
rect 35044 29276 35048 29332
rect 34984 29272 35048 29276
rect 35064 29332 35128 29336
rect 35064 29276 35068 29332
rect 35068 29276 35124 29332
rect 35124 29276 35128 29332
rect 35064 29272 35128 29276
rect 35144 29332 35208 29336
rect 35144 29276 35148 29332
rect 35148 29276 35204 29332
rect 35204 29276 35208 29332
rect 35144 29272 35208 29276
rect 35224 29332 35288 29336
rect 35224 29276 35228 29332
rect 35228 29276 35284 29332
rect 35284 29276 35288 29332
rect 35224 29272 35288 29276
rect 19624 28666 19688 28670
rect 19624 28610 19628 28666
rect 19628 28610 19684 28666
rect 19684 28610 19688 28666
rect 19624 28606 19688 28610
rect 19704 28666 19768 28670
rect 19704 28610 19708 28666
rect 19708 28610 19764 28666
rect 19764 28610 19768 28666
rect 19704 28606 19768 28610
rect 19784 28666 19848 28670
rect 19784 28610 19788 28666
rect 19788 28610 19844 28666
rect 19844 28610 19848 28666
rect 19784 28606 19848 28610
rect 19864 28666 19928 28670
rect 19864 28610 19868 28666
rect 19868 28610 19924 28666
rect 19924 28610 19928 28666
rect 19864 28606 19928 28610
rect 50344 28666 50408 28670
rect 50344 28610 50348 28666
rect 50348 28610 50404 28666
rect 50404 28610 50408 28666
rect 50344 28606 50408 28610
rect 50424 28666 50488 28670
rect 50424 28610 50428 28666
rect 50428 28610 50484 28666
rect 50484 28610 50488 28666
rect 50424 28606 50488 28610
rect 50504 28666 50568 28670
rect 50504 28610 50508 28666
rect 50508 28610 50564 28666
rect 50564 28610 50568 28666
rect 50504 28606 50568 28610
rect 50584 28666 50648 28670
rect 50584 28610 50588 28666
rect 50588 28610 50644 28666
rect 50644 28610 50648 28666
rect 50584 28606 50648 28610
rect 4264 28000 4328 28004
rect 4264 27944 4268 28000
rect 4268 27944 4324 28000
rect 4324 27944 4328 28000
rect 4264 27940 4328 27944
rect 4344 28000 4408 28004
rect 4344 27944 4348 28000
rect 4348 27944 4404 28000
rect 4404 27944 4408 28000
rect 4344 27940 4408 27944
rect 4424 28000 4488 28004
rect 4424 27944 4428 28000
rect 4428 27944 4484 28000
rect 4484 27944 4488 28000
rect 4424 27940 4488 27944
rect 4504 28000 4568 28004
rect 4504 27944 4508 28000
rect 4508 27944 4564 28000
rect 4564 27944 4568 28000
rect 4504 27940 4568 27944
rect 34984 28000 35048 28004
rect 34984 27944 34988 28000
rect 34988 27944 35044 28000
rect 35044 27944 35048 28000
rect 34984 27940 35048 27944
rect 35064 28000 35128 28004
rect 35064 27944 35068 28000
rect 35068 27944 35124 28000
rect 35124 27944 35128 28000
rect 35064 27940 35128 27944
rect 35144 28000 35208 28004
rect 35144 27944 35148 28000
rect 35148 27944 35204 28000
rect 35204 27944 35208 28000
rect 35144 27940 35208 27944
rect 35224 28000 35288 28004
rect 35224 27944 35228 28000
rect 35228 27944 35284 28000
rect 35284 27944 35288 28000
rect 35224 27940 35288 27944
rect 19624 27334 19688 27338
rect 19624 27278 19628 27334
rect 19628 27278 19684 27334
rect 19684 27278 19688 27334
rect 19624 27274 19688 27278
rect 19704 27334 19768 27338
rect 19704 27278 19708 27334
rect 19708 27278 19764 27334
rect 19764 27278 19768 27334
rect 19704 27274 19768 27278
rect 19784 27334 19848 27338
rect 19784 27278 19788 27334
rect 19788 27278 19844 27334
rect 19844 27278 19848 27334
rect 19784 27274 19848 27278
rect 19864 27334 19928 27338
rect 19864 27278 19868 27334
rect 19868 27278 19924 27334
rect 19924 27278 19928 27334
rect 19864 27274 19928 27278
rect 50344 27334 50408 27338
rect 50344 27278 50348 27334
rect 50348 27278 50404 27334
rect 50404 27278 50408 27334
rect 50344 27274 50408 27278
rect 50424 27334 50488 27338
rect 50424 27278 50428 27334
rect 50428 27278 50484 27334
rect 50484 27278 50488 27334
rect 50424 27274 50488 27278
rect 50504 27334 50568 27338
rect 50504 27278 50508 27334
rect 50508 27278 50564 27334
rect 50564 27278 50568 27334
rect 50504 27274 50568 27278
rect 50584 27334 50648 27338
rect 50584 27278 50588 27334
rect 50588 27278 50644 27334
rect 50644 27278 50648 27334
rect 50584 27274 50648 27278
rect 4264 26668 4328 26672
rect 4264 26612 4268 26668
rect 4268 26612 4324 26668
rect 4324 26612 4328 26668
rect 4264 26608 4328 26612
rect 4344 26668 4408 26672
rect 4344 26612 4348 26668
rect 4348 26612 4404 26668
rect 4404 26612 4408 26668
rect 4344 26608 4408 26612
rect 4424 26668 4488 26672
rect 4424 26612 4428 26668
rect 4428 26612 4484 26668
rect 4484 26612 4488 26668
rect 4424 26608 4488 26612
rect 4504 26668 4568 26672
rect 4504 26612 4508 26668
rect 4508 26612 4564 26668
rect 4564 26612 4568 26668
rect 4504 26608 4568 26612
rect 34984 26668 35048 26672
rect 34984 26612 34988 26668
rect 34988 26612 35044 26668
rect 35044 26612 35048 26668
rect 34984 26608 35048 26612
rect 35064 26668 35128 26672
rect 35064 26612 35068 26668
rect 35068 26612 35124 26668
rect 35124 26612 35128 26668
rect 35064 26608 35128 26612
rect 35144 26668 35208 26672
rect 35144 26612 35148 26668
rect 35148 26612 35204 26668
rect 35204 26612 35208 26668
rect 35144 26608 35208 26612
rect 35224 26668 35288 26672
rect 35224 26612 35228 26668
rect 35228 26612 35284 26668
rect 35284 26612 35288 26668
rect 35224 26608 35288 26612
rect 19624 26002 19688 26006
rect 19624 25946 19628 26002
rect 19628 25946 19684 26002
rect 19684 25946 19688 26002
rect 19624 25942 19688 25946
rect 19704 26002 19768 26006
rect 19704 25946 19708 26002
rect 19708 25946 19764 26002
rect 19764 25946 19768 26002
rect 19704 25942 19768 25946
rect 19784 26002 19848 26006
rect 19784 25946 19788 26002
rect 19788 25946 19844 26002
rect 19844 25946 19848 26002
rect 19784 25942 19848 25946
rect 19864 26002 19928 26006
rect 19864 25946 19868 26002
rect 19868 25946 19924 26002
rect 19924 25946 19928 26002
rect 19864 25942 19928 25946
rect 50344 26002 50408 26006
rect 50344 25946 50348 26002
rect 50348 25946 50404 26002
rect 50404 25946 50408 26002
rect 50344 25942 50408 25946
rect 50424 26002 50488 26006
rect 50424 25946 50428 26002
rect 50428 25946 50484 26002
rect 50484 25946 50488 26002
rect 50424 25942 50488 25946
rect 50504 26002 50568 26006
rect 50504 25946 50508 26002
rect 50508 25946 50564 26002
rect 50564 25946 50568 26002
rect 50504 25942 50568 25946
rect 50584 26002 50648 26006
rect 50584 25946 50588 26002
rect 50588 25946 50644 26002
rect 50644 25946 50648 26002
rect 50584 25942 50648 25946
rect 4264 25336 4328 25340
rect 4264 25280 4268 25336
rect 4268 25280 4324 25336
rect 4324 25280 4328 25336
rect 4264 25276 4328 25280
rect 4344 25336 4408 25340
rect 4344 25280 4348 25336
rect 4348 25280 4404 25336
rect 4404 25280 4408 25336
rect 4344 25276 4408 25280
rect 4424 25336 4488 25340
rect 4424 25280 4428 25336
rect 4428 25280 4484 25336
rect 4484 25280 4488 25336
rect 4424 25276 4488 25280
rect 4504 25336 4568 25340
rect 4504 25280 4508 25336
rect 4508 25280 4564 25336
rect 4564 25280 4568 25336
rect 4504 25276 4568 25280
rect 34984 25336 35048 25340
rect 34984 25280 34988 25336
rect 34988 25280 35044 25336
rect 35044 25280 35048 25336
rect 34984 25276 35048 25280
rect 35064 25336 35128 25340
rect 35064 25280 35068 25336
rect 35068 25280 35124 25336
rect 35124 25280 35128 25336
rect 35064 25276 35128 25280
rect 35144 25336 35208 25340
rect 35144 25280 35148 25336
rect 35148 25280 35204 25336
rect 35204 25280 35208 25336
rect 35144 25276 35208 25280
rect 35224 25336 35288 25340
rect 35224 25280 35228 25336
rect 35228 25280 35284 25336
rect 35284 25280 35288 25336
rect 35224 25276 35288 25280
rect 19624 24670 19688 24674
rect 19624 24614 19628 24670
rect 19628 24614 19684 24670
rect 19684 24614 19688 24670
rect 19624 24610 19688 24614
rect 19704 24670 19768 24674
rect 19704 24614 19708 24670
rect 19708 24614 19764 24670
rect 19764 24614 19768 24670
rect 19704 24610 19768 24614
rect 19784 24670 19848 24674
rect 19784 24614 19788 24670
rect 19788 24614 19844 24670
rect 19844 24614 19848 24670
rect 19784 24610 19848 24614
rect 19864 24670 19928 24674
rect 19864 24614 19868 24670
rect 19868 24614 19924 24670
rect 19924 24614 19928 24670
rect 19864 24610 19928 24614
rect 50344 24670 50408 24674
rect 50344 24614 50348 24670
rect 50348 24614 50404 24670
rect 50404 24614 50408 24670
rect 50344 24610 50408 24614
rect 50424 24670 50488 24674
rect 50424 24614 50428 24670
rect 50428 24614 50484 24670
rect 50484 24614 50488 24670
rect 50424 24610 50488 24614
rect 50504 24670 50568 24674
rect 50504 24614 50508 24670
rect 50508 24614 50564 24670
rect 50564 24614 50568 24670
rect 50504 24610 50568 24614
rect 50584 24670 50648 24674
rect 50584 24614 50588 24670
rect 50588 24614 50644 24670
rect 50644 24614 50648 24670
rect 50584 24610 50648 24614
rect 4264 24004 4328 24008
rect 4264 23948 4268 24004
rect 4268 23948 4324 24004
rect 4324 23948 4328 24004
rect 4264 23944 4328 23948
rect 4344 24004 4408 24008
rect 4344 23948 4348 24004
rect 4348 23948 4404 24004
rect 4404 23948 4408 24004
rect 4344 23944 4408 23948
rect 4424 24004 4488 24008
rect 4424 23948 4428 24004
rect 4428 23948 4484 24004
rect 4484 23948 4488 24004
rect 4424 23944 4488 23948
rect 4504 24004 4568 24008
rect 4504 23948 4508 24004
rect 4508 23948 4564 24004
rect 4564 23948 4568 24004
rect 4504 23944 4568 23948
rect 34984 24004 35048 24008
rect 34984 23948 34988 24004
rect 34988 23948 35044 24004
rect 35044 23948 35048 24004
rect 34984 23944 35048 23948
rect 35064 24004 35128 24008
rect 35064 23948 35068 24004
rect 35068 23948 35124 24004
rect 35124 23948 35128 24004
rect 35064 23944 35128 23948
rect 35144 24004 35208 24008
rect 35144 23948 35148 24004
rect 35148 23948 35204 24004
rect 35204 23948 35208 24004
rect 35144 23944 35208 23948
rect 35224 24004 35288 24008
rect 35224 23948 35228 24004
rect 35228 23948 35284 24004
rect 35284 23948 35288 24004
rect 35224 23944 35288 23948
rect 19624 23338 19688 23342
rect 19624 23282 19628 23338
rect 19628 23282 19684 23338
rect 19684 23282 19688 23338
rect 19624 23278 19688 23282
rect 19704 23338 19768 23342
rect 19704 23282 19708 23338
rect 19708 23282 19764 23338
rect 19764 23282 19768 23338
rect 19704 23278 19768 23282
rect 19784 23338 19848 23342
rect 19784 23282 19788 23338
rect 19788 23282 19844 23338
rect 19844 23282 19848 23338
rect 19784 23278 19848 23282
rect 19864 23338 19928 23342
rect 19864 23282 19868 23338
rect 19868 23282 19924 23338
rect 19924 23282 19928 23338
rect 19864 23278 19928 23282
rect 50344 23338 50408 23342
rect 50344 23282 50348 23338
rect 50348 23282 50404 23338
rect 50404 23282 50408 23338
rect 50344 23278 50408 23282
rect 50424 23338 50488 23342
rect 50424 23282 50428 23338
rect 50428 23282 50484 23338
rect 50484 23282 50488 23338
rect 50424 23278 50488 23282
rect 50504 23338 50568 23342
rect 50504 23282 50508 23338
rect 50508 23282 50564 23338
rect 50564 23282 50568 23338
rect 50504 23278 50568 23282
rect 50584 23338 50648 23342
rect 50584 23282 50588 23338
rect 50588 23282 50644 23338
rect 50644 23282 50648 23338
rect 50584 23278 50648 23282
rect 4264 22672 4328 22676
rect 4264 22616 4268 22672
rect 4268 22616 4324 22672
rect 4324 22616 4328 22672
rect 4264 22612 4328 22616
rect 4344 22672 4408 22676
rect 4344 22616 4348 22672
rect 4348 22616 4404 22672
rect 4404 22616 4408 22672
rect 4344 22612 4408 22616
rect 4424 22672 4488 22676
rect 4424 22616 4428 22672
rect 4428 22616 4484 22672
rect 4484 22616 4488 22672
rect 4424 22612 4488 22616
rect 4504 22672 4568 22676
rect 4504 22616 4508 22672
rect 4508 22616 4564 22672
rect 4564 22616 4568 22672
rect 4504 22612 4568 22616
rect 34984 22672 35048 22676
rect 34984 22616 34988 22672
rect 34988 22616 35044 22672
rect 35044 22616 35048 22672
rect 34984 22612 35048 22616
rect 35064 22672 35128 22676
rect 35064 22616 35068 22672
rect 35068 22616 35124 22672
rect 35124 22616 35128 22672
rect 35064 22612 35128 22616
rect 35144 22672 35208 22676
rect 35144 22616 35148 22672
rect 35148 22616 35204 22672
rect 35204 22616 35208 22672
rect 35144 22612 35208 22616
rect 35224 22672 35288 22676
rect 35224 22616 35228 22672
rect 35228 22616 35284 22672
rect 35284 22616 35288 22672
rect 35224 22612 35288 22616
rect 19624 22006 19688 22010
rect 19624 21950 19628 22006
rect 19628 21950 19684 22006
rect 19684 21950 19688 22006
rect 19624 21946 19688 21950
rect 19704 22006 19768 22010
rect 19704 21950 19708 22006
rect 19708 21950 19764 22006
rect 19764 21950 19768 22006
rect 19704 21946 19768 21950
rect 19784 22006 19848 22010
rect 19784 21950 19788 22006
rect 19788 21950 19844 22006
rect 19844 21950 19848 22006
rect 19784 21946 19848 21950
rect 19864 22006 19928 22010
rect 19864 21950 19868 22006
rect 19868 21950 19924 22006
rect 19924 21950 19928 22006
rect 19864 21946 19928 21950
rect 50344 22006 50408 22010
rect 50344 21950 50348 22006
rect 50348 21950 50404 22006
rect 50404 21950 50408 22006
rect 50344 21946 50408 21950
rect 50424 22006 50488 22010
rect 50424 21950 50428 22006
rect 50428 21950 50484 22006
rect 50484 21950 50488 22006
rect 50424 21946 50488 21950
rect 50504 22006 50568 22010
rect 50504 21950 50508 22006
rect 50508 21950 50564 22006
rect 50564 21950 50568 22006
rect 50504 21946 50568 21950
rect 50584 22006 50648 22010
rect 50584 21950 50588 22006
rect 50588 21950 50644 22006
rect 50644 21950 50648 22006
rect 50584 21946 50648 21950
rect 4264 21340 4328 21344
rect 4264 21284 4268 21340
rect 4268 21284 4324 21340
rect 4324 21284 4328 21340
rect 4264 21280 4328 21284
rect 4344 21340 4408 21344
rect 4344 21284 4348 21340
rect 4348 21284 4404 21340
rect 4404 21284 4408 21340
rect 4344 21280 4408 21284
rect 4424 21340 4488 21344
rect 4424 21284 4428 21340
rect 4428 21284 4484 21340
rect 4484 21284 4488 21340
rect 4424 21280 4488 21284
rect 4504 21340 4568 21344
rect 4504 21284 4508 21340
rect 4508 21284 4564 21340
rect 4564 21284 4568 21340
rect 4504 21280 4568 21284
rect 34984 21340 35048 21344
rect 34984 21284 34988 21340
rect 34988 21284 35044 21340
rect 35044 21284 35048 21340
rect 34984 21280 35048 21284
rect 35064 21340 35128 21344
rect 35064 21284 35068 21340
rect 35068 21284 35124 21340
rect 35124 21284 35128 21340
rect 35064 21280 35128 21284
rect 35144 21340 35208 21344
rect 35144 21284 35148 21340
rect 35148 21284 35204 21340
rect 35204 21284 35208 21340
rect 35144 21280 35208 21284
rect 35224 21340 35288 21344
rect 35224 21284 35228 21340
rect 35228 21284 35284 21340
rect 35284 21284 35288 21340
rect 35224 21280 35288 21284
rect 19624 20674 19688 20678
rect 19624 20618 19628 20674
rect 19628 20618 19684 20674
rect 19684 20618 19688 20674
rect 19624 20614 19688 20618
rect 19704 20674 19768 20678
rect 19704 20618 19708 20674
rect 19708 20618 19764 20674
rect 19764 20618 19768 20674
rect 19704 20614 19768 20618
rect 19784 20674 19848 20678
rect 19784 20618 19788 20674
rect 19788 20618 19844 20674
rect 19844 20618 19848 20674
rect 19784 20614 19848 20618
rect 19864 20674 19928 20678
rect 19864 20618 19868 20674
rect 19868 20618 19924 20674
rect 19924 20618 19928 20674
rect 19864 20614 19928 20618
rect 50344 20674 50408 20678
rect 50344 20618 50348 20674
rect 50348 20618 50404 20674
rect 50404 20618 50408 20674
rect 50344 20614 50408 20618
rect 50424 20674 50488 20678
rect 50424 20618 50428 20674
rect 50428 20618 50484 20674
rect 50484 20618 50488 20674
rect 50424 20614 50488 20618
rect 50504 20674 50568 20678
rect 50504 20618 50508 20674
rect 50508 20618 50564 20674
rect 50564 20618 50568 20674
rect 50504 20614 50568 20618
rect 50584 20674 50648 20678
rect 50584 20618 50588 20674
rect 50588 20618 50644 20674
rect 50644 20618 50648 20674
rect 50584 20614 50648 20618
rect 4264 20008 4328 20012
rect 4264 19952 4268 20008
rect 4268 19952 4324 20008
rect 4324 19952 4328 20008
rect 4264 19948 4328 19952
rect 4344 20008 4408 20012
rect 4344 19952 4348 20008
rect 4348 19952 4404 20008
rect 4404 19952 4408 20008
rect 4344 19948 4408 19952
rect 4424 20008 4488 20012
rect 4424 19952 4428 20008
rect 4428 19952 4484 20008
rect 4484 19952 4488 20008
rect 4424 19948 4488 19952
rect 4504 20008 4568 20012
rect 4504 19952 4508 20008
rect 4508 19952 4564 20008
rect 4564 19952 4568 20008
rect 4504 19948 4568 19952
rect 34984 20008 35048 20012
rect 34984 19952 34988 20008
rect 34988 19952 35044 20008
rect 35044 19952 35048 20008
rect 34984 19948 35048 19952
rect 35064 20008 35128 20012
rect 35064 19952 35068 20008
rect 35068 19952 35124 20008
rect 35124 19952 35128 20008
rect 35064 19948 35128 19952
rect 35144 20008 35208 20012
rect 35144 19952 35148 20008
rect 35148 19952 35204 20008
rect 35204 19952 35208 20008
rect 35144 19948 35208 19952
rect 35224 20008 35288 20012
rect 35224 19952 35228 20008
rect 35228 19952 35284 20008
rect 35284 19952 35288 20008
rect 35224 19948 35288 19952
rect 19624 19342 19688 19346
rect 19624 19286 19628 19342
rect 19628 19286 19684 19342
rect 19684 19286 19688 19342
rect 19624 19282 19688 19286
rect 19704 19342 19768 19346
rect 19704 19286 19708 19342
rect 19708 19286 19764 19342
rect 19764 19286 19768 19342
rect 19704 19282 19768 19286
rect 19784 19342 19848 19346
rect 19784 19286 19788 19342
rect 19788 19286 19844 19342
rect 19844 19286 19848 19342
rect 19784 19282 19848 19286
rect 19864 19342 19928 19346
rect 19864 19286 19868 19342
rect 19868 19286 19924 19342
rect 19924 19286 19928 19342
rect 19864 19282 19928 19286
rect 50344 19342 50408 19346
rect 50344 19286 50348 19342
rect 50348 19286 50404 19342
rect 50404 19286 50408 19342
rect 50344 19282 50408 19286
rect 50424 19342 50488 19346
rect 50424 19286 50428 19342
rect 50428 19286 50484 19342
rect 50484 19286 50488 19342
rect 50424 19282 50488 19286
rect 50504 19342 50568 19346
rect 50504 19286 50508 19342
rect 50508 19286 50564 19342
rect 50564 19286 50568 19342
rect 50504 19282 50568 19286
rect 50584 19342 50648 19346
rect 50584 19286 50588 19342
rect 50588 19286 50644 19342
rect 50644 19286 50648 19342
rect 50584 19282 50648 19286
rect 4264 18676 4328 18680
rect 4264 18620 4268 18676
rect 4268 18620 4324 18676
rect 4324 18620 4328 18676
rect 4264 18616 4328 18620
rect 4344 18676 4408 18680
rect 4344 18620 4348 18676
rect 4348 18620 4404 18676
rect 4404 18620 4408 18676
rect 4344 18616 4408 18620
rect 4424 18676 4488 18680
rect 4424 18620 4428 18676
rect 4428 18620 4484 18676
rect 4484 18620 4488 18676
rect 4424 18616 4488 18620
rect 4504 18676 4568 18680
rect 4504 18620 4508 18676
rect 4508 18620 4564 18676
rect 4564 18620 4568 18676
rect 4504 18616 4568 18620
rect 34984 18676 35048 18680
rect 34984 18620 34988 18676
rect 34988 18620 35044 18676
rect 35044 18620 35048 18676
rect 34984 18616 35048 18620
rect 35064 18676 35128 18680
rect 35064 18620 35068 18676
rect 35068 18620 35124 18676
rect 35124 18620 35128 18676
rect 35064 18616 35128 18620
rect 35144 18676 35208 18680
rect 35144 18620 35148 18676
rect 35148 18620 35204 18676
rect 35204 18620 35208 18676
rect 35144 18616 35208 18620
rect 35224 18676 35288 18680
rect 35224 18620 35228 18676
rect 35228 18620 35284 18676
rect 35284 18620 35288 18676
rect 35224 18616 35288 18620
rect 19624 18010 19688 18014
rect 19624 17954 19628 18010
rect 19628 17954 19684 18010
rect 19684 17954 19688 18010
rect 19624 17950 19688 17954
rect 19704 18010 19768 18014
rect 19704 17954 19708 18010
rect 19708 17954 19764 18010
rect 19764 17954 19768 18010
rect 19704 17950 19768 17954
rect 19784 18010 19848 18014
rect 19784 17954 19788 18010
rect 19788 17954 19844 18010
rect 19844 17954 19848 18010
rect 19784 17950 19848 17954
rect 19864 18010 19928 18014
rect 19864 17954 19868 18010
rect 19868 17954 19924 18010
rect 19924 17954 19928 18010
rect 19864 17950 19928 17954
rect 50344 18010 50408 18014
rect 50344 17954 50348 18010
rect 50348 17954 50404 18010
rect 50404 17954 50408 18010
rect 50344 17950 50408 17954
rect 50424 18010 50488 18014
rect 50424 17954 50428 18010
rect 50428 17954 50484 18010
rect 50484 17954 50488 18010
rect 50424 17950 50488 17954
rect 50504 18010 50568 18014
rect 50504 17954 50508 18010
rect 50508 17954 50564 18010
rect 50564 17954 50568 18010
rect 50504 17950 50568 17954
rect 50584 18010 50648 18014
rect 50584 17954 50588 18010
rect 50588 17954 50644 18010
rect 50644 17954 50648 18010
rect 50584 17950 50648 17954
rect 4264 17344 4328 17348
rect 4264 17288 4268 17344
rect 4268 17288 4324 17344
rect 4324 17288 4328 17344
rect 4264 17284 4328 17288
rect 4344 17344 4408 17348
rect 4344 17288 4348 17344
rect 4348 17288 4404 17344
rect 4404 17288 4408 17344
rect 4344 17284 4408 17288
rect 4424 17344 4488 17348
rect 4424 17288 4428 17344
rect 4428 17288 4484 17344
rect 4484 17288 4488 17344
rect 4424 17284 4488 17288
rect 4504 17344 4568 17348
rect 4504 17288 4508 17344
rect 4508 17288 4564 17344
rect 4564 17288 4568 17344
rect 4504 17284 4568 17288
rect 34984 17344 35048 17348
rect 34984 17288 34988 17344
rect 34988 17288 35044 17344
rect 35044 17288 35048 17344
rect 34984 17284 35048 17288
rect 35064 17344 35128 17348
rect 35064 17288 35068 17344
rect 35068 17288 35124 17344
rect 35124 17288 35128 17344
rect 35064 17284 35128 17288
rect 35144 17344 35208 17348
rect 35144 17288 35148 17344
rect 35148 17288 35204 17344
rect 35204 17288 35208 17344
rect 35144 17284 35208 17288
rect 35224 17344 35288 17348
rect 35224 17288 35228 17344
rect 35228 17288 35284 17344
rect 35284 17288 35288 17344
rect 35224 17284 35288 17288
rect 19624 16678 19688 16682
rect 19624 16622 19628 16678
rect 19628 16622 19684 16678
rect 19684 16622 19688 16678
rect 19624 16618 19688 16622
rect 19704 16678 19768 16682
rect 19704 16622 19708 16678
rect 19708 16622 19764 16678
rect 19764 16622 19768 16678
rect 19704 16618 19768 16622
rect 19784 16678 19848 16682
rect 19784 16622 19788 16678
rect 19788 16622 19844 16678
rect 19844 16622 19848 16678
rect 19784 16618 19848 16622
rect 19864 16678 19928 16682
rect 19864 16622 19868 16678
rect 19868 16622 19924 16678
rect 19924 16622 19928 16678
rect 19864 16618 19928 16622
rect 50344 16678 50408 16682
rect 50344 16622 50348 16678
rect 50348 16622 50404 16678
rect 50404 16622 50408 16678
rect 50344 16618 50408 16622
rect 50424 16678 50488 16682
rect 50424 16622 50428 16678
rect 50428 16622 50484 16678
rect 50484 16622 50488 16678
rect 50424 16618 50488 16622
rect 50504 16678 50568 16682
rect 50504 16622 50508 16678
rect 50508 16622 50564 16678
rect 50564 16622 50568 16678
rect 50504 16618 50568 16622
rect 50584 16678 50648 16682
rect 50584 16622 50588 16678
rect 50588 16622 50644 16678
rect 50644 16622 50648 16678
rect 50584 16618 50648 16622
rect 4264 16012 4328 16016
rect 4264 15956 4268 16012
rect 4268 15956 4324 16012
rect 4324 15956 4328 16012
rect 4264 15952 4328 15956
rect 4344 16012 4408 16016
rect 4344 15956 4348 16012
rect 4348 15956 4404 16012
rect 4404 15956 4408 16012
rect 4344 15952 4408 15956
rect 4424 16012 4488 16016
rect 4424 15956 4428 16012
rect 4428 15956 4484 16012
rect 4484 15956 4488 16012
rect 4424 15952 4488 15956
rect 4504 16012 4568 16016
rect 4504 15956 4508 16012
rect 4508 15956 4564 16012
rect 4564 15956 4568 16012
rect 4504 15952 4568 15956
rect 34984 16012 35048 16016
rect 34984 15956 34988 16012
rect 34988 15956 35044 16012
rect 35044 15956 35048 16012
rect 34984 15952 35048 15956
rect 35064 16012 35128 16016
rect 35064 15956 35068 16012
rect 35068 15956 35124 16012
rect 35124 15956 35128 16012
rect 35064 15952 35128 15956
rect 35144 16012 35208 16016
rect 35144 15956 35148 16012
rect 35148 15956 35204 16012
rect 35204 15956 35208 16012
rect 35144 15952 35208 15956
rect 35224 16012 35288 16016
rect 35224 15956 35228 16012
rect 35228 15956 35284 16012
rect 35284 15956 35288 16012
rect 35224 15952 35288 15956
rect 19624 15346 19688 15350
rect 19624 15290 19628 15346
rect 19628 15290 19684 15346
rect 19684 15290 19688 15346
rect 19624 15286 19688 15290
rect 19704 15346 19768 15350
rect 19704 15290 19708 15346
rect 19708 15290 19764 15346
rect 19764 15290 19768 15346
rect 19704 15286 19768 15290
rect 19784 15346 19848 15350
rect 19784 15290 19788 15346
rect 19788 15290 19844 15346
rect 19844 15290 19848 15346
rect 19784 15286 19848 15290
rect 19864 15346 19928 15350
rect 19864 15290 19868 15346
rect 19868 15290 19924 15346
rect 19924 15290 19928 15346
rect 19864 15286 19928 15290
rect 50344 15346 50408 15350
rect 50344 15290 50348 15346
rect 50348 15290 50404 15346
rect 50404 15290 50408 15346
rect 50344 15286 50408 15290
rect 50424 15346 50488 15350
rect 50424 15290 50428 15346
rect 50428 15290 50484 15346
rect 50484 15290 50488 15346
rect 50424 15286 50488 15290
rect 50504 15346 50568 15350
rect 50504 15290 50508 15346
rect 50508 15290 50564 15346
rect 50564 15290 50568 15346
rect 50504 15286 50568 15290
rect 50584 15346 50648 15350
rect 50584 15290 50588 15346
rect 50588 15290 50644 15346
rect 50644 15290 50648 15346
rect 50584 15286 50648 15290
rect 4264 14680 4328 14684
rect 4264 14624 4268 14680
rect 4268 14624 4324 14680
rect 4324 14624 4328 14680
rect 4264 14620 4328 14624
rect 4344 14680 4408 14684
rect 4344 14624 4348 14680
rect 4348 14624 4404 14680
rect 4404 14624 4408 14680
rect 4344 14620 4408 14624
rect 4424 14680 4488 14684
rect 4424 14624 4428 14680
rect 4428 14624 4484 14680
rect 4484 14624 4488 14680
rect 4424 14620 4488 14624
rect 4504 14680 4568 14684
rect 4504 14624 4508 14680
rect 4508 14624 4564 14680
rect 4564 14624 4568 14680
rect 4504 14620 4568 14624
rect 34984 14680 35048 14684
rect 34984 14624 34988 14680
rect 34988 14624 35044 14680
rect 35044 14624 35048 14680
rect 34984 14620 35048 14624
rect 35064 14680 35128 14684
rect 35064 14624 35068 14680
rect 35068 14624 35124 14680
rect 35124 14624 35128 14680
rect 35064 14620 35128 14624
rect 35144 14680 35208 14684
rect 35144 14624 35148 14680
rect 35148 14624 35204 14680
rect 35204 14624 35208 14680
rect 35144 14620 35208 14624
rect 35224 14680 35288 14684
rect 35224 14624 35228 14680
rect 35228 14624 35284 14680
rect 35284 14624 35288 14680
rect 35224 14620 35288 14624
rect 19624 14014 19688 14018
rect 19624 13958 19628 14014
rect 19628 13958 19684 14014
rect 19684 13958 19688 14014
rect 19624 13954 19688 13958
rect 19704 14014 19768 14018
rect 19704 13958 19708 14014
rect 19708 13958 19764 14014
rect 19764 13958 19768 14014
rect 19704 13954 19768 13958
rect 19784 14014 19848 14018
rect 19784 13958 19788 14014
rect 19788 13958 19844 14014
rect 19844 13958 19848 14014
rect 19784 13954 19848 13958
rect 19864 14014 19928 14018
rect 19864 13958 19868 14014
rect 19868 13958 19924 14014
rect 19924 13958 19928 14014
rect 19864 13954 19928 13958
rect 50344 14014 50408 14018
rect 50344 13958 50348 14014
rect 50348 13958 50404 14014
rect 50404 13958 50408 14014
rect 50344 13954 50408 13958
rect 50424 14014 50488 14018
rect 50424 13958 50428 14014
rect 50428 13958 50484 14014
rect 50484 13958 50488 14014
rect 50424 13954 50488 13958
rect 50504 14014 50568 14018
rect 50504 13958 50508 14014
rect 50508 13958 50564 14014
rect 50564 13958 50568 14014
rect 50504 13954 50568 13958
rect 50584 14014 50648 14018
rect 50584 13958 50588 14014
rect 50588 13958 50644 14014
rect 50644 13958 50648 14014
rect 50584 13954 50648 13958
rect 4264 13348 4328 13352
rect 4264 13292 4268 13348
rect 4268 13292 4324 13348
rect 4324 13292 4328 13348
rect 4264 13288 4328 13292
rect 4344 13348 4408 13352
rect 4344 13292 4348 13348
rect 4348 13292 4404 13348
rect 4404 13292 4408 13348
rect 4344 13288 4408 13292
rect 4424 13348 4488 13352
rect 4424 13292 4428 13348
rect 4428 13292 4484 13348
rect 4484 13292 4488 13348
rect 4424 13288 4488 13292
rect 4504 13348 4568 13352
rect 4504 13292 4508 13348
rect 4508 13292 4564 13348
rect 4564 13292 4568 13348
rect 4504 13288 4568 13292
rect 34984 13348 35048 13352
rect 34984 13292 34988 13348
rect 34988 13292 35044 13348
rect 35044 13292 35048 13348
rect 34984 13288 35048 13292
rect 35064 13348 35128 13352
rect 35064 13292 35068 13348
rect 35068 13292 35124 13348
rect 35124 13292 35128 13348
rect 35064 13288 35128 13292
rect 35144 13348 35208 13352
rect 35144 13292 35148 13348
rect 35148 13292 35204 13348
rect 35204 13292 35208 13348
rect 35144 13288 35208 13292
rect 35224 13348 35288 13352
rect 35224 13292 35228 13348
rect 35228 13292 35284 13348
rect 35284 13292 35288 13348
rect 35224 13288 35288 13292
rect 19624 12682 19688 12686
rect 19624 12626 19628 12682
rect 19628 12626 19684 12682
rect 19684 12626 19688 12682
rect 19624 12622 19688 12626
rect 19704 12682 19768 12686
rect 19704 12626 19708 12682
rect 19708 12626 19764 12682
rect 19764 12626 19768 12682
rect 19704 12622 19768 12626
rect 19784 12682 19848 12686
rect 19784 12626 19788 12682
rect 19788 12626 19844 12682
rect 19844 12626 19848 12682
rect 19784 12622 19848 12626
rect 19864 12682 19928 12686
rect 19864 12626 19868 12682
rect 19868 12626 19924 12682
rect 19924 12626 19928 12682
rect 19864 12622 19928 12626
rect 50344 12682 50408 12686
rect 50344 12626 50348 12682
rect 50348 12626 50404 12682
rect 50404 12626 50408 12682
rect 50344 12622 50408 12626
rect 50424 12682 50488 12686
rect 50424 12626 50428 12682
rect 50428 12626 50484 12682
rect 50484 12626 50488 12682
rect 50424 12622 50488 12626
rect 50504 12682 50568 12686
rect 50504 12626 50508 12682
rect 50508 12626 50564 12682
rect 50564 12626 50568 12682
rect 50504 12622 50568 12626
rect 50584 12682 50648 12686
rect 50584 12626 50588 12682
rect 50588 12626 50644 12682
rect 50644 12626 50648 12682
rect 50584 12622 50648 12626
rect 4264 12016 4328 12020
rect 4264 11960 4268 12016
rect 4268 11960 4324 12016
rect 4324 11960 4328 12016
rect 4264 11956 4328 11960
rect 4344 12016 4408 12020
rect 4344 11960 4348 12016
rect 4348 11960 4404 12016
rect 4404 11960 4408 12016
rect 4344 11956 4408 11960
rect 4424 12016 4488 12020
rect 4424 11960 4428 12016
rect 4428 11960 4484 12016
rect 4484 11960 4488 12016
rect 4424 11956 4488 11960
rect 4504 12016 4568 12020
rect 4504 11960 4508 12016
rect 4508 11960 4564 12016
rect 4564 11960 4568 12016
rect 4504 11956 4568 11960
rect 34984 12016 35048 12020
rect 34984 11960 34988 12016
rect 34988 11960 35044 12016
rect 35044 11960 35048 12016
rect 34984 11956 35048 11960
rect 35064 12016 35128 12020
rect 35064 11960 35068 12016
rect 35068 11960 35124 12016
rect 35124 11960 35128 12016
rect 35064 11956 35128 11960
rect 35144 12016 35208 12020
rect 35144 11960 35148 12016
rect 35148 11960 35204 12016
rect 35204 11960 35208 12016
rect 35144 11956 35208 11960
rect 35224 12016 35288 12020
rect 35224 11960 35228 12016
rect 35228 11960 35284 12016
rect 35284 11960 35288 12016
rect 35224 11956 35288 11960
rect 19624 11350 19688 11354
rect 19624 11294 19628 11350
rect 19628 11294 19684 11350
rect 19684 11294 19688 11350
rect 19624 11290 19688 11294
rect 19704 11350 19768 11354
rect 19704 11294 19708 11350
rect 19708 11294 19764 11350
rect 19764 11294 19768 11350
rect 19704 11290 19768 11294
rect 19784 11350 19848 11354
rect 19784 11294 19788 11350
rect 19788 11294 19844 11350
rect 19844 11294 19848 11350
rect 19784 11290 19848 11294
rect 19864 11350 19928 11354
rect 19864 11294 19868 11350
rect 19868 11294 19924 11350
rect 19924 11294 19928 11350
rect 19864 11290 19928 11294
rect 50344 11350 50408 11354
rect 50344 11294 50348 11350
rect 50348 11294 50404 11350
rect 50404 11294 50408 11350
rect 50344 11290 50408 11294
rect 50424 11350 50488 11354
rect 50424 11294 50428 11350
rect 50428 11294 50484 11350
rect 50484 11294 50488 11350
rect 50424 11290 50488 11294
rect 50504 11350 50568 11354
rect 50504 11294 50508 11350
rect 50508 11294 50564 11350
rect 50564 11294 50568 11350
rect 50504 11290 50568 11294
rect 50584 11350 50648 11354
rect 50584 11294 50588 11350
rect 50588 11294 50644 11350
rect 50644 11294 50648 11350
rect 50584 11290 50648 11294
rect 4264 10684 4328 10688
rect 4264 10628 4268 10684
rect 4268 10628 4324 10684
rect 4324 10628 4328 10684
rect 4264 10624 4328 10628
rect 4344 10684 4408 10688
rect 4344 10628 4348 10684
rect 4348 10628 4404 10684
rect 4404 10628 4408 10684
rect 4344 10624 4408 10628
rect 4424 10684 4488 10688
rect 4424 10628 4428 10684
rect 4428 10628 4484 10684
rect 4484 10628 4488 10684
rect 4424 10624 4488 10628
rect 4504 10684 4568 10688
rect 4504 10628 4508 10684
rect 4508 10628 4564 10684
rect 4564 10628 4568 10684
rect 4504 10624 4568 10628
rect 34984 10684 35048 10688
rect 34984 10628 34988 10684
rect 34988 10628 35044 10684
rect 35044 10628 35048 10684
rect 34984 10624 35048 10628
rect 35064 10684 35128 10688
rect 35064 10628 35068 10684
rect 35068 10628 35124 10684
rect 35124 10628 35128 10684
rect 35064 10624 35128 10628
rect 35144 10684 35208 10688
rect 35144 10628 35148 10684
rect 35148 10628 35204 10684
rect 35204 10628 35208 10684
rect 35144 10624 35208 10628
rect 35224 10684 35288 10688
rect 35224 10628 35228 10684
rect 35228 10628 35284 10684
rect 35284 10628 35288 10684
rect 35224 10624 35288 10628
rect 19624 10018 19688 10022
rect 19624 9962 19628 10018
rect 19628 9962 19684 10018
rect 19684 9962 19688 10018
rect 19624 9958 19688 9962
rect 19704 10018 19768 10022
rect 19704 9962 19708 10018
rect 19708 9962 19764 10018
rect 19764 9962 19768 10018
rect 19704 9958 19768 9962
rect 19784 10018 19848 10022
rect 19784 9962 19788 10018
rect 19788 9962 19844 10018
rect 19844 9962 19848 10018
rect 19784 9958 19848 9962
rect 19864 10018 19928 10022
rect 19864 9962 19868 10018
rect 19868 9962 19924 10018
rect 19924 9962 19928 10018
rect 19864 9958 19928 9962
rect 50344 10018 50408 10022
rect 50344 9962 50348 10018
rect 50348 9962 50404 10018
rect 50404 9962 50408 10018
rect 50344 9958 50408 9962
rect 50424 10018 50488 10022
rect 50424 9962 50428 10018
rect 50428 9962 50484 10018
rect 50484 9962 50488 10018
rect 50424 9958 50488 9962
rect 50504 10018 50568 10022
rect 50504 9962 50508 10018
rect 50508 9962 50564 10018
rect 50564 9962 50568 10018
rect 50504 9958 50568 9962
rect 50584 10018 50648 10022
rect 50584 9962 50588 10018
rect 50588 9962 50644 10018
rect 50644 9962 50648 10018
rect 50584 9958 50648 9962
rect 4264 9352 4328 9356
rect 4264 9296 4268 9352
rect 4268 9296 4324 9352
rect 4324 9296 4328 9352
rect 4264 9292 4328 9296
rect 4344 9352 4408 9356
rect 4344 9296 4348 9352
rect 4348 9296 4404 9352
rect 4404 9296 4408 9352
rect 4344 9292 4408 9296
rect 4424 9352 4488 9356
rect 4424 9296 4428 9352
rect 4428 9296 4484 9352
rect 4484 9296 4488 9352
rect 4424 9292 4488 9296
rect 4504 9352 4568 9356
rect 4504 9296 4508 9352
rect 4508 9296 4564 9352
rect 4564 9296 4568 9352
rect 4504 9292 4568 9296
rect 34984 9352 35048 9356
rect 34984 9296 34988 9352
rect 34988 9296 35044 9352
rect 35044 9296 35048 9352
rect 34984 9292 35048 9296
rect 35064 9352 35128 9356
rect 35064 9296 35068 9352
rect 35068 9296 35124 9352
rect 35124 9296 35128 9352
rect 35064 9292 35128 9296
rect 35144 9352 35208 9356
rect 35144 9296 35148 9352
rect 35148 9296 35204 9352
rect 35204 9296 35208 9352
rect 35144 9292 35208 9296
rect 35224 9352 35288 9356
rect 35224 9296 35228 9352
rect 35228 9296 35284 9352
rect 35284 9296 35288 9352
rect 35224 9292 35288 9296
rect 19624 8686 19688 8690
rect 19624 8630 19628 8686
rect 19628 8630 19684 8686
rect 19684 8630 19688 8686
rect 19624 8626 19688 8630
rect 19704 8686 19768 8690
rect 19704 8630 19708 8686
rect 19708 8630 19764 8686
rect 19764 8630 19768 8686
rect 19704 8626 19768 8630
rect 19784 8686 19848 8690
rect 19784 8630 19788 8686
rect 19788 8630 19844 8686
rect 19844 8630 19848 8686
rect 19784 8626 19848 8630
rect 19864 8686 19928 8690
rect 19864 8630 19868 8686
rect 19868 8630 19924 8686
rect 19924 8630 19928 8686
rect 19864 8626 19928 8630
rect 50344 8686 50408 8690
rect 50344 8630 50348 8686
rect 50348 8630 50404 8686
rect 50404 8630 50408 8686
rect 50344 8626 50408 8630
rect 50424 8686 50488 8690
rect 50424 8630 50428 8686
rect 50428 8630 50484 8686
rect 50484 8630 50488 8686
rect 50424 8626 50488 8630
rect 50504 8686 50568 8690
rect 50504 8630 50508 8686
rect 50508 8630 50564 8686
rect 50564 8630 50568 8686
rect 50504 8626 50568 8630
rect 50584 8686 50648 8690
rect 50584 8630 50588 8686
rect 50588 8630 50644 8686
rect 50644 8630 50648 8686
rect 50584 8626 50648 8630
rect 4264 8020 4328 8024
rect 4264 7964 4268 8020
rect 4268 7964 4324 8020
rect 4324 7964 4328 8020
rect 4264 7960 4328 7964
rect 4344 8020 4408 8024
rect 4344 7964 4348 8020
rect 4348 7964 4404 8020
rect 4404 7964 4408 8020
rect 4344 7960 4408 7964
rect 4424 8020 4488 8024
rect 4424 7964 4428 8020
rect 4428 7964 4484 8020
rect 4484 7964 4488 8020
rect 4424 7960 4488 7964
rect 4504 8020 4568 8024
rect 4504 7964 4508 8020
rect 4508 7964 4564 8020
rect 4564 7964 4568 8020
rect 4504 7960 4568 7964
rect 34984 8020 35048 8024
rect 34984 7964 34988 8020
rect 34988 7964 35044 8020
rect 35044 7964 35048 8020
rect 34984 7960 35048 7964
rect 35064 8020 35128 8024
rect 35064 7964 35068 8020
rect 35068 7964 35124 8020
rect 35124 7964 35128 8020
rect 35064 7960 35128 7964
rect 35144 8020 35208 8024
rect 35144 7964 35148 8020
rect 35148 7964 35204 8020
rect 35204 7964 35208 8020
rect 35144 7960 35208 7964
rect 35224 8020 35288 8024
rect 35224 7964 35228 8020
rect 35228 7964 35284 8020
rect 35284 7964 35288 8020
rect 35224 7960 35288 7964
rect 19624 7354 19688 7358
rect 19624 7298 19628 7354
rect 19628 7298 19684 7354
rect 19684 7298 19688 7354
rect 19624 7294 19688 7298
rect 19704 7354 19768 7358
rect 19704 7298 19708 7354
rect 19708 7298 19764 7354
rect 19764 7298 19768 7354
rect 19704 7294 19768 7298
rect 19784 7354 19848 7358
rect 19784 7298 19788 7354
rect 19788 7298 19844 7354
rect 19844 7298 19848 7354
rect 19784 7294 19848 7298
rect 19864 7354 19928 7358
rect 19864 7298 19868 7354
rect 19868 7298 19924 7354
rect 19924 7298 19928 7354
rect 19864 7294 19928 7298
rect 50344 7354 50408 7358
rect 50344 7298 50348 7354
rect 50348 7298 50404 7354
rect 50404 7298 50408 7354
rect 50344 7294 50408 7298
rect 50424 7354 50488 7358
rect 50424 7298 50428 7354
rect 50428 7298 50484 7354
rect 50484 7298 50488 7354
rect 50424 7294 50488 7298
rect 50504 7354 50568 7358
rect 50504 7298 50508 7354
rect 50508 7298 50564 7354
rect 50564 7298 50568 7354
rect 50504 7294 50568 7298
rect 50584 7354 50648 7358
rect 50584 7298 50588 7354
rect 50588 7298 50644 7354
rect 50644 7298 50648 7354
rect 50584 7294 50648 7298
rect 4264 6688 4328 6692
rect 4264 6632 4268 6688
rect 4268 6632 4324 6688
rect 4324 6632 4328 6688
rect 4264 6628 4328 6632
rect 4344 6688 4408 6692
rect 4344 6632 4348 6688
rect 4348 6632 4404 6688
rect 4404 6632 4408 6688
rect 4344 6628 4408 6632
rect 4424 6688 4488 6692
rect 4424 6632 4428 6688
rect 4428 6632 4484 6688
rect 4484 6632 4488 6688
rect 4424 6628 4488 6632
rect 4504 6688 4568 6692
rect 4504 6632 4508 6688
rect 4508 6632 4564 6688
rect 4564 6632 4568 6688
rect 4504 6628 4568 6632
rect 34984 6688 35048 6692
rect 34984 6632 34988 6688
rect 34988 6632 35044 6688
rect 35044 6632 35048 6688
rect 34984 6628 35048 6632
rect 35064 6688 35128 6692
rect 35064 6632 35068 6688
rect 35068 6632 35124 6688
rect 35124 6632 35128 6688
rect 35064 6628 35128 6632
rect 35144 6688 35208 6692
rect 35144 6632 35148 6688
rect 35148 6632 35204 6688
rect 35204 6632 35208 6688
rect 35144 6628 35208 6632
rect 35224 6688 35288 6692
rect 35224 6632 35228 6688
rect 35228 6632 35284 6688
rect 35284 6632 35288 6688
rect 35224 6628 35288 6632
rect 19624 6022 19688 6026
rect 19624 5966 19628 6022
rect 19628 5966 19684 6022
rect 19684 5966 19688 6022
rect 19624 5962 19688 5966
rect 19704 6022 19768 6026
rect 19704 5966 19708 6022
rect 19708 5966 19764 6022
rect 19764 5966 19768 6022
rect 19704 5962 19768 5966
rect 19784 6022 19848 6026
rect 19784 5966 19788 6022
rect 19788 5966 19844 6022
rect 19844 5966 19848 6022
rect 19784 5962 19848 5966
rect 19864 6022 19928 6026
rect 19864 5966 19868 6022
rect 19868 5966 19924 6022
rect 19924 5966 19928 6022
rect 19864 5962 19928 5966
rect 50344 6022 50408 6026
rect 50344 5966 50348 6022
rect 50348 5966 50404 6022
rect 50404 5966 50408 6022
rect 50344 5962 50408 5966
rect 50424 6022 50488 6026
rect 50424 5966 50428 6022
rect 50428 5966 50484 6022
rect 50484 5966 50488 6022
rect 50424 5962 50488 5966
rect 50504 6022 50568 6026
rect 50504 5966 50508 6022
rect 50508 5966 50564 6022
rect 50564 5966 50568 6022
rect 50504 5962 50568 5966
rect 50584 6022 50648 6026
rect 50584 5966 50588 6022
rect 50588 5966 50644 6022
rect 50644 5966 50648 6022
rect 50584 5962 50648 5966
rect 4264 5356 4328 5360
rect 4264 5300 4268 5356
rect 4268 5300 4324 5356
rect 4324 5300 4328 5356
rect 4264 5296 4328 5300
rect 4344 5356 4408 5360
rect 4344 5300 4348 5356
rect 4348 5300 4404 5356
rect 4404 5300 4408 5356
rect 4344 5296 4408 5300
rect 4424 5356 4488 5360
rect 4424 5300 4428 5356
rect 4428 5300 4484 5356
rect 4484 5300 4488 5356
rect 4424 5296 4488 5300
rect 4504 5356 4568 5360
rect 4504 5300 4508 5356
rect 4508 5300 4564 5356
rect 4564 5300 4568 5356
rect 4504 5296 4568 5300
rect 34984 5356 35048 5360
rect 34984 5300 34988 5356
rect 34988 5300 35044 5356
rect 35044 5300 35048 5356
rect 34984 5296 35048 5300
rect 35064 5356 35128 5360
rect 35064 5300 35068 5356
rect 35068 5300 35124 5356
rect 35124 5300 35128 5356
rect 35064 5296 35128 5300
rect 35144 5356 35208 5360
rect 35144 5300 35148 5356
rect 35148 5300 35204 5356
rect 35204 5300 35208 5356
rect 35144 5296 35208 5300
rect 35224 5356 35288 5360
rect 35224 5300 35228 5356
rect 35228 5300 35284 5356
rect 35284 5300 35288 5356
rect 35224 5296 35288 5300
rect 19624 4690 19688 4694
rect 19624 4634 19628 4690
rect 19628 4634 19684 4690
rect 19684 4634 19688 4690
rect 19624 4630 19688 4634
rect 19704 4690 19768 4694
rect 19704 4634 19708 4690
rect 19708 4634 19764 4690
rect 19764 4634 19768 4690
rect 19704 4630 19768 4634
rect 19784 4690 19848 4694
rect 19784 4634 19788 4690
rect 19788 4634 19844 4690
rect 19844 4634 19848 4690
rect 19784 4630 19848 4634
rect 19864 4690 19928 4694
rect 19864 4634 19868 4690
rect 19868 4634 19924 4690
rect 19924 4634 19928 4690
rect 19864 4630 19928 4634
rect 50344 4690 50408 4694
rect 50344 4634 50348 4690
rect 50348 4634 50404 4690
rect 50404 4634 50408 4690
rect 50344 4630 50408 4634
rect 50424 4690 50488 4694
rect 50424 4634 50428 4690
rect 50428 4634 50484 4690
rect 50484 4634 50488 4690
rect 50424 4630 50488 4634
rect 50504 4690 50568 4694
rect 50504 4634 50508 4690
rect 50508 4634 50564 4690
rect 50564 4634 50568 4690
rect 50504 4630 50568 4634
rect 50584 4690 50648 4694
rect 50584 4634 50588 4690
rect 50588 4634 50644 4690
rect 50644 4634 50648 4690
rect 50584 4630 50648 4634
rect 4264 4024 4328 4028
rect 4264 3968 4268 4024
rect 4268 3968 4324 4024
rect 4324 3968 4328 4024
rect 4264 3964 4328 3968
rect 4344 4024 4408 4028
rect 4344 3968 4348 4024
rect 4348 3968 4404 4024
rect 4404 3968 4408 4024
rect 4344 3964 4408 3968
rect 4424 4024 4488 4028
rect 4424 3968 4428 4024
rect 4428 3968 4484 4024
rect 4484 3968 4488 4024
rect 4424 3964 4488 3968
rect 4504 4024 4568 4028
rect 4504 3968 4508 4024
rect 4508 3968 4564 4024
rect 4564 3968 4568 4024
rect 4504 3964 4568 3968
rect 34984 4024 35048 4028
rect 34984 3968 34988 4024
rect 34988 3968 35044 4024
rect 35044 3968 35048 4024
rect 34984 3964 35048 3968
rect 35064 4024 35128 4028
rect 35064 3968 35068 4024
rect 35068 3968 35124 4024
rect 35124 3968 35128 4024
rect 35064 3964 35128 3968
rect 35144 4024 35208 4028
rect 35144 3968 35148 4024
rect 35148 3968 35204 4024
rect 35204 3968 35208 4024
rect 35144 3964 35208 3968
rect 35224 4024 35288 4028
rect 35224 3968 35228 4024
rect 35228 3968 35284 4024
rect 35284 3968 35288 4024
rect 35224 3964 35288 3968
rect 19624 3358 19688 3362
rect 19624 3302 19628 3358
rect 19628 3302 19684 3358
rect 19684 3302 19688 3358
rect 19624 3298 19688 3302
rect 19704 3358 19768 3362
rect 19704 3302 19708 3358
rect 19708 3302 19764 3358
rect 19764 3302 19768 3358
rect 19704 3298 19768 3302
rect 19784 3358 19848 3362
rect 19784 3302 19788 3358
rect 19788 3302 19844 3358
rect 19844 3302 19848 3358
rect 19784 3298 19848 3302
rect 19864 3358 19928 3362
rect 19864 3302 19868 3358
rect 19868 3302 19924 3358
rect 19924 3302 19928 3358
rect 19864 3298 19928 3302
rect 50344 3358 50408 3362
rect 50344 3302 50348 3358
rect 50348 3302 50404 3358
rect 50404 3302 50408 3358
rect 50344 3298 50408 3302
rect 50424 3358 50488 3362
rect 50424 3302 50428 3358
rect 50428 3302 50484 3358
rect 50484 3302 50488 3358
rect 50424 3298 50488 3302
rect 50504 3358 50568 3362
rect 50504 3302 50508 3358
rect 50508 3302 50564 3358
rect 50564 3302 50568 3358
rect 50504 3298 50568 3302
rect 50584 3358 50648 3362
rect 50584 3302 50588 3358
rect 50588 3302 50644 3358
rect 50644 3302 50648 3358
rect 50584 3298 50648 3302
rect 4264 2692 4328 2696
rect 4264 2636 4268 2692
rect 4268 2636 4324 2692
rect 4324 2636 4328 2692
rect 4264 2632 4328 2636
rect 4344 2692 4408 2696
rect 4344 2636 4348 2692
rect 4348 2636 4404 2692
rect 4404 2636 4408 2692
rect 4344 2632 4408 2636
rect 4424 2692 4488 2696
rect 4424 2636 4428 2692
rect 4428 2636 4484 2692
rect 4484 2636 4488 2692
rect 4424 2632 4488 2636
rect 4504 2692 4568 2696
rect 4504 2636 4508 2692
rect 4508 2636 4564 2692
rect 4564 2636 4568 2692
rect 4504 2632 4568 2636
rect 34984 2692 35048 2696
rect 34984 2636 34988 2692
rect 34988 2636 35044 2692
rect 35044 2636 35048 2692
rect 34984 2632 35048 2636
rect 35064 2692 35128 2696
rect 35064 2636 35068 2692
rect 35068 2636 35124 2692
rect 35124 2636 35128 2692
rect 35064 2632 35128 2636
rect 35144 2692 35208 2696
rect 35144 2636 35148 2692
rect 35148 2636 35204 2692
rect 35204 2636 35208 2692
rect 35144 2632 35208 2636
rect 35224 2692 35288 2696
rect 35224 2636 35228 2692
rect 35228 2636 35284 2692
rect 35284 2636 35288 2692
rect 35224 2632 35288 2636
<< metal4 >>
rect 4256 57308 4576 57324
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 55976 4576 57244
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 54644 4576 55912
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 53312 4576 54580
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 51980 4576 53248
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 50648 4576 51916
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 49316 4576 50584
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 47984 4576 49252
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 46652 4576 47920
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 45320 4576 46588
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 43988 4576 45256
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 42656 4576 43924
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 41324 4576 42592
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 39992 4576 41260
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 38660 4576 39928
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 37328 4576 38596
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 35996 4576 37264
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 34664 4576 35932
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 33332 4576 34600
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 32000 4576 33268
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 30668 4576 31936
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 29336 4576 30604
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 28004 4576 29272
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 26672 4576 27940
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 25340 4576 26608
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 24008 4576 25276
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 22676 4576 23944
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 21344 4576 22612
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 20012 4576 21280
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 18680 4576 19948
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 17348 4576 18616
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 16016 4576 17284
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 14684 4576 15952
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 13352 4576 14620
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 12020 4576 13288
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 10688 4576 11956
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 9356 4576 10624
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 8024 4576 9292
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 6692 4576 7960
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 5360 4576 6628
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 4028 4576 5296
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 2696 4576 3964
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4916 2664 5236 57276
rect 5576 2664 5896 57276
rect 6236 2664 6556 57276
rect 19616 56642 19936 57324
rect 34976 57308 35296 57324
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 55310 19936 56578
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 53978 19936 55246
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 52646 19936 53914
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 51314 19936 52582
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 49982 19936 51250
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 48650 19936 49918
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 47318 19936 48586
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 45986 19936 47254
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 44654 19936 45922
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 43322 19936 44590
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 41990 19936 43258
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 40658 19936 41926
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 39326 19936 40594
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 37994 19936 39262
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 36662 19936 37930
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 35330 19936 36598
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 33998 19936 35266
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 32666 19936 33934
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 31334 19936 32602
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 30002 19936 31270
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 28670 19936 29938
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 27338 19936 28606
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 26006 19936 27274
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 24674 19936 25942
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 23342 19936 24610
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 22010 19936 23278
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 20678 19936 21946
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 19346 19936 20614
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 18014 19936 19282
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 16682 19936 17950
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 15350 19936 16618
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 14018 19936 15286
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 12686 19936 13954
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 11354 19936 12622
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 10022 19936 11290
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 8690 19936 9958
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 7358 19936 8626
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 6026 19936 7294
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 4694 19936 5962
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 3362 19936 4630
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 4256 2616 4576 2632
rect 19616 2616 19936 3298
rect 20276 2664 20596 57276
rect 20936 2664 21256 57276
rect 21596 2664 21916 57276
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 55976 35296 57244
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 54644 35296 55912
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 53312 35296 54580
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 51980 35296 53248
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 50648 35296 51916
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 49316 35296 50584
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 47984 35296 49252
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 46652 35296 47920
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 45320 35296 46588
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 43988 35296 45256
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 42656 35296 43924
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 41324 35296 42592
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 39992 35296 41260
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 38660 35296 39928
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 37328 35296 38596
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 35996 35296 37264
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 34664 35296 35932
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 33332 35296 34600
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 32000 35296 33268
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 30668 35296 31936
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 29336 35296 30604
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 28004 35296 29272
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 26672 35296 27940
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 25340 35296 26608
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 24008 35296 25276
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 22676 35296 23944
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 21344 35296 22612
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 20012 35296 21280
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 18680 35296 19948
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 17348 35296 18616
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 16016 35296 17284
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 14684 35296 15952
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 13352 35296 14620
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 12020 35296 13288
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 10688 35296 11956
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 9356 35296 10624
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 8024 35296 9292
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 6692 35296 7960
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 5360 35296 6628
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 4028 35296 5296
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 2696 35296 3964
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 35636 2664 35956 57276
rect 36296 2664 36616 57276
rect 36956 2664 37276 57276
rect 50336 56642 50656 57324
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 55310 50656 56578
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 53978 50656 55246
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 52646 50656 53914
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 51314 50656 52582
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 49982 50656 51250
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 48650 50656 49918
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 47318 50656 48586
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 45986 50656 47254
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 44654 50656 45922
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 43322 50656 44590
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 41990 50656 43258
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 40658 50656 41926
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 39326 50656 40594
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 37994 50656 39262
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 36662 50656 37930
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 35330 50656 36598
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 33998 50656 35266
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 32666 50656 33934
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 31334 50656 32602
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 30002 50656 31270
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 28670 50656 29938
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 27338 50656 28606
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 26006 50656 27274
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 24674 50656 25942
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 23342 50656 24610
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 22010 50656 23278
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 20678 50656 21946
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 19346 50656 20614
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 18014 50656 19282
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 16682 50656 17950
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 15350 50656 16618
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 14018 50656 15286
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 12686 50656 13954
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 11354 50656 12622
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 10022 50656 11290
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 8690 50656 9958
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 7358 50656 8626
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 6026 50656 7294
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 4694 50656 5962
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 3362 50656 4630
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 34976 2616 35296 2632
rect 50336 2616 50656 3298
rect 50996 2664 51316 57276
rect 51656 2664 51976 57276
rect 52316 2664 52636 57276
use sky130_fd_sc_ls__clkbuf_1  input296 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input295
timestamp 1621261055
transform 1 0 1536 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_0
timestamp 1621261055
transform 1 0 1152 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_8
timestamp 1621261055
transform 1 0 1920 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_8
timestamp 1621261055
transform 1 0 1920 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input319
timestamp 1621261055
transform 1 0 2304 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input297
timestamp 1621261055
transform 1 0 2304 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_16
timestamp 1621261055
transform 1 0 2688 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_16
timestamp 1621261055
transform 1 0 2688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input323
timestamp 1621261055
transform 1 0 3072 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input322
timestamp 1621261055
transform 1 0 3072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_24
timestamp 1621261055
transform 1 0 3456 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3936 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_24
timestamp 1621261055
transform 1 0 3456 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input324
timestamp 1621261055
transform 1 0 3840 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_164 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3840 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_32
timestamp 1621261055
transform 1 0 4224 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 4704 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input325
timestamp 1621261055
transform 1 0 4608 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_40
timestamp 1621261055
transform 1 0 4992 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input298
timestamp 1621261055
transform 1 0 4896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_44
timestamp 1621261055
transform 1 0 5376 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_43
timestamp 1621261055
transform 1 0 5280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input300
timestamp 1621261055
transform 1 0 5568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_50
timestamp 1621261055
transform 1 0 5952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_51
timestamp 1621261055
transform 1 0 6048 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input299
timestamp 1621261055
transform 1 0 5664 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_56
timestamp 1621261055
transform 1 0 6528 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_54 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 6336 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_0_55
timestamp 1621261055
transform 1 0 6432 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_185
timestamp 1621261055
transform 1 0 6432 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_165
timestamp 1621261055
transform 1 0 6528 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_57
timestamp 1621261055
transform 1 0 6624 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input302
timestamp 1621261055
transform 1 0 6912 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input301
timestamp 1621261055
transform 1 0 7008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_64
timestamp 1621261055
transform 1 0 7296 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_65
timestamp 1621261055
transform 1 0 7392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_72
timestamp 1621261055
transform 1 0 8064 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input304
timestamp 1621261055
transform 1 0 7680 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input303
timestamp 1621261055
transform 1 0 7776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_73
timestamp 1621261055
transform 1 0 8160 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input306
timestamp 1621261055
transform 1 0 8448 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 8544 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_80
timestamp 1621261055
transform 1 0 8832 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_80
timestamp 1621261055
transform 1 0 8832 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input309
timestamp 1621261055
transform 1 0 9216 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_166
timestamp 1621261055
transform 1 0 9216 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_88
timestamp 1621261055
transform 1 0 9600 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_85
timestamp 1621261055
transform 1 0 9312 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input311
timestamp 1621261055
transform 1 0 9984 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input307
timestamp 1621261055
transform 1 0 9696 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_96
timestamp 1621261055
transform 1 0 10368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_101
timestamp 1621261055
transform 1 0 10848 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_93
timestamp 1621261055
transform 1 0 10080 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input313
timestamp 1621261055
transform 1 0 10752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input310
timestamp 1621261055
transform 1 0 10464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_104
timestamp 1621261055
transform 1 0 11136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_111
timestamp 1621261055
transform 1 0 11808 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_108
timestamp 1621261055
transform 1 0 11520 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_113
timestamp 1621261055
transform 1 0 12000 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_0_111
timestamp 1621261055
transform 1 0 11808 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_109
timestamp 1621261055
transform 1 0 11616 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_23 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform -1 0 12192 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_186
timestamp 1621261055
transform 1 0 11712 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_167
timestamp 1621261055
transform 1 0 11904 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_118
timestamp 1621261055
transform 1 0 12480 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_121
timestamp 1621261055
transform 1 0 12768 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input167
timestamp 1621261055
transform 1 0 12864 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _013_
timestamp 1621261055
transform -1 0 12480 0 1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_126
timestamp 1621261055
transform 1 0 13248 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input39
timestamp 1621261055
transform 1 0 12960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_127
timestamp 1621261055
transform 1 0 13344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input89
timestamp 1621261055
transform 1 0 13632 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_134
timestamp 1621261055
transform 1 0 14016 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_135
timestamp 1621261055
transform 1 0 14112 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input78
timestamp 1621261055
transform 1 0 13728 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_139
timestamp 1621261055
transform 1 0 14496 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input100
timestamp 1621261055
transform 1 0 14400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_168
timestamp 1621261055
transform 1 0 14592 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_142
timestamp 1621261055
transform 1 0 14784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_141
timestamp 1621261055
transform 1 0 14688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input111
timestamp 1621261055
transform 1 0 15072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input122
timestamp 1621261055
transform 1 0 15168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_150
timestamp 1621261055
transform 1 0 15552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_149
timestamp 1621261055
transform 1 0 15456 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input133
timestamp 1621261055
transform 1 0 15936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_164
timestamp 1621261055
transform 1 0 16896 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_162
timestamp 1621261055
transform 1 0 16704 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_158
timestamp 1621261055
transform 1 0 16320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_164
timestamp 1621261055
transform 1 0 16896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_159
timestamp 1621261055
transform 1 0 16416 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_157
timestamp 1621261055
transform 1 0 16224 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input50
timestamp 1621261055
transform 1 0 16512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_166
timestamp 1621261055
transform 1 0 17088 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_187
timestamp 1621261055
transform 1 0 16992 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_169
timestamp 1621261055
transform 1 0 17280 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_174
timestamp 1621261055
transform 1 0 17856 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_169
timestamp 1621261055
transform 1 0 17376 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input70
timestamp 1621261055
transform 1 0 17472 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input61
timestamp 1621261055
transform 1 0 17760 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_182
timestamp 1621261055
transform 1 0 18624 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_185
timestamp 1621261055
transform 1 0 18912 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_177
timestamp 1621261055
transform 1 0 18144 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input72
timestamp 1621261055
transform 1 0 18240 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input71
timestamp 1621261055
transform 1 0 18528 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input73
timestamp 1621261055
transform 1 0 19008 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_190
timestamp 1621261055
transform 1 0 19392 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_193
timestamp 1621261055
transform 1 0 19680 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_198
timestamp 1621261055
transform 1 0 20160 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_197
timestamp 1621261055
transform 1 0 20064 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_195
timestamp 1621261055
transform 1 0 19872 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input75
timestamp 1621261055
transform 1 0 19776 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_170
timestamp 1621261055
transform 1 0 19968 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input77
timestamp 1621261055
transform 1 0 20544 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input74
timestamp 1621261055
transform 1 0 20448 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_206
timestamp 1621261055
transform 1 0 20928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_205
timestamp 1621261055
transform 1 0 20832 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input80
timestamp 1621261055
transform 1 0 21312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input76
timestamp 1621261055
transform 1 0 21216 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_218
timestamp 1621261055
transform 1 0 22080 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_214
timestamp 1621261055
transform 1 0 21696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_213
timestamp 1621261055
transform 1 0 21600 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_1_221
timestamp 1621261055
transform 1 0 22368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_225
timestamp 1621261055
transform 1 0 22752 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_223
timestamp 1621261055
transform 1 0 22560 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_221
timestamp 1621261055
transform 1 0 22368 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input84
timestamp 1621261055
transform 1 0 22752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_188
timestamp 1621261055
transform 1 0 22272 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_171
timestamp 1621261055
transform 1 0 22656 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_229
timestamp 1621261055
transform 1 0 23136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input82
timestamp 1621261055
transform 1 0 23136 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_237
timestamp 1621261055
transform 1 0 23904 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_233
timestamp 1621261055
transform 1 0 23520 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input86
timestamp 1621261055
transform 1 0 23520 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input85
timestamp 1621261055
transform 1 0 23904 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_245
timestamp 1621261055
transform 1 0 24672 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_241
timestamp 1621261055
transform 1 0 24288 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input88
timestamp 1621261055
transform 1 0 24288 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_251
timestamp 1621261055
transform 1 0 25248 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_249
timestamp 1621261055
transform 1 0 25056 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input91
timestamp 1621261055
transform 1 0 25056 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_172
timestamp 1621261055
transform 1 0 25344 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_253
timestamp 1621261055
transform 1 0 25440 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_253
timestamp 1621261055
transform 1 0 25440 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input92
timestamp 1621261055
transform 1 0 25824 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input90
timestamp 1621261055
transform 1 0 25824 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_269
timestamp 1621261055
transform 1 0 26976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_261
timestamp 1621261055
transform 1 0 26208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_269
timestamp 1621261055
transform 1 0 26976 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_261
timestamp 1621261055
transform 1 0 26208 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input95
timestamp 1621261055
transform 1 0 26592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input93
timestamp 1621261055
transform 1 0 26592 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_273
timestamp 1621261055
transform 1 0 27360 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_276
timestamp 1621261055
transform 1 0 27648 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_277
timestamp 1621261055
transform 1 0 27744 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_189
timestamp 1621261055
transform 1 0 27552 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_281
timestamp 1621261055
transform 1 0 28128 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_279
timestamp 1621261055
transform 1 0 27936 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input99
timestamp 1621261055
transform 1 0 28032 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_173
timestamp 1621261055
transform 1 0 28032 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_284
timestamp 1621261055
transform 1 0 28416 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input98
timestamp 1621261055
transform 1 0 28512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_292
timestamp 1621261055
transform 1 0 29184 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_289
timestamp 1621261055
transform 1 0 28896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input102
timestamp 1621261055
transform 1 0 28800 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input101
timestamp 1621261055
transform 1 0 29280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_300
timestamp 1621261055
transform 1 0 29952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_297
timestamp 1621261055
transform 1 0 29664 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input104
timestamp 1621261055
transform 1 0 29568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_308
timestamp 1621261055
transform 1 0 30720 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_309
timestamp 1621261055
transform 1 0 30816 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_307
timestamp 1621261055
transform 1 0 30624 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_305
timestamp 1621261055
transform 1 0 30432 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input106
timestamp 1621261055
transform 1 0 30336 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_174
timestamp 1621261055
transform 1 0 30720 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input108
timestamp 1621261055
transform 1 0 31104 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input107
timestamp 1621261055
transform 1 0 31200 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_316
timestamp 1621261055
transform 1 0 31488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_317
timestamp 1621261055
transform 1 0 31584 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input112
timestamp 1621261055
transform 1 0 31872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input109
timestamp 1621261055
transform 1 0 31968 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_331
timestamp 1621261055
transform 1 0 32928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_328
timestamp 1621261055
transform 1 0 32640 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_324
timestamp 1621261055
transform 1 0 32256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_325
timestamp 1621261055
transform 1 0 32352 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_190
timestamp 1621261055
transform 1 0 32832 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_0_335
timestamp 1621261055
transform 1 0 33312 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_333
timestamp 1621261055
transform 1 0 33120 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input115
timestamp 1621261055
transform 1 0 33312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_175
timestamp 1621261055
transform 1 0 33408 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_339
timestamp 1621261055
transform 1 0 33696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_337
timestamp 1621261055
transform 1 0 33504 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_345
timestamp 1621261055
transform 1 0 34272 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input118
timestamp 1621261055
transform 1 0 34080 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input114
timestamp 1621261055
transform 1 0 33888 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_347
timestamp 1621261055
transform 1 0 34464 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input117
timestamp 1621261055
transform 1 0 34656 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_355
timestamp 1621261055
transform 1 0 35232 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_353
timestamp 1621261055
transform 1 0 35040 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_66
timestamp 1621261055
transform 1 0 35232 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input120
timestamp 1621261055
transform 1 0 34848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _049_
timestamp 1621261055
transform 1 0 35424 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_360
timestamp 1621261055
transform 1 0 35712 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input123
timestamp 1621261055
transform 1 0 35616 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_363
timestamp 1621261055
transform 1 0 36000 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_365
timestamp 1621261055
transform 1 0 36192 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_176
timestamp 1621261055
transform 1 0 36096 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_371
timestamp 1621261055
transform 1 0 36768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input125
timestamp 1621261055
transform 1 0 36384 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input124
timestamp 1621261055
transform 1 0 36576 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_373
timestamp 1621261055
transform 1 0 36960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input127
timestamp 1621261055
transform 1 0 37152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input126
timestamp 1621261055
transform 1 0 37344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_386
timestamp 1621261055
transform 1 0 38208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_383
timestamp 1621261055
transform 1 0 37920 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_379
timestamp 1621261055
transform 1 0 37536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_381
timestamp 1621261055
transform 1 0 37728 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_191
timestamp 1621261055
transform 1 0 38112 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_394
timestamp 1621261055
transform 1 0 38976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_393
timestamp 1621261055
transform 1 0 38880 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_391
timestamp 1621261055
transform 1 0 38688 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_389
timestamp 1621261055
transform 1 0 38496 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input131
timestamp 1621261055
transform 1 0 38592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_177
timestamp 1621261055
transform 1 0 38784 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input134
timestamp 1621261055
transform 1 0 39360 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input130
timestamp 1621261055
transform 1 0 39264 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_402
timestamp 1621261055
transform 1 0 39744 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_401
timestamp 1621261055
transform 1 0 39648 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input136
timestamp 1621261055
transform 1 0 40128 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input132
timestamp 1621261055
transform 1 0 40032 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_410
timestamp 1621261055
transform 1 0 40512 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_409
timestamp 1621261055
transform 1 0 40416 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _105_
timestamp 1621261055
transform 1 0 40800 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_418
timestamp 1621261055
transform 1 0 41280 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_416
timestamp 1621261055
transform 1 0 41088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input138
timestamp 1621261055
transform 1 0 40896 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_178
timestamp 1621261055
transform 1 0 41472 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_421
timestamp 1621261055
transform 1 0 41568 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input140
timestamp 1621261055
transform 1 0 41664 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input139
timestamp 1621261055
transform 1 0 41952 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_426
timestamp 1621261055
transform 1 0 42048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_429
timestamp 1621261055
transform 1 0 42336 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_434
timestamp 1621261055
transform 1 0 42816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input142
timestamp 1621261055
transform 1 0 42432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input141
timestamp 1621261055
transform 1 0 42720 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_438
timestamp 1621261055
transform 1 0 43200 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_437
timestamp 1621261055
transform 1 0 43104 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_441
timestamp 1621261055
transform 1 0 43488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_192
timestamp 1621261055
transform 1 0 43392 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _217_
timestamp 1621261055
transform 1 0 43488 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_444
timestamp 1621261055
transform 1 0 43776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input146
timestamp 1621261055
transform 1 0 43872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_449
timestamp 1621261055
transform 1 0 44256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_449
timestamp 1621261055
transform 1 0 44256 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_179
timestamp 1621261055
transform 1 0 44160 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input149
timestamp 1621261055
transform 1 0 44640 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input147
timestamp 1621261055
transform 1 0 44640 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_457
timestamp 1621261055
transform 1 0 45024 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_457
timestamp 1621261055
transform 1 0 45024 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input151
timestamp 1621261055
transform 1 0 45408 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input150
timestamp 1621261055
transform 1 0 45408 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_465
timestamp 1621261055
transform 1 0 45792 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_465
timestamp 1621261055
transform 1 0 45792 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input153
timestamp 1621261055
transform 1 0 46176 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _188_
timestamp 1621261055
transform 1 0 46176 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_473
timestamp 1621261055
transform 1 0 46560 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_472
timestamp 1621261055
transform 1 0 46464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_180
timestamp 1621261055
transform 1 0 46848 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_481
timestamp 1621261055
transform 1 0 47328 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_477
timestamp 1621261055
transform 1 0 46944 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input156
timestamp 1621261055
transform 1 0 46944 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input154
timestamp 1621261055
transform 1 0 47328 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_489
timestamp 1621261055
transform 1 0 48096 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_485
timestamp 1621261055
transform 1 0 47712 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input159
timestamp 1621261055
transform 1 0 47712 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input157
timestamp 1621261055
transform 1 0 48096 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_496
timestamp 1621261055
transform 1 0 48768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_493
timestamp 1621261055
transform 1 0 48480 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_500
timestamp 1621261055
transform 1 0 49152 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_493
timestamp 1621261055
transform 1 0 48480 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input162
timestamp 1621261055
transform 1 0 49152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_193
timestamp 1621261055
transform 1 0 48672 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _180_
timestamp 1621261055
transform 1 0 48864 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_1_504
timestamp 1621261055
transform 1 0 49536 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_181
timestamp 1621261055
transform 1 0 49536 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_505
timestamp 1621261055
transform 1 0 49632 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input40
timestamp 1621261055
transform 1 0 50016 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_512
timestamp 1621261055
transform 1 0 50304 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_513
timestamp 1621261055
transform 1 0 50400 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input42
timestamp 1621261055
transform 1 0 50400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_517
timestamp 1621261055
transform 1 0 50784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input41
timestamp 1621261055
transform 1 0 50784 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_521
timestamp 1621261055
transform 1 0 51168 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input43
timestamp 1621261055
transform 1 0 51168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_525
timestamp 1621261055
transform 1 0 51552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _168_
timestamp 1621261055
transform 1 0 51552 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_533
timestamp 1621261055
transform 1 0 52320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_533
timestamp 1621261055
transform 1 0 52320 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_528
timestamp 1621261055
transform 1 0 51840 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input44
timestamp 1621261055
transform 1 0 51936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_182
timestamp 1621261055
transform 1 0 52224 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_541
timestamp 1621261055
transform 1 0 53088 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_541
timestamp 1621261055
transform 1 0 53088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input46
timestamp 1621261055
transform 1 0 52704 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input45
timestamp 1621261055
transform 1 0 52704 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input47
timestamp 1621261055
transform 1 0 53472 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_551
timestamp 1621261055
transform 1 0 54048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_549
timestamp 1621261055
transform 1 0 53856 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_0_549
timestamp 1621261055
transform 1 0 53856 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input51
timestamp 1621261055
transform 1 0 54432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_194
timestamp 1621261055
transform 1 0 53952 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_559
timestamp 1621261055
transform 1 0 54816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_561
timestamp 1621261055
transform 1 0 55008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_559
timestamp 1621261055
transform 1 0 54816 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_557
timestamp 1621261055
transform 1 0 54624 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input54
timestamp 1621261055
transform 1 0 55200 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_183
timestamp 1621261055
transform 1 0 54912 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_567
timestamp 1621261055
transform 1 0 55584 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input52
timestamp 1621261055
transform 1 0 55392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_575
timestamp 1621261055
transform 1 0 56352 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_569
timestamp 1621261055
transform 1 0 55776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input56
timestamp 1621261055
transform 1 0 55968 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input55
timestamp 1621261055
transform 1 0 56160 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_583
timestamp 1621261055
transform 1 0 57120 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_577
timestamp 1621261055
transform 1 0 56544 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input58
timestamp 1621261055
transform 1 0 56736 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_587
timestamp 1621261055
transform 1 0 57504 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_585
timestamp 1621261055
transform 1 0 57312 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input59
timestamp 1621261055
transform 1 0 57504 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_184
timestamp 1621261055
transform 1 0 57600 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_1
timestamp 1621261055
transform -1 0 58848 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_3
timestamp 1621261055
transform -1 0 58848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_589
timestamp 1621261055
transform 1 0 57696 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_1_591
timestamp 1621261055
transform 1 0 57888 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_595
timestamp 1621261055
transform 1 0 58272 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_4
timestamp 1621261055
transform 1 0 1152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input308
timestamp 1621261055
transform 1 0 1536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input330
timestamp 1621261055
transform 1 0 2304 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input341
timestamp 1621261055
transform 1 0 3072 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_8
timestamp 1621261055
transform 1 0 1920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_16
timestamp 1621261055
transform 1 0 2688 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_195
timestamp 1621261055
transform 1 0 3840 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input326
timestamp 1621261055
transform 1 0 4320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input328
timestamp 1621261055
transform 1 0 5088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_24
timestamp 1621261055
transform 1 0 3456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_29
timestamp 1621261055
transform 1 0 3936 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_37
timestamp 1621261055
transform 1 0 4704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input331
timestamp 1621261055
transform 1 0 5856 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input333
timestamp 1621261055
transform 1 0 6624 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_45
timestamp 1621261055
transform 1 0 5472 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_53
timestamp 1621261055
transform 1 0 6240 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_61
timestamp 1621261055
transform 1 0 7008 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_196
timestamp 1621261055
transform 1 0 9120 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input305
timestamp 1621261055
transform 1 0 7392 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input335
timestamp 1621261055
transform 1 0 8160 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_69
timestamp 1621261055
transform 1 0 7776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_77
timestamp 1621261055
transform 1 0 8544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_81
timestamp 1621261055
transform 1 0 8928 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_84
timestamp 1621261055
transform 1 0 9216 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input312
timestamp 1621261055
transform 1 0 9600 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input314
timestamp 1621261055
transform 1 0 10368 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input315
timestamp 1621261055
transform 1 0 11136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_92
timestamp 1621261055
transform 1 0 9984 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_100
timestamp 1621261055
transform 1 0 10752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input316
timestamp 1621261055
transform 1 0 11904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input317
timestamp 1621261055
transform 1 0 12672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_108
timestamp 1621261055
transform 1 0 11520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_116
timestamp 1621261055
transform 1 0 12288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_124
timestamp 1621261055
transform 1 0 13056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_197
timestamp 1621261055
transform 1 0 14400 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input206
timestamp 1621261055
transform 1 0 13536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_128
timestamp 1621261055
transform 1 0 13440 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_133
timestamp 1621261055
transform 1 0 13920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_137
timestamp 1621261055
transform 1 0 14304 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_139
timestamp 1621261055
transform 1 0 14496 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_147
timestamp 1621261055
transform 1 0 15264 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input144
timestamp 1621261055
transform 1 0 15456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input155
timestamp 1621261055
transform 1 0 16224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input166
timestamp 1621261055
transform 1 0 16992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_153
timestamp 1621261055
transform 1 0 15840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_161
timestamp 1621261055
transform 1 0 16608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input178
timestamp 1621261055
transform 1 0 17760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input198
timestamp 1621261055
transform 1 0 18528 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_169
timestamp 1621261055
transform 1 0 17376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_177
timestamp 1621261055
transform 1 0 18144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_185
timestamp 1621261055
transform 1 0 18912 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_198
timestamp 1621261055
transform 1 0 19680 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input79
timestamp 1621261055
transform 1 0 20256 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input81
timestamp 1621261055
transform 1 0 21024 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_194
timestamp 1621261055
transform 1 0 19776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_198
timestamp 1621261055
transform 1 0 20160 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_203
timestamp 1621261055
transform 1 0 20640 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input83
timestamp 1621261055
transform 1 0 21792 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input87
timestamp 1621261055
transform 1 0 23232 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_211
timestamp 1621261055
transform 1 0 21408 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_219
timestamp 1621261055
transform 1 0 22176 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_227
timestamp 1621261055
transform 1 0 22944 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_229
timestamp 1621261055
transform 1 0 23136 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_199
timestamp 1621261055
transform 1 0 24960 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input211
timestamp 1621261055
transform 1 0 24000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_234
timestamp 1621261055
transform 1 0 23616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_242
timestamp 1621261055
transform 1 0 24384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_246
timestamp 1621261055
transform 1 0 24768 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_249
timestamp 1621261055
transform 1 0 25056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input94
timestamp 1621261055
transform 1 0 25440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input96
timestamp 1621261055
transform 1 0 26208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input97
timestamp 1621261055
transform 1 0 26976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_257
timestamp 1621261055
transform 1 0 25824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_265
timestamp 1621261055
transform 1 0 26592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_273
timestamp 1621261055
transform 1 0 27360 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input103
timestamp 1621261055
transform 1 0 28320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input105
timestamp 1621261055
transform 1 0 29088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_281
timestamp 1621261055
transform 1 0 28128 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_287
timestamp 1621261055
transform 1 0 28704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_200
timestamp 1621261055
transform 1 0 30240 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input110
timestamp 1621261055
transform 1 0 30912 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_295
timestamp 1621261055
transform 1 0 29472 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_304
timestamp 1621261055
transform 1 0 30336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_308
timestamp 1621261055
transform 1 0 30720 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_314
timestamp 1621261055
transform 1 0 31296 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input113
timestamp 1621261055
transform 1 0 31680 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input116
timestamp 1621261055
transform 1 0 32736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_322
timestamp 1621261055
transform 1 0 32064 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_326
timestamp 1621261055
transform 1 0 32448 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_328
timestamp 1621261055
transform 1 0 32640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_333
timestamp 1621261055
transform 1 0 33120 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input119
timestamp 1621261055
transform 1 0 33888 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input121
timestamp 1621261055
transform 1 0 34656 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_345
timestamp 1621261055
transform 1 0 34272 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_353
timestamp 1621261055
transform 1 0 35040 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_357
timestamp 1621261055
transform 1 0 35424 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_201
timestamp 1621261055
transform 1 0 35520 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input128
timestamp 1621261055
transform 1 0 36768 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input247
timestamp 1621261055
transform 1 0 36000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_359
timestamp 1621261055
transform 1 0 35616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_367
timestamp 1621261055
transform 1 0 36384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_375
timestamp 1621261055
transform 1 0 37152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input129
timestamp 1621261055
transform 1 0 37536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input135
timestamp 1621261055
transform 1 0 38976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_383
timestamp 1621261055
transform 1 0 37920 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_391
timestamp 1621261055
transform 1 0 38688 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_393
timestamp 1621261055
transform 1 0 38880 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_398
timestamp 1621261055
transform 1 0 39360 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _024_
timestamp 1621261055
transform 1 0 41280 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_202
timestamp 1621261055
transform 1 0 40800 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input137
timestamp 1621261055
transform 1 0 39744 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_0
timestamp 1621261055
transform 1 0 41088 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_406
timestamp 1621261055
transform 1 0 40128 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_410
timestamp 1621261055
transform 1 0 40512 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_412
timestamp 1621261055
transform 1 0 40704 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_414
timestamp 1621261055
transform 1 0 40896 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input143
timestamp 1621261055
transform 1 0 41952 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input145
timestamp 1621261055
transform 1 0 42720 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input148
timestamp 1621261055
transform 1 0 43488 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_421
timestamp 1621261055
transform 1 0 41568 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_429
timestamp 1621261055
transform 1 0 42336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_437
timestamp 1621261055
transform 1 0 43104 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _131_
timestamp 1621261055
transform 1 0 44256 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input152
timestamp 1621261055
transform 1 0 44928 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_445
timestamp 1621261055
transform 1 0 43872 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_452
timestamp 1621261055
transform 1 0 44544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_460
timestamp 1621261055
transform 1 0 45312 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_203
timestamp 1621261055
transform 1 0 46080 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input158
timestamp 1621261055
transform 1 0 46752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input160
timestamp 1621261055
transform 1 0 47520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_469
timestamp 1621261055
transform 1 0 46176 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_473
timestamp 1621261055
transform 1 0 46560 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_479
timestamp 1621261055
transform 1 0 47136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input161
timestamp 1621261055
transform 1 0 48288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input163
timestamp 1621261055
transform 1 0 49056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_487
timestamp 1621261055
transform 1 0 47904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_495
timestamp 1621261055
transform 1 0 48672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_503
timestamp 1621261055
transform 1 0 49440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_204
timestamp 1621261055
transform 1 0 51360 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input164
timestamp 1621261055
transform 1 0 49824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input168
timestamp 1621261055
transform 1 0 50592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_511
timestamp 1621261055
transform 1 0 50208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_519
timestamp 1621261055
transform 1 0 50976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_524
timestamp 1621261055
transform 1 0 51456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input48
timestamp 1621261055
transform 1 0 52608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input49
timestamp 1621261055
transform 1 0 53376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input171
timestamp 1621261055
transform 1 0 51840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_532
timestamp 1621261055
transform 1 0 52224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_540
timestamp 1621261055
transform 1 0 52992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _161_
timestamp 1621261055
transform 1 0 54912 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input53
timestamp 1621261055
transform 1 0 54144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input57
timestamp 1621261055
transform 1 0 55584 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_548
timestamp 1621261055
transform 1 0 53760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_556
timestamp 1621261055
transform 1 0 54528 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_563
timestamp 1621261055
transform 1 0 55200 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_205
timestamp 1621261055
transform 1 0 56640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input60
timestamp 1621261055
transform 1 0 57120 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_571
timestamp 1621261055
transform 1 0 55968 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_575
timestamp 1621261055
transform 1 0 56352 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_577
timestamp 1621261055
transform 1 0 56544 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_579
timestamp 1621261055
transform 1 0 56736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_587
timestamp 1621261055
transform 1 0 57504 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_5
timestamp 1621261055
transform -1 0 58848 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_595
timestamp 1621261055
transform 1 0 58272 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_6
timestamp 1621261055
transform 1 0 1152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input329
timestamp 1621261055
transform 1 0 1536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input352
timestamp 1621261055
transform 1 0 2304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input355
timestamp 1621261055
transform 1 0 3072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_8
timestamp 1621261055
transform 1 0 1920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_16
timestamp 1621261055
transform 1 0 2688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input327
timestamp 1621261055
transform 1 0 4128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_24
timestamp 1621261055
transform 1 0 3456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_28
timestamp 1621261055
transform 1 0 3840 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_30
timestamp 1621261055
transform 1 0 4032 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_3_35
timestamp 1621261055
transform 1 0 4512 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_206
timestamp 1621261055
transform 1 0 6432 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input332
timestamp 1621261055
transform 1 0 5376 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input334
timestamp 1621261055
transform 1 0 6912 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_43
timestamp 1621261055
transform 1 0 5280 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_3_48
timestamp 1621261055
transform 1 0 5760 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_52
timestamp 1621261055
transform 1 0 6144 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_54
timestamp 1621261055
transform 1 0 6336 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_3_56
timestamp 1621261055
transform 1 0 6528 0 1 4662
box -38 -49 422 715
use AND2X1  AND2X1
timestamp 1624196784
transform 1 0 7680 0 1 4662
box 0 -48 1152 714
use sky130_fd_sc_ls__clkbuf_1  input339
timestamp 1621261055
transform 1 0 9216 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_78
timestamp 1621261055
transform 1 0 7488 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_64
timestamp 1621261055
transform 1 0 7296 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_80
timestamp 1621261055
transform 1 0 8832 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input340
timestamp 1621261055
transform 1 0 9984 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input343
timestamp 1621261055
transform 1 0 10752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_88
timestamp 1621261055
transform 1 0 9600 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_96
timestamp 1621261055
transform 1 0 10368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_104
timestamp 1621261055
transform 1 0 11136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_207
timestamp 1621261055
transform 1 0 11712 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input318
timestamp 1621261055
transform 1 0 12192 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input320
timestamp 1621261055
transform 1 0 12960 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_108
timestamp 1621261055
transform 1 0 11520 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_111
timestamp 1621261055
transform 1 0 11808 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_119
timestamp 1621261055
transform 1 0 12576 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input217
timestamp 1621261055
transform 1 0 13920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input228
timestamp 1621261055
transform 1 0 14688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_127
timestamp 1621261055
transform 1 0 13344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_131
timestamp 1621261055
transform 1 0 13728 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_137
timestamp 1621261055
transform 1 0 14304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_145
timestamp 1621261055
transform 1 0 15072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_208
timestamp 1621261055
transform 1 0 16992 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input239
timestamp 1621261055
transform 1 0 15456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input261
timestamp 1621261055
transform 1 0 16224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_153
timestamp 1621261055
transform 1 0 15840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_161
timestamp 1621261055
transform 1 0 16608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_166
timestamp 1621261055
transform 1 0 17088 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input189
timestamp 1621261055
transform 1 0 17472 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input199
timestamp 1621261055
transform 1 0 18240 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input200
timestamp 1621261055
transform 1 0 19008 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_174
timestamp 1621261055
transform 1 0 17856 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_182
timestamp 1621261055
transform 1 0 18624 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input202
timestamp 1621261055
transform 1 0 19776 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input203
timestamp 1621261055
transform 1 0 20544 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input205
timestamp 1621261055
transform 1 0 21312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_190
timestamp 1621261055
transform 1 0 19392 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_198
timestamp 1621261055
transform 1 0 20160 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_206
timestamp 1621261055
transform 1 0 20928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_209
timestamp 1621261055
transform 1 0 22272 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input209
timestamp 1621261055
transform 1 0 22752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_214
timestamp 1621261055
transform 1 0 21696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_218
timestamp 1621261055
transform 1 0 22080 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_221
timestamp 1621261055
transform 1 0 22368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_229
timestamp 1621261055
transform 1 0 23136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input212
timestamp 1621261055
transform 1 0 23520 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input214
timestamp 1621261055
transform 1 0 24288 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input216
timestamp 1621261055
transform 1 0 25056 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_237
timestamp 1621261055
transform 1 0 23904 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_245
timestamp 1621261055
transform 1 0 24672 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input218
timestamp 1621261055
transform 1 0 25824 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input220
timestamp 1621261055
transform 1 0 26592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_253
timestamp 1621261055
transform 1 0 25440 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_261
timestamp 1621261055
transform 1 0 26208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_269
timestamp 1621261055
transform 1 0 26976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_273
timestamp 1621261055
transform 1 0 27360 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_210
timestamp 1621261055
transform 1 0 27552 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input224
timestamp 1621261055
transform 1 0 28032 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input227
timestamp 1621261055
transform 1 0 28800 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_276
timestamp 1621261055
transform 1 0 27648 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_284
timestamp 1621261055
transform 1 0 28416 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_292
timestamp 1621261055
transform 1 0 29184 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input230
timestamp 1621261055
transform 1 0 29568 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input232
timestamp 1621261055
transform 1 0 30336 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input233
timestamp 1621261055
transform 1 0 31104 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_300
timestamp 1621261055
transform 1 0 29952 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_308
timestamp 1621261055
transform 1 0 30720 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_211
timestamp 1621261055
transform 1 0 32832 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input236
timestamp 1621261055
transform 1 0 31872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input241
timestamp 1621261055
transform 1 0 33312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_316
timestamp 1621261055
transform 1 0 31488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_324
timestamp 1621261055
transform 1 0 32256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_328
timestamp 1621261055
transform 1 0 32640 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_331
timestamp 1621261055
transform 1 0 32928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input243
timestamp 1621261055
transform 1 0 34080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input245
timestamp 1621261055
transform 1 0 34848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_339
timestamp 1621261055
transform 1 0 33696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_347
timestamp 1621261055
transform 1 0 34464 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_355
timestamp 1621261055
transform 1 0 35232 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input248
timestamp 1621261055
transform 1 0 35616 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input249
timestamp 1621261055
transform 1 0 36384 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input252
timestamp 1621261055
transform 1 0 37152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_363
timestamp 1621261055
transform 1 0 36000 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_371
timestamp 1621261055
transform 1 0 36768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_212
timestamp 1621261055
transform 1 0 38112 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input256
timestamp 1621261055
transform 1 0 38592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input258
timestamp 1621261055
transform 1 0 39360 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_379
timestamp 1621261055
transform 1 0 37536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_383
timestamp 1621261055
transform 1 0 37920 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_386
timestamp 1621261055
transform 1 0 38208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_394
timestamp 1621261055
transform 1 0 38976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input260
timestamp 1621261055
transform 1 0 40128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input264
timestamp 1621261055
transform 1 0 40896 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_402
timestamp 1621261055
transform 1 0 39744 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_410
timestamp 1621261055
transform 1 0 40512 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_418
timestamp 1621261055
transform 1 0 41280 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_213
timestamp 1621261055
transform 1 0 43392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input265
timestamp 1621261055
transform 1 0 41664 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input268
timestamp 1621261055
transform 1 0 42432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_426
timestamp 1621261055
transform 1 0 42048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_434
timestamp 1621261055
transform 1 0 42816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_438
timestamp 1621261055
transform 1 0 43200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_441
timestamp 1621261055
transform 1 0 43488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input273
timestamp 1621261055
transform 1 0 43872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input275
timestamp 1621261055
transform 1 0 44640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input277
timestamp 1621261055
transform 1 0 45408 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_449
timestamp 1621261055
transform 1 0 44256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_457
timestamp 1621261055
transform 1 0 45024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input279
timestamp 1621261055
transform 1 0 46176 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input280
timestamp 1621261055
transform 1 0 46944 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_465
timestamp 1621261055
transform 1 0 45792 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_473
timestamp 1621261055
transform 1 0 46560 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_481
timestamp 1621261055
transform 1 0 47328 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_214
timestamp 1621261055
transform 1 0 48672 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input165
timestamp 1621261055
transform 1 0 49344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input284
timestamp 1621261055
transform 1 0 47712 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_489
timestamp 1621261055
transform 1 0 48096 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_493
timestamp 1621261055
transform 1 0 48480 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_496
timestamp 1621261055
transform 1 0 48768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_500
timestamp 1621261055
transform 1 0 49152 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input169
timestamp 1621261055
transform 1 0 50304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input170
timestamp 1621261055
transform 1 0 51072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_506
timestamp 1621261055
transform 1 0 49728 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_510
timestamp 1621261055
transform 1 0 50112 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_516
timestamp 1621261055
transform 1 0 50688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_524
timestamp 1621261055
transform 1 0 51456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input172
timestamp 1621261055
transform 1 0 51840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input173
timestamp 1621261055
transform 1 0 52608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_532
timestamp 1621261055
transform 1 0 52224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_540
timestamp 1621261055
transform 1 0 52992 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_215
timestamp 1621261055
transform 1 0 53952 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input68
timestamp 1621261055
transform 1 0 55488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input177
timestamp 1621261055
transform 1 0 54432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_548
timestamp 1621261055
transform 1 0 53760 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_551
timestamp 1621261055
transform 1 0 54048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_559
timestamp 1621261055
transform 1 0 54816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_563
timestamp 1621261055
transform 1 0 55200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_565
timestamp 1621261055
transform 1 0 55392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input62
timestamp 1621261055
transform 1 0 57024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input64
timestamp 1621261055
transform 1 0 56256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_570
timestamp 1621261055
transform 1 0 55872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_578
timestamp 1621261055
transform 1 0 56640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_586
timestamp 1621261055
transform 1 0 57408 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _184_
timestamp 1621261055
transform 1 0 57792 0 1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_7
timestamp 1621261055
transform -1 0 58848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_593
timestamp 1621261055
transform 1 0 58080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_8
timestamp 1621261055
transform 1 0 1152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input356
timestamp 1621261055
transform 1 0 2784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input362
timestamp 1621261055
transform 1 0 1536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_8
timestamp 1621261055
transform 1 0 1920 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_4_16
timestamp 1621261055
transform 1 0 2688 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_21
timestamp 1621261055
transform 1 0 3168 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_216
timestamp 1621261055
transform 1 0 3840 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input358
timestamp 1621261055
transform 1 0 4320 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input360
timestamp 1621261055
transform 1 0 5088 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_25
timestamp 1621261055
transform 1 0 3552 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_27
timestamp 1621261055
transform 1 0 3744 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_29
timestamp 1621261055
transform 1 0 3936 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_37
timestamp 1621261055
transform 1 0 4704 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input336
timestamp 1621261055
transform 1 0 6816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output574 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform -1 0 6240 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_214
timestamp 1621261055
transform -1 0 5856 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_45
timestamp 1621261055
transform 1 0 5472 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_53
timestamp 1621261055
transform 1 0 6240 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_57
timestamp 1621261055
transform 1 0 6624 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_63
timestamp 1621261055
transform 1 0 7200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_217
timestamp 1621261055
transform 1 0 9120 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input337
timestamp 1621261055
transform 1 0 7584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input338
timestamp 1621261055
transform 1 0 8352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_71
timestamp 1621261055
transform 1 0 7968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_79
timestamp 1621261055
transform 1 0 8736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_84
timestamp 1621261055
transform 1 0 9216 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input342
timestamp 1621261055
transform 1 0 9600 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input345
timestamp 1621261055
transform 1 0 10368 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input347
timestamp 1621261055
transform 1 0 11136 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_92
timestamp 1621261055
transform 1 0 9984 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_100
timestamp 1621261055
transform 1 0 10752 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input321
timestamp 1621261055
transform 1 0 12576 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_108
timestamp 1621261055
transform 1 0 11520 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_116
timestamp 1621261055
transform 1 0 12288 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_118
timestamp 1621261055
transform 1 0 12480 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_123
timestamp 1621261055
transform 1 0 12960 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_218
timestamp 1621261055
transform 1 0 14400 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input250
timestamp 1621261055
transform 1 0 14976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input351
timestamp 1621261055
transform 1 0 13344 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_131
timestamp 1621261055
transform 1 0 13728 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_135
timestamp 1621261055
transform 1 0 14112 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_137
timestamp 1621261055
transform 1 0 14304 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_139
timestamp 1621261055
transform 1 0 14496 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_143
timestamp 1621261055
transform 1 0 14880 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input272
timestamp 1621261055
transform 1 0 15744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input283
timestamp 1621261055
transform 1 0 16512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input294
timestamp 1621261055
transform 1 0 17280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_148
timestamp 1621261055
transform 1 0 15360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_156
timestamp 1621261055
transform 1 0 16128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_164
timestamp 1621261055
transform 1 0 16896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input201
timestamp 1621261055
transform 1 0 18720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_172
timestamp 1621261055
transform 1 0 17664 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_180
timestamp 1621261055
transform 1 0 18432 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_182
timestamp 1621261055
transform 1 0 18624 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_187
timestamp 1621261055
transform 1 0 19104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_219
timestamp 1621261055
transform 1 0 19680 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input204
timestamp 1621261055
transform 1 0 20160 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input207
timestamp 1621261055
transform 1 0 20928 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_191
timestamp 1621261055
transform 1 0 19488 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_194
timestamp 1621261055
transform 1 0 19776 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_202
timestamp 1621261055
transform 1 0 20544 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_210
timestamp 1621261055
transform 1 0 21312 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input208
timestamp 1621261055
transform 1 0 21696 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input210
timestamp 1621261055
transform 1 0 22464 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input213
timestamp 1621261055
transform 1 0 23232 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_218
timestamp 1621261055
transform 1 0 22080 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_226
timestamp 1621261055
transform 1 0 22848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_220
timestamp 1621261055
transform 1 0 24960 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input215
timestamp 1621261055
transform 1 0 24000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_234
timestamp 1621261055
transform 1 0 23616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_242
timestamp 1621261055
transform 1 0 24384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_246
timestamp 1621261055
transform 1 0 24768 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_249
timestamp 1621261055
transform 1 0 25056 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input219
timestamp 1621261055
transform 1 0 25440 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input221
timestamp 1621261055
transform 1 0 26208 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input223
timestamp 1621261055
transform 1 0 26976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_257
timestamp 1621261055
transform 1 0 25824 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_265
timestamp 1621261055
transform 1 0 26592 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_273
timestamp 1621261055
transform 1 0 27360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input226
timestamp 1621261055
transform 1 0 27744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input229
timestamp 1621261055
transform 1 0 28512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input231
timestamp 1621261055
transform 1 0 29280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_281
timestamp 1621261055
transform 1 0 28128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_289
timestamp 1621261055
transform 1 0 28896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_221
timestamp 1621261055
transform 1 0 30240 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input235
timestamp 1621261055
transform 1 0 30720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_297
timestamp 1621261055
transform 1 0 29664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_301
timestamp 1621261055
transform 1 0 30048 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_304
timestamp 1621261055
transform 1 0 30336 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_312
timestamp 1621261055
transform 1 0 31104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input237
timestamp 1621261055
transform 1 0 31488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input240
timestamp 1621261055
transform 1 0 32256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input242
timestamp 1621261055
transform 1 0 33024 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_320
timestamp 1621261055
transform 1 0 31872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_328
timestamp 1621261055
transform 1 0 32640 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_336
timestamp 1621261055
transform 1 0 33408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input244
timestamp 1621261055
transform 1 0 33792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input246
timestamp 1621261055
transform 1 0 34560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_344
timestamp 1621261055
transform 1 0 34176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_352
timestamp 1621261055
transform 1 0 34944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_356
timestamp 1621261055
transform 1 0 35328 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_222
timestamp 1621261055
transform 1 0 35520 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input251
timestamp 1621261055
transform 1 0 36000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input253
timestamp 1621261055
transform 1 0 36768 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_359
timestamp 1621261055
transform 1 0 35616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_367
timestamp 1621261055
transform 1 0 36384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_375
timestamp 1621261055
transform 1 0 37152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input255
timestamp 1621261055
transform 1 0 37536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input257
timestamp 1621261055
transform 1 0 38304 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input259
timestamp 1621261055
transform 1 0 39072 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_383
timestamp 1621261055
transform 1 0 37920 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_391
timestamp 1621261055
transform 1 0 38688 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_399
timestamp 1621261055
transform 1 0 39456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_223
timestamp 1621261055
transform 1 0 40800 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input263
timestamp 1621261055
transform 1 0 39840 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input267
timestamp 1621261055
transform 1 0 41280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_407
timestamp 1621261055
transform 1 0 40224 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_411
timestamp 1621261055
transform 1 0 40608 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_414
timestamp 1621261055
transform 1 0 40896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input269
timestamp 1621261055
transform 1 0 42048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input271
timestamp 1621261055
transform 1 0 42816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_422
timestamp 1621261055
transform 1 0 41664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_430
timestamp 1621261055
transform 1 0 42432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_438
timestamp 1621261055
transform 1 0 43200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input274
timestamp 1621261055
transform 1 0 43584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input276
timestamp 1621261055
transform 1 0 44352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input278
timestamp 1621261055
transform 1 0 45120 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_446
timestamp 1621261055
transform 1 0 43968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_454
timestamp 1621261055
transform 1 0 44736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_462
timestamp 1621261055
transform 1 0 45504 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_224
timestamp 1621261055
transform 1 0 46080 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input282
timestamp 1621261055
transform 1 0 46560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input285
timestamp 1621261055
transform 1 0 47328 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_466
timestamp 1621261055
transform 1 0 45888 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_469
timestamp 1621261055
transform 1 0 46176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_477
timestamp 1621261055
transform 1 0 46944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input287
timestamp 1621261055
transform 1 0 48096 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input289
timestamp 1621261055
transform 1 0 48864 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_485
timestamp 1621261055
transform 1 0 47712 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_493
timestamp 1621261055
transform 1 0 48480 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_501
timestamp 1621261055
transform 1 0 49248 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_225
timestamp 1621261055
transform 1 0 51360 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input290
timestamp 1621261055
transform 1 0 49632 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input292
timestamp 1621261055
transform 1 0 50400 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_509
timestamp 1621261055
transform 1 0 50016 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_517
timestamp 1621261055
transform 1 0 50784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_521
timestamp 1621261055
transform 1 0 51168 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_524
timestamp 1621261055
transform 1 0 51456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input174
timestamp 1621261055
transform 1 0 52128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input175
timestamp 1621261055
transform 1 0 52896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_528
timestamp 1621261055
transform 1 0 51840 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_530
timestamp 1621261055
transform 1 0 52032 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_535
timestamp 1621261055
transform 1 0 52512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_543
timestamp 1621261055
transform 1 0 53280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _101_
timestamp 1621261055
transform 1 0 55200 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input176
timestamp 1621261055
transform 1 0 53664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input179
timestamp 1621261055
transform 1 0 54432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_551
timestamp 1621261055
transform 1 0 54048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_559
timestamp 1621261055
transform 1 0 54816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_566
timestamp 1621261055
transform 1 0 55488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_226
timestamp 1621261055
transform 1 0 56640 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input63
timestamp 1621261055
transform 1 0 57408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input69
timestamp 1621261055
transform 1 0 55872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_574
timestamp 1621261055
transform 1 0 56256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_579
timestamp 1621261055
transform 1 0 56736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_583
timestamp 1621261055
transform 1 0 57120 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_585
timestamp 1621261055
transform 1 0 57312 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_9
timestamp 1621261055
transform -1 0 58848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_590
timestamp 1621261055
transform 1 0 57792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_594
timestamp 1621261055
transform 1 0 58176 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_596
timestamp 1621261055
transform 1 0 58368 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_10
timestamp 1621261055
transform 1 0 1152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input357
timestamp 1621261055
transform 1 0 3168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input363
timestamp 1621261055
transform 1 0 1536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input364
timestamp 1621261055
transform 1 0 2304 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_8
timestamp 1621261055
transform 1 0 1920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_16
timestamp 1621261055
transform 1 0 2688 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_20
timestamp 1621261055
transform 1 0 3072 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input359
timestamp 1621261055
transform 1 0 3936 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input361
timestamp 1621261055
transform 1 0 4704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_25
timestamp 1621261055
transform 1 0 3552 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_33
timestamp 1621261055
transform 1 0 4320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_41
timestamp 1621261055
transform 1 0 5088 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_227
timestamp 1621261055
transform 1 0 6432 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output575
timestamp 1621261055
transform 1 0 5472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output577
timestamp 1621261055
transform 1 0 6912 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_216
timestamp 1621261055
transform 1 0 5280 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_218
timestamp 1621261055
transform 1 0 6720 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_49
timestamp 1621261055
transform 1 0 5856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_53
timestamp 1621261055
transform 1 0 6240 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_56
timestamp 1621261055
transform 1 0 6528 0 1 5994
box -38 -49 230 715
use AND2X2  AND2X2
timestamp 1624196784
transform 1 0 7680 0 1 5994
box 0 -48 1152 714
use sky130_fd_sc_ls__diode_2  ANTENNA_99
timestamp 1621261055
transform 1 0 7488 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_64
timestamp 1621261055
transform 1 0 7296 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_80
timestamp 1621261055
transform 1 0 8832 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_84
timestamp 1621261055
transform 1 0 9216 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input344
timestamp 1621261055
transform 1 0 9408 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input346
timestamp 1621261055
transform 1 0 10176 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input348
timestamp 1621261055
transform 1 0 10944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_90
timestamp 1621261055
transform 1 0 9792 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_98
timestamp 1621261055
transform 1 0 10560 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_228
timestamp 1621261055
transform 1 0 11712 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input350
timestamp 1621261055
transform 1 0 12192 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input353
timestamp 1621261055
transform 1 0 12960 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_106
timestamp 1621261055
transform 1 0 11328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_111
timestamp 1621261055
transform 1 0 11808 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_119
timestamp 1621261055
transform 1 0 12576 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output444
timestamp 1621261055
transform 1 0 13728 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output494
timestamp 1621261055
transform 1 0 14496 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output505
timestamp 1621261055
transform 1 0 15264 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_173
timestamp 1621261055
transform 1 0 15072 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_127
timestamp 1621261055
transform 1 0 13344 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_135
timestamp 1621261055
transform 1 0 14112 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_143
timestamp 1621261055
transform 1 0 14880 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_229
timestamp 1621261055
transform 1 0 16992 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output527
timestamp 1621261055
transform -1 0 16416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_111
timestamp 1621261055
transform 1 0 17280 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_186
timestamp 1621261055
transform -1 0 16032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_151
timestamp 1621261055
transform 1 0 15648 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_159
timestamp 1621261055
transform 1 0 16416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_163
timestamp 1621261055
transform 1 0 16800 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_166
timestamp 1621261055
transform 1 0 17088 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output455
timestamp 1621261055
transform 1 0 17472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output475
timestamp 1621261055
transform 1 0 18240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output477
timestamp 1621261055
transform 1 0 19008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_131
timestamp 1621261055
transform 1 0 18048 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_135
timestamp 1621261055
transform 1 0 18816 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_174
timestamp 1621261055
transform 1 0 17856 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_182
timestamp 1621261055
transform 1 0 18624 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output479
timestamp 1621261055
transform 1 0 19776 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output480
timestamp 1621261055
transform 1 0 20544 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output482
timestamp 1621261055
transform 1 0 21312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_137
timestamp 1621261055
transform 1 0 20352 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_190
timestamp 1621261055
transform 1 0 19392 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_198
timestamp 1621261055
transform 1 0 20160 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_206
timestamp 1621261055
transform 1 0 20928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_230
timestamp 1621261055
transform 1 0 22272 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output487
timestamp 1621261055
transform 1 0 22752 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_145
timestamp 1621261055
transform -1 0 23520 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_214
timestamp 1621261055
transform 1 0 21696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_218
timestamp 1621261055
transform 1 0 22080 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_221
timestamp 1621261055
transform 1 0 22368 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_229
timestamp 1621261055
transform 1 0 23136 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output489
timestamp 1621261055
transform -1 0 23904 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output491
timestamp 1621261055
transform -1 0 24672 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_149
timestamp 1621261055
transform -1 0 24288 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_237
timestamp 1621261055
transform 1 0 23904 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_245
timestamp 1621261055
transform 1 0 24672 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input222
timestamp 1621261055
transform 1 0 25632 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input225
timestamp 1621261055
transform 1 0 26784 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_253
timestamp 1621261055
transform 1 0 25440 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_259
timestamp 1621261055
transform 1 0 26016 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_5_271
timestamp 1621261055
transform 1 0 27168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_231
timestamp 1621261055
transform 1 0 27552 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output501
timestamp 1621261055
transform -1 0 28416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output504
timestamp 1621261055
transform 1 0 28800 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_167
timestamp 1621261055
transform -1 0 28032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_171
timestamp 1621261055
transform 1 0 28608 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_276
timestamp 1621261055
transform 1 0 27648 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_284
timestamp 1621261055
transform 1 0 28416 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_292
timestamp 1621261055
transform 1 0 29184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input234
timestamp 1621261055
transform 1 0 29664 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input238
timestamp 1621261055
transform 1 0 31200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output509
timestamp 1621261055
transform 1 0 30432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_296
timestamp 1621261055
transform 1 0 29568 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_301
timestamp 1621261055
transform 1 0 30048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_309
timestamp 1621261055
transform 1 0 30816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_232
timestamp 1621261055
transform 1 0 32832 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output513
timestamp 1621261055
transform 1 0 31968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output518
timestamp 1621261055
transform -1 0 33696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_183
timestamp 1621261055
transform -1 0 33312 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_317
timestamp 1621261055
transform 1 0 31584 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_325
timestamp 1621261055
transform 1 0 32352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_329
timestamp 1621261055
transform 1 0 32736 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_331
timestamp 1621261055
transform 1 0 32928 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output520
timestamp 1621261055
transform 1 0 34080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output522
timestamp 1621261055
transform -1 0 35232 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_184
timestamp 1621261055
transform -1 0 34848 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_339
timestamp 1621261055
transform 1 0 33696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_347
timestamp 1621261055
transform 1 0 34464 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_355
timestamp 1621261055
transform 1 0 35232 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _115_
timestamp 1621261055
transform 1 0 35616 0 1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input254
timestamp 1621261055
transform 1 0 36288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output529
timestamp 1621261055
transform -1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_187
timestamp 1621261055
transform -1 0 37056 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_362
timestamp 1621261055
transform 1 0 35904 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_370
timestamp 1621261055
transform 1 0 36672 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_378
timestamp 1621261055
transform 1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_233
timestamp 1621261055
transform 1 0 38112 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input262
timestamp 1621261055
transform 1 0 38880 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_382
timestamp 1621261055
transform 1 0 37824 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_384
timestamp 1621261055
transform 1 0 38016 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_386
timestamp 1621261055
transform 1 0 38208 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_390
timestamp 1621261055
transform 1 0 38592 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_392
timestamp 1621261055
transform 1 0 38784 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_5_397
timestamp 1621261055
transform 1 0 39264 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input266
timestamp 1621261055
transform 1 0 40320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output540
timestamp 1621261055
transform -1 0 41472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_196
timestamp 1621261055
transform -1 0 41088 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_405
timestamp 1621261055
transform 1 0 40032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_407
timestamp 1621261055
transform 1 0 40224 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_412
timestamp 1621261055
transform 1 0 40704 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_420
timestamp 1621261055
transform 1 0 41472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_234
timestamp 1621261055
transform 1 0 43392 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input270
timestamp 1621261055
transform 1 0 41856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output544
timestamp 1621261055
transform 1 0 42624 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_428
timestamp 1621261055
transform 1 0 42240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_436
timestamp 1621261055
transform 1 0 43008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_441
timestamp 1621261055
transform 1 0 43488 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input281
timestamp 1621261055
transform 1 0 45504 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output548
timestamp 1621261055
transform 1 0 43872 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output552
timestamp 1621261055
transform 1 0 44640 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_449
timestamp 1621261055
transform 1 0 44256 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_457
timestamp 1621261055
transform 1 0 45024 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_461
timestamp 1621261055
transform 1 0 45408 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input286
timestamp 1621261055
transform 1 0 46944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_466
timestamp 1621261055
transform 1 0 45888 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_474
timestamp 1621261055
transform 1 0 46656 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_476
timestamp 1621261055
transform 1 0 46848 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_481
timestamp 1621261055
transform 1 0 47328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_235
timestamp 1621261055
transform 1 0 48672 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input288
timestamp 1621261055
transform 1 0 47712 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input291
timestamp 1621261055
transform 1 0 49152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_489
timestamp 1621261055
transform 1 0 48096 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_493
timestamp 1621261055
transform 1 0 48480 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_496
timestamp 1621261055
transform 1 0 48768 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_504
timestamp 1621261055
transform 1 0 49536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input293
timestamp 1621261055
transform 1 0 49920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output445
timestamp 1621261055
transform -1 0 51072 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output447
timestamp 1621261055
transform -1 0 51840 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_105
timestamp 1621261055
transform -1 0 50688 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_107
timestamp 1621261055
transform -1 0 51456 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_512
timestamp 1621261055
transform 1 0 50304 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_520
timestamp 1621261055
transform 1 0 51072 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input192
timestamp 1621261055
transform 1 0 53184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output448
timestamp 1621261055
transform 1 0 52224 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_528
timestamp 1621261055
transform 1 0 51840 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_536
timestamp 1621261055
transform 1 0 52608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_540
timestamp 1621261055
transform 1 0 52992 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_546
timestamp 1621261055
transform 1 0 53568 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_236
timestamp 1621261055
transform 1 0 53952 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input180
timestamp 1621261055
transform 1 0 54432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input181
timestamp 1621261055
transform 1 0 55200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_551
timestamp 1621261055
transform 1 0 54048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_559
timestamp 1621261055
transform 1 0 54816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_567
timestamp 1621261055
transform 1 0 55584 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input67
timestamp 1621261055
transform 1 0 56928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input183
timestamp 1621261055
transform 1 0 55968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_575
timestamp 1621261055
transform 1 0 56352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_579
timestamp 1621261055
transform 1 0 56736 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_585
timestamp 1621261055
transform 1 0 57312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_11
timestamp 1621261055
transform -1 0 58848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input65
timestamp 1621261055
transform 1 0 57696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_593
timestamp 1621261055
transform 1 0 58080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_12
timestamp 1621261055
transform 1 0 1152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input365
timestamp 1621261055
transform 1 0 2496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input366
timestamp 1621261055
transform 1 0 1536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_8
timestamp 1621261055
transform 1 0 1920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_12
timestamp 1621261055
transform 1 0 2304 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_18
timestamp 1621261055
transform 1 0 2880 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_237
timestamp 1621261055
transform 1 0 3840 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output598
timestamp 1621261055
transform 1 0 4320 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output601
timestamp 1621261055
transform 1 0 5088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_234
timestamp 1621261055
transform 1 0 4128 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_26
timestamp 1621261055
transform 1 0 3648 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_29
timestamp 1621261055
transform 1 0 3936 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_37
timestamp 1621261055
transform 1 0 4704 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output576
timestamp 1621261055
transform 1 0 5856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output578
timestamp 1621261055
transform 1 0 6624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_220
timestamp 1621261055
transform 1 0 6432 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_45
timestamp 1621261055
transform 1 0 5472 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_53
timestamp 1621261055
transform 1 0 6240 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_61
timestamp 1621261055
transform 1 0 7008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_238
timestamp 1621261055
transform 1 0 9120 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output579
timestamp 1621261055
transform 1 0 7392 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output580
timestamp 1621261055
transform 1 0 8160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_69
timestamp 1621261055
transform 1 0 7776 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_77
timestamp 1621261055
transform 1 0 8544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_81
timestamp 1621261055
transform 1 0 8928 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_84
timestamp 1621261055
transform 1 0 9216 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input349
timestamp 1621261055
transform 1 0 11232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output582
timestamp 1621261055
transform 1 0 9600 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output585
timestamp 1621261055
transform 1 0 10368 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_222
timestamp 1621261055
transform 1 0 10176 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_92
timestamp 1621261055
transform 1 0 9984 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_100
timestamp 1621261055
transform 1 0 10752 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_104
timestamp 1621261055
transform 1 0 11136 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input354
timestamp 1621261055
transform 1 0 12672 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_109
timestamp 1621261055
transform 1 0 11616 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_117
timestamp 1621261055
transform 1 0 12384 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_119
timestamp 1621261055
transform 1 0 12576 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_124
timestamp 1621261055
transform 1 0 13056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_239
timestamp 1621261055
transform 1 0 14400 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output483
timestamp 1621261055
transform 1 0 13440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output516
timestamp 1621261055
transform -1 0 15264 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_181
timestamp 1621261055
transform -1 0 14880 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_132
timestamp 1621261055
transform 1 0 13824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_136
timestamp 1621261055
transform 1 0 14208 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_139
timestamp 1621261055
transform 1 0 14496 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_147
timestamp 1621261055
transform 1 0 15264 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _042_
timestamp 1621261055
transform 1 0 16416 0 -1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output466
timestamp 1621261055
transform 1 0 17088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output538
timestamp 1621261055
transform 1 0 15648 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_43
timestamp 1621261055
transform 1 0 16224 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_155
timestamp 1621261055
transform 1 0 16032 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_162
timestamp 1621261055
transform 1 0 16704 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output476
timestamp 1621261055
transform 1 0 17856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output478
timestamp 1621261055
transform 1 0 18624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_133
timestamp 1621261055
transform 1 0 17664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_170
timestamp 1621261055
transform 1 0 17472 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_178
timestamp 1621261055
transform 1 0 18240 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_186
timestamp 1621261055
transform 1 0 19008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_240
timestamp 1621261055
transform 1 0 19680 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output481
timestamp 1621261055
transform -1 0 20544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output484
timestamp 1621261055
transform 1 0 20928 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_139
timestamp 1621261055
transform -1 0 20160 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_190
timestamp 1621261055
transform 1 0 19392 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_192
timestamp 1621261055
transform 1 0 19584 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_194
timestamp 1621261055
transform 1 0 19776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_202
timestamp 1621261055
transform 1 0 20544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_210
timestamp 1621261055
transform 1 0 21312 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output486
timestamp 1621261055
transform 1 0 21696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output488
timestamp 1621261055
transform 1 0 22464 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output490
timestamp 1621261055
transform -1 0 23616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_141
timestamp 1621261055
transform 1 0 21504 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_143
timestamp 1621261055
transform 1 0 22272 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_147
timestamp 1621261055
transform -1 0 23232 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_218
timestamp 1621261055
transform 1 0 22080 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_226
timestamp 1621261055
transform 1 0 22848 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_241
timestamp 1621261055
transform 1 0 24960 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output492
timestamp 1621261055
transform -1 0 24384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_151
timestamp 1621261055
transform -1 0 24000 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_157
timestamp 1621261055
transform 1 0 25248 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_234
timestamp 1621261055
transform 1 0 23616 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_242
timestamp 1621261055
transform 1 0 24384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_246
timestamp 1621261055
transform 1 0 24768 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_249
timestamp 1621261055
transform 1 0 25056 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output496
timestamp 1621261055
transform 1 0 25440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output498
timestamp 1621261055
transform 1 0 26208 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output500
timestamp 1621261055
transform -1 0 27360 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_161
timestamp 1621261055
transform 1 0 26016 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_165
timestamp 1621261055
transform -1 0 26976 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_257
timestamp 1621261055
transform 1 0 25824 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_265
timestamp 1621261055
transform 1 0 26592 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_273
timestamp 1621261055
transform 1 0 27360 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output503
timestamp 1621261055
transform 1 0 27744 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output506
timestamp 1621261055
transform 1 0 28512 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output508
timestamp 1621261055
transform 1 0 29280 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_169
timestamp 1621261055
transform 1 0 27552 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_281
timestamp 1621261055
transform 1 0 28128 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_289
timestamp 1621261055
transform 1 0 28896 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_242
timestamp 1621261055
transform 1 0 30240 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output512
timestamp 1621261055
transform -1 0 31104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_177
timestamp 1621261055
transform -1 0 30720 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_179
timestamp 1621261055
transform -1 0 31488 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_297
timestamp 1621261055
transform 1 0 29664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_301
timestamp 1621261055
transform 1 0 30048 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_304
timestamp 1621261055
transform 1 0 30336 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_312
timestamp 1621261055
transform 1 0 31104 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output514
timestamp 1621261055
transform -1 0 31872 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output517
timestamp 1621261055
transform 1 0 32256 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output519
timestamp 1621261055
transform 1 0 33024 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_320
timestamp 1621261055
transform 1 0 31872 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_328
timestamp 1621261055
transform 1 0 32640 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_336
timestamp 1621261055
transform 1 0 33408 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output521
timestamp 1621261055
transform 1 0 33792 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output524
timestamp 1621261055
transform 1 0 34560 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_344
timestamp 1621261055
transform 1 0 34176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_352
timestamp 1621261055
transform 1 0 34944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_356
timestamp 1621261055
transform 1 0 35328 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_243
timestamp 1621261055
transform 1 0 35520 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output528
timestamp 1621261055
transform 1 0 36000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output531
timestamp 1621261055
transform 1 0 36768 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_359
timestamp 1621261055
transform 1 0 35616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_367
timestamp 1621261055
transform 1 0 36384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_375
timestamp 1621261055
transform 1 0 37152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output533
timestamp 1621261055
transform 1 0 37536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output534
timestamp 1621261055
transform -1 0 38688 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output535
timestamp 1621261055
transform 1 0 39072 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_191
timestamp 1621261055
transform -1 0 38304 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_383
timestamp 1621261055
transform 1 0 37920 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_391
timestamp 1621261055
transform 1 0 38688 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_399
timestamp 1621261055
transform 1 0 39456 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_244
timestamp 1621261055
transform 1 0 40800 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output537
timestamp 1621261055
transform -1 0 40224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output542
timestamp 1621261055
transform 1 0 41280 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_193
timestamp 1621261055
transform -1 0 39840 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_407
timestamp 1621261055
transform 1 0 40224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_411
timestamp 1621261055
transform 1 0 40608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_414
timestamp 1621261055
transform 1 0 40896 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output545
timestamp 1621261055
transform -1 0 42432 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output547
timestamp 1621261055
transform 1 0 42816 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_200
timestamp 1621261055
transform -1 0 42048 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_203
timestamp 1621261055
transform -1 0 43584 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_422
timestamp 1621261055
transform 1 0 41664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_430
timestamp 1621261055
transform 1 0 42432 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_438
timestamp 1621261055
transform 1 0 43200 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output551
timestamp 1621261055
transform -1 0 43968 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output553
timestamp 1621261055
transform -1 0 44736 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output555
timestamp 1621261055
transform -1 0 45504 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_204
timestamp 1621261055
transform -1 0 44352 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_205
timestamp 1621261055
transform -1 0 45120 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_446
timestamp 1621261055
transform 1 0 43968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_454
timestamp 1621261055
transform 1 0 44736 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_462
timestamp 1621261055
transform 1 0 45504 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_245
timestamp 1621261055
transform 1 0 46080 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output558
timestamp 1621261055
transform 1 0 46560 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output561
timestamp 1621261055
transform 1 0 47328 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_466
timestamp 1621261055
transform 1 0 45888 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_469
timestamp 1621261055
transform 1 0 46176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_477
timestamp 1621261055
transform 1 0 46944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output563
timestamp 1621261055
transform 1 0 48096 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output565
timestamp 1621261055
transform 1 0 48864 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_485
timestamp 1621261055
transform 1 0 47712 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_493
timestamp 1621261055
transform 1 0 48480 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_501
timestamp 1621261055
transform 1 0 49248 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_246
timestamp 1621261055
transform 1 0 51360 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output446
timestamp 1621261055
transform 1 0 50112 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_509
timestamp 1621261055
transform 1 0 50016 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_6_514
timestamp 1621261055
transform 1 0 50496 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_6_522
timestamp 1621261055
transform 1 0 51264 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_524
timestamp 1621261055
transform 1 0 51456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output449
timestamp 1621261055
transform 1 0 51840 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output451
timestamp 1621261055
transform 1 0 52608 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_532
timestamp 1621261055
transform 1 0 52224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_540
timestamp 1621261055
transform 1 0 52992 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input182
timestamp 1621261055
transform 1 0 54720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input184
timestamp 1621261055
transform 1 0 55488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input196
timestamp 1621261055
transform 1 0 53952 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_548
timestamp 1621261055
transform 1 0 53760 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_554
timestamp 1621261055
transform 1 0 54336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_562
timestamp 1621261055
transform 1 0 55104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_247
timestamp 1621261055
transform 1 0 56640 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_6_570
timestamp 1621261055
transform 1 0 55872 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_6_579
timestamp 1621261055
transform 1 0 56736 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_587
timestamp 1621261055
transform 1 0 57504 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_13
timestamp 1621261055
transform -1 0 58848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input66
timestamp 1621261055
transform 1 0 57696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_593
timestamp 1621261055
transform 1 0 58080 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output572
timestamp 1621261055
transform 1 0 1536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input367
timestamp 1621261055
transform 1 0 1536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_16
timestamp 1621261055
transform 1 0 1152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_14
timestamp 1621261055
transform 1 0 1152 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_8
timestamp 1621261055
transform 1 0 1920 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_212
timestamp 1621261055
transform 1 0 1920 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_10
timestamp 1621261055
transform 1 0 2112 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output584
timestamp 1621261055
transform 1 0 2304 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output573
timestamp 1621261055
transform 1 0 2304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_16
timestamp 1621261055
transform 1 0 2688 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_16
timestamp 1621261055
transform 1 0 2688 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_236
timestamp 1621261055
transform 1 0 2880 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_232
timestamp 1621261055
transform 1 0 2880 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output599
timestamp 1621261055
transform 1 0 3072 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output595
timestamp 1621261055
transform 1 0 3072 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_29
timestamp 1621261055
transform 1 0 3936 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_24
timestamp 1621261055
transform 1 0 3456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_24
timestamp 1621261055
transform 1 0 3456 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output600
timestamp 1621261055
transform 1 0 3840 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_258
timestamp 1621261055
transform 1 0 3840 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_37
timestamp 1621261055
transform 1 0 4704 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_32
timestamp 1621261055
transform 1 0 4224 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_238
timestamp 1621261055
transform 1 0 4128 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output603
timestamp 1621261055
transform 1 0 4320 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output602
timestamp 1621261055
transform 1 0 4608 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_40
timestamp 1621261055
transform 1 0 4992 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_240
timestamp 1621261055
transform 1 0 5184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_45
timestamp 1621261055
transform 1 0 5472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output604
timestamp 1621261055
transform 1 0 5376 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_49
timestamp 1621261055
transform 1 0 5856 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_48
timestamp 1621261055
transform 1 0 5760 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _139_
timestamp 1621261055
transform 1 0 5952 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_8_53
timestamp 1621261055
transform 1 0 6240 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_56
timestamp 1621261055
transform 1 0 6528 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_54
timestamp 1621261055
transform 1 0 6336 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_52
timestamp 1621261055
transform 1 0 6144 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_248
timestamp 1621261055
transform 1 0 6432 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_61
timestamp 1621261055
transform 1 0 7008 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_57
timestamp 1621261055
transform 1 0 6624 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _202_
timestamp 1621261055
transform 1 0 6720 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _119_
timestamp 1621261055
transform 1 0 6912 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_63
timestamp 1621261055
transform 1 0 7200 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_72
timestamp 1621261055
transform 1 0 8064 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_67
timestamp 1621261055
transform 1 0 7584 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_65
timestamp 1621261055
transform 1 0 7392 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_7_65
timestamp 1621261055
transform 1 0 7392 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_103
timestamp 1621261055
transform 1 0 7488 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output581
timestamp 1621261055
transform 1 0 7680 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_84
timestamp 1621261055
transform 1 0 9216 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_82
timestamp 1621261055
transform 1 0 9024 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_80
timestamp 1621261055
transform 1 0 8832 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_80
timestamp 1621261055
transform 1 0 8832 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output583
timestamp 1621261055
transform 1 0 9216 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_259
timestamp 1621261055
transform 1 0 9120 0 -1 8658
box -38 -49 134 715
use AOI21X1  AOI21X1
timestamp 1624196784
transform 1 0 7680 0 1 7326
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_4  FILLER_7_88
timestamp 1621261055
transform 1 0 9600 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_224
timestamp 1621261055
transform 1 0 9408 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output587
timestamp 1621261055
transform 1 0 9600 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_92
timestamp 1621261055
transform 1 0 9984 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output586
timestamp 1621261055
transform 1 0 9984 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_96
timestamp 1621261055
transform 1 0 10368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output589
timestamp 1621261055
transform 1 0 10368 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_100
timestamp 1621261055
transform 1 0 10752 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_226
timestamp 1621261055
transform 1 0 10944 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output588
timestamp 1621261055
transform 1 0 10752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_104
timestamp 1621261055
transform 1 0 11136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output590
timestamp 1621261055
transform 1 0 11136 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_108
timestamp 1621261055
transform 1 0 11520 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_108
timestamp 1621261055
transform 1 0 11520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_111
timestamp 1621261055
transform 1 0 11808 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_228
timestamp 1621261055
transform 1 0 11712 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output592
timestamp 1621261055
transform 1 0 11904 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_249
timestamp 1621261055
transform 1 0 11712 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_116
timestamp 1621261055
transform 1 0 12288 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_119
timestamp 1621261055
transform 1 0 12576 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output591
timestamp 1621261055
transform 1 0 12192 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_124
timestamp 1621261055
transform 1 0 13056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_230
timestamp 1621261055
transform 1 0 12768 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output594
timestamp 1621261055
transform 1 0 12672 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output593
timestamp 1621261055
transform 1 0 12960 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_132
timestamp 1621261055
transform 1 0 13824 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_127
timestamp 1621261055
transform 1 0 13344 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output597
timestamp 1621261055
transform 1 0 13440 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output596
timestamp 1621261055
transform 1 0 13728 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_139
timestamp 1621261055
transform 1 0 14496 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_136
timestamp 1621261055
transform 1 0 14208 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_7_143
timestamp 1621261055
transform 1 0 14880 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_7_135
timestamp 1621261055
transform 1 0 14112 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_260
timestamp 1621261055
transform 1 0 14400 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_147
timestamp 1621261055
transform 1 0 15264 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_147
timestamp 1621261055
transform 1 0 15264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _098_
timestamp 1621261055
transform 1 0 14976 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_7_155
timestamp 1621261055
transform 1 0 16032 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_202
timestamp 1621261055
transform 1 0 15456 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output560
timestamp 1621261055
transform 1 0 16032 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output549
timestamp 1621261055
transform 1 0 15648 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_159
timestamp 1621261055
transform 1 0 16416 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_163
timestamp 1621261055
transform 1 0 16800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output571
timestamp 1621261055
transform 1 0 16800 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_167
timestamp 1621261055
transform 1 0 17184 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_166
timestamp 1621261055
transform 1 0 17088 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_250
timestamp 1621261055
transform 1 0 16992 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _125_
timestamp 1621261055
transform 1 0 17568 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_7_174
timestamp 1621261055
transform 1 0 17856 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_182
timestamp 1621261055
transform 1 0 18624 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_174
timestamp 1621261055
transform 1 0 17856 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_182
timestamp 1621261055
transform 1 0 18624 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_194
timestamp 1621261055
transform 1 0 19776 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_192
timestamp 1621261055
transform 1 0 19584 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_190
timestamp 1621261055
transform 1 0 19392 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_190
timestamp 1621261055
transform 1 0 19392 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_261
timestamp 1621261055
transform 1 0 19680 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_202
timestamp 1621261055
transform 1 0 20544 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_202
timestamp 1621261055
transform 1 0 20544 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_198
timestamp 1621261055
transform 1 0 20160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output485
timestamp 1621261055
transform 1 0 20736 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_210
timestamp 1621261055
transform 1 0 21312 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_208
timestamp 1621261055
transform 1 0 21120 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_214
timestamp 1621261055
transform 1 0 21696 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_215
timestamp 1621261055
transform 1 0 21792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _199_
timestamp 1621261055
transform 1 0 21504 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _148_
timestamp 1621261055
transform 1 0 21888 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_227
timestamp 1621261055
transform 1 0 22944 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_219
timestamp 1621261055
transform 1 0 22176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_227
timestamp 1621261055
transform 1 0 22944 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_225
timestamp 1621261055
transform 1 0 22752 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_221
timestamp 1621261055
transform 1 0 22368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_219
timestamp 1621261055
transform 1 0 22176 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_251
timestamp 1621261055
transform 1 0 22272 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_231
timestamp 1621261055
transform 1 0 23328 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _103_
timestamp 1621261055
transform 1 0 23040 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_235
timestamp 1621261055
transform 1 0 23712 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_239
timestamp 1621261055
transform 1 0 24096 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_153
timestamp 1621261055
transform 1 0 23520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output493
timestamp 1621261055
transform 1 0 23712 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_247
timestamp 1621261055
transform 1 0 24864 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_243
timestamp 1621261055
transform 1 0 24480 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_247
timestamp 1621261055
transform 1 0 24864 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_155
timestamp 1621261055
transform -1 0 24480 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output495
timestamp 1621261055
transform -1 0 24864 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_262
timestamp 1621261055
transform 1 0 24960 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_249
timestamp 1621261055
transform 1 0 25056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_159
timestamp 1621261055
transform 1 0 25056 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output497
timestamp 1621261055
transform 1 0 25248 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_259
timestamp 1621261055
transform 1 0 26016 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_255
timestamp 1621261055
transform 1 0 25632 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_253
timestamp 1621261055
transform 1 0 25440 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_255
timestamp 1621261055
transform 1 0 25632 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_163
timestamp 1621261055
transform -1 0 26016 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output499
timestamp 1621261055
transform -1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _110_
timestamp 1621261055
transform 1 0 25728 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_267
timestamp 1621261055
transform 1 0 26784 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_263
timestamp 1621261055
transform 1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output502
timestamp 1621261055
transform 1 0 26784 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_271
timestamp 1621261055
transform 1 0 27168 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_275
timestamp 1621261055
transform 1 0 27552 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_280
timestamp 1621261055
transform 1 0 28032 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_276
timestamp 1621261055
transform 1 0 27648 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output507
timestamp 1621261055
transform 1 0 28128 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_252
timestamp 1621261055
transform 1 0 27552 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_283
timestamp 1621261055
transform 1 0 28320 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_289
timestamp 1621261055
transform 1 0 28896 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_285
timestamp 1621261055
transform 1 0 28512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_175
timestamp 1621261055
transform -1 0 29184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_291
timestamp 1621261055
transform 1 0 29088 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output510
timestamp 1621261055
transform -1 0 29568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_299
timestamp 1621261055
transform 1 0 29856 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_296
timestamp 1621261055
transform 1 0 29568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output511
timestamp 1621261055
transform 1 0 29952 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_304
timestamp 1621261055
transform 1 0 30336 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_310
timestamp 1621261055
transform 1 0 30912 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_308
timestamp 1621261055
transform 1 0 30720 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_304
timestamp 1621261055
transform 1 0 30336 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output515
timestamp 1621261055
transform 1 0 31008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_263
timestamp 1621261055
transform 1 0 30240 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_312
timestamp 1621261055
transform 1 0 31104 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_315
timestamp 1621261055
transform 1 0 31392 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _151_
timestamp 1621261055
transform 1 0 32160 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _204_
timestamp 1621261055
transform 1 0 33408 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_253
timestamp 1621261055
transform 1 0 32832 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_326
timestamp 1621261055
transform 1 0 32448 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_331
timestamp 1621261055
transform 1 0 32928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_335
timestamp 1621261055
transform 1 0 33312 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_320
timestamp 1621261055
transform 1 0 31872 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_328
timestamp 1621261055
transform 1 0 32640 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_339
timestamp 1621261055
transform 1 0 33696 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_7_337
timestamp 1621261055
transform 1 0 33504 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output523
timestamp 1621261055
transform 1 0 33600 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_341
timestamp 1621261055
transform 1 0 33888 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_342
timestamp 1621261055
transform 1 0 33984 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_21
timestamp 1621261055
transform -1 0 34176 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _011_
timestamp 1621261055
transform -1 0 34464 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_8_347
timestamp 1621261055
transform 1 0 34464 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_350
timestamp 1621261055
transform 1 0 34752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output525
timestamp 1621261055
transform 1 0 34368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_354
timestamp 1621261055
transform 1 0 35136 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output526
timestamp 1621261055
transform 1 0 35136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _171_
timestamp 1621261055
transform 1 0 34848 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_359
timestamp 1621261055
transform 1 0 35616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_358
timestamp 1621261055
transform 1 0 35520 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output530
timestamp 1621261055
transform 1 0 35904 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_264
timestamp 1621261055
transform 1 0 35520 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_367
timestamp 1621261055
transform 1 0 36384 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_374
timestamp 1621261055
transform 1 0 37056 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_366
timestamp 1621261055
transform 1 0 36288 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_189
timestamp 1621261055
transform -1 0 36672 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output532
timestamp 1621261055
transform -1 0 37056 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_375
timestamp 1621261055
transform 1 0 37152 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_383
timestamp 1621261055
transform 1 0 37920 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_386
timestamp 1621261055
transform 1 0 38208 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_384
timestamp 1621261055
transform 1 0 38016 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_382
timestamp 1621261055
transform 1 0 37824 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_254
timestamp 1621261055
transform 1 0 38112 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_391
timestamp 1621261055
transform 1 0 38688 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_394
timestamp 1621261055
transform 1 0 38976 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output536
timestamp 1621261055
transform 1 0 38592 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_239
timestamp 1621261055
transform -1 0 39648 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_195
timestamp 1621261055
transform -1 0 39360 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output539
timestamp 1621261055
transform -1 0 39744 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_404
timestamp 1621261055
transform 1 0 39936 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_402
timestamp 1621261055
transform 1 0 39744 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_198
timestamp 1621261055
transform -1 0 40128 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output541
timestamp 1621261055
transform -1 0 40512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _196_
timestamp 1621261055
transform -1 0 39936 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_414
timestamp 1621261055
transform 1 0 40896 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_412
timestamp 1621261055
transform 1 0 40704 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_410
timestamp 1621261055
transform 1 0 40512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output543
timestamp 1621261055
transform 1 0 40896 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_265
timestamp 1621261055
transform 1 0 40800 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_418
timestamp 1621261055
transform 1 0 41280 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_424
timestamp 1621261055
transform 1 0 41856 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_422
timestamp 1621261055
transform 1 0 41664 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_426
timestamp 1621261055
transform 1 0 42048 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_39
timestamp 1621261055
transform -1 0 42144 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output546
timestamp 1621261055
transform 1 0 41664 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _041_
timestamp 1621261055
transform -1 0 42432 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_430
timestamp 1621261055
transform 1 0 42432 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_434
timestamp 1621261055
transform 1 0 42816 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output550
timestamp 1621261055
transform 1 0 42432 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_438
timestamp 1621261055
transform 1 0 43200 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_441
timestamp 1621261055
transform 1 0 43488 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_438
timestamp 1621261055
transform 1 0 43200 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_255
timestamp 1621261055
transform 1 0 43392 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output554
timestamp 1621261055
transform 1 0 43872 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output556
timestamp 1621261055
transform 1 0 44640 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output557
timestamp 1621261055
transform 1 0 45408 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_449
timestamp 1621261055
transform 1 0 44256 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_457
timestamp 1621261055
transform 1 0 45024 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_446
timestamp 1621261055
transform 1 0 43968 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_454
timestamp 1621261055
transform 1 0 44736 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_8_462
timestamp 1621261055
transform 1 0 45504 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_469
timestamp 1621261055
transform 1 0 46176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_466
timestamp 1621261055
transform 1 0 45888 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_465
timestamp 1621261055
transform 1 0 45792 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_207
timestamp 1621261055
transform 1 0 45984 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output559
timestamp 1621261055
transform 1 0 46176 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_266
timestamp 1621261055
transform 1 0 46080 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_477
timestamp 1621261055
transform 1 0 46944 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_473
timestamp 1621261055
transform 1 0 46560 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_209
timestamp 1621261055
transform 1 0 46752 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output562
timestamp 1621261055
transform 1 0 46944 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_481
timestamp 1621261055
transform 1 0 47328 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_487
timestamp 1621261055
transform 1 0 47904 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_485
timestamp 1621261055
transform 1 0 47712 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output566
timestamp 1621261055
transform 1 0 48000 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output564
timestamp 1621261055
transform 1 0 47712 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_492
timestamp 1621261055
transform 1 0 48384 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_489
timestamp 1621261055
transform 1 0 48096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_496
timestamp 1621261055
transform 1 0 48768 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_493
timestamp 1621261055
transform 1 0 48480 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_210
timestamp 1621261055
transform -1 0 48768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output568
timestamp 1621261055
transform -1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_256
timestamp 1621261055
transform 1 0 48672 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_500
timestamp 1621261055
transform 1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output567
timestamp 1621261055
transform 1 0 49152 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_504
timestamp 1621261055
transform 1 0 49536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output570
timestamp 1621261055
transform 1 0 49536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_508
timestamp 1621261055
transform 1 0 49920 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_512
timestamp 1621261055
transform 1 0 50304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output569
timestamp 1621261055
transform 1 0 49920 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_520
timestamp 1621261055
transform 1 0 51072 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_516
timestamp 1621261055
transform 1 0 50688 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_516
timestamp 1621261055
transform 1 0 50688 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output473
timestamp 1621261055
transform 1 0 50880 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_524
timestamp 1621261055
transform 1 0 51456 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_522
timestamp 1621261055
transform 1 0 51264 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_522
timestamp 1621261055
transform 1 0 51264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_109
timestamp 1621261055
transform -1 0 51648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_267
timestamp 1621261055
transform 1 0 51360 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_530
timestamp 1621261055
transform 1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output450
timestamp 1621261055
transform -1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_532
timestamp 1621261055
transform 1 0 52224 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output472
timestamp 1621261055
transform 1 0 52320 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output452
timestamp 1621261055
transform 1 0 52416 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_537
timestamp 1621261055
transform 1 0 52704 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_538
timestamp 1621261055
transform 1 0 52800 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output454
timestamp 1621261055
transform 1 0 53088 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output453
timestamp 1621261055
transform 1 0 53184 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_545
timestamp 1621261055
transform 1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_546
timestamp 1621261055
transform 1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_553
timestamp 1621261055
transform 1 0 54240 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_551
timestamp 1621261055
transform 1 0 54048 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output456
timestamp 1621261055
transform 1 0 53856 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_257
timestamp 1621261055
transform 1 0 53952 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_561
timestamp 1621261055
transform 1 0 55008 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_559
timestamp 1621261055
transform 1 0 54816 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input197
timestamp 1621261055
transform 1 0 55104 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input194
timestamp 1621261055
transform 1 0 55008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_566
timestamp 1621261055
transform 1 0 55488 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_565
timestamp 1621261055
transform 1 0 55392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_574
timestamp 1621261055
transform 1 0 56256 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_573
timestamp 1621261055
transform 1 0 56160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input193
timestamp 1621261055
transform 1 0 55872 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input185
timestamp 1621261055
transform 1 0 55776 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_579
timestamp 1621261055
transform 1 0 56736 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_581
timestamp 1621261055
transform 1 0 56928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input188
timestamp 1621261055
transform 1 0 57120 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input186
timestamp 1621261055
transform 1 0 56544 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_268
timestamp 1621261055
transform 1 0 56640 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_587
timestamp 1621261055
transform 1 0 57504 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input187
timestamp 1621261055
transform 1 0 57312 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_15
timestamp 1621261055
transform -1 0 58848 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_17
timestamp 1621261055
transform -1 0 58848 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_589
timestamp 1621261055
transform 1 0 57696 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_595
timestamp 1621261055
transform 1 0 58272 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _143_
timestamp 1621261055
transform 1 0 2880 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_18
timestamp 1621261055
transform 1 0 1152 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_4
timestamp 1621261055
transform 1 0 1536 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_12
timestamp 1621261055
transform 1 0 2304 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_16
timestamp 1621261055
transform 1 0 2688 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_21
timestamp 1621261055
transform 1 0 3168 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_29
timestamp 1621261055
transform 1 0 3936 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_37
timestamp 1621261055
transform 1 0 4704 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_269
timestamp 1621261055
transform 1 0 6432 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_45
timestamp 1621261055
transform 1 0 5472 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_53
timestamp 1621261055
transform 1 0 6240 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_56
timestamp 1621261055
transform 1 0 6528 0 1 8658
box -38 -49 806 715
use BUFX2  BUFX2
timestamp 1624196784
transform 1 0 7680 0 1 8658
box 0 -48 864 714
use sky130_fd_sc_ls__diode_2  ANTENNA_41
timestamp 1621261055
transform 1 0 7488 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_64
timestamp 1621261055
transform 1 0 7296 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_77
timestamp 1621261055
transform 1 0 8544 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_85
timestamp 1621261055
transform 1 0 9312 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_93
timestamp 1621261055
transform 1 0 10080 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_101
timestamp 1621261055
transform 1 0 10848 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_270
timestamp 1621261055
transform 1 0 11712 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_9_109
timestamp 1621261055
transform 1 0 11616 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_111
timestamp 1621261055
transform 1 0 11808 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_119
timestamp 1621261055
transform 1 0 12576 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_127
timestamp 1621261055
transform 1 0 13344 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_135
timestamp 1621261055
transform 1 0 14112 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_143
timestamp 1621261055
transform 1 0 14880 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_271
timestamp 1621261055
transform 1 0 16992 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_151
timestamp 1621261055
transform 1 0 15648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_159
timestamp 1621261055
transform 1 0 16416 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_163
timestamp 1621261055
transform 1 0 16800 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_166
timestamp 1621261055
transform 1 0 17088 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_174
timestamp 1621261055
transform 1 0 17856 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_182
timestamp 1621261055
transform 1 0 18624 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_190
timestamp 1621261055
transform 1 0 19392 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_198
timestamp 1621261055
transform 1 0 20160 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_206
timestamp 1621261055
transform 1 0 20928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_272
timestamp 1621261055
transform 1 0 22272 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_214
timestamp 1621261055
transform 1 0 21696 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_218
timestamp 1621261055
transform 1 0 22080 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_221
timestamp 1621261055
transform 1 0 22368 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_229
timestamp 1621261055
transform 1 0 23136 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_237
timestamp 1621261055
transform 1 0 23904 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_245
timestamp 1621261055
transform 1 0 24672 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_253
timestamp 1621261055
transform 1 0 25440 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_261
timestamp 1621261055
transform 1 0 26208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_269
timestamp 1621261055
transform 1 0 26976 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_273
timestamp 1621261055
transform 1 0 27360 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_273
timestamp 1621261055
transform 1 0 27552 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_276
timestamp 1621261055
transform 1 0 27648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_284
timestamp 1621261055
transform 1 0 28416 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_292
timestamp 1621261055
transform 1 0 29184 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _007_
timestamp 1621261055
transform -1 0 30432 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_15
timestamp 1621261055
transform -1 0 30144 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_305
timestamp 1621261055
transform 1 0 30432 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_313
timestamp 1621261055
transform 1 0 31200 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_274
timestamp 1621261055
transform 1 0 32832 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_321
timestamp 1621261055
transform 1 0 31968 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_9_329
timestamp 1621261055
transform 1 0 32736 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_331
timestamp 1621261055
transform 1 0 32928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_339
timestamp 1621261055
transform 1 0 33696 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_347
timestamp 1621261055
transform 1 0 34464 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_355
timestamp 1621261055
transform 1 0 35232 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _016_
timestamp 1621261055
transform -1 0 36864 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _175_
timestamp 1621261055
transform 1 0 37248 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_29
timestamp 1621261055
transform -1 0 36576 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_9_363
timestamp 1621261055
transform 1 0 36000 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_9_372
timestamp 1621261055
transform 1 0 36864 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_275
timestamp 1621261055
transform 1 0 38112 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_379
timestamp 1621261055
transform 1 0 37536 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_383
timestamp 1621261055
transform 1 0 37920 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_386
timestamp 1621261055
transform 1 0 38208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_394
timestamp 1621261055
transform 1 0 38976 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_402
timestamp 1621261055
transform 1 0 39744 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_410
timestamp 1621261055
transform 1 0 40512 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_418
timestamp 1621261055
transform 1 0 41280 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_276
timestamp 1621261055
transform 1 0 43392 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_426
timestamp 1621261055
transform 1 0 42048 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_434
timestamp 1621261055
transform 1 0 42816 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_438
timestamp 1621261055
transform 1 0 43200 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_9_441
timestamp 1621261055
transform 1 0 43488 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _136_
timestamp 1621261055
transform 1 0 43872 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_9_448
timestamp 1621261055
transform 1 0 44160 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_456
timestamp 1621261055
transform 1 0 44928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_464
timestamp 1621261055
transform 1 0 45696 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_472
timestamp 1621261055
transform 1 0 46464 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_480
timestamp 1621261055
transform 1 0 47232 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _221_
timestamp 1621261055
transform 1 0 49152 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_277
timestamp 1621261055
transform 1 0 48672 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_488
timestamp 1621261055
transform 1 0 48000 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_492
timestamp 1621261055
transform 1 0 48384 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_494
timestamp 1621261055
transform 1 0 48576 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_496
timestamp 1621261055
transform 1 0 48768 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_503
timestamp 1621261055
transform 1 0 49440 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_511
timestamp 1621261055
transform 1 0 50208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_519
timestamp 1621261055
transform 1 0 50976 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output469
timestamp 1621261055
transform 1 0 53184 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_527
timestamp 1621261055
transform 1 0 51744 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_535
timestamp 1621261055
transform 1 0 52512 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_539
timestamp 1621261055
transform 1 0 52896 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_541
timestamp 1621261055
transform 1 0 53088 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_546
timestamp 1621261055
transform 1 0 53568 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_278
timestamp 1621261055
transform 1 0 53952 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output457
timestamp 1621261055
transform 1 0 54432 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output459
timestamp 1621261055
transform 1 0 55200 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_9_551
timestamp 1621261055
transform 1 0 54048 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_9_559
timestamp 1621261055
transform 1 0 54816 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_567
timestamp 1621261055
transform 1 0 55584 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input190
timestamp 1621261055
transform 1 0 57216 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input195
timestamp 1621261055
transform 1 0 56448 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_575
timestamp 1621261055
transform 1 0 56352 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_580
timestamp 1621261055
transform 1 0 56832 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_588
timestamp 1621261055
transform 1 0 57600 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_19
timestamp 1621261055
transform -1 0 58848 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_596
timestamp 1621261055
transform 1 0 58368 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_20
timestamp 1621261055
transform 1 0 1152 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_4
timestamp 1621261055
transform 1 0 1536 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_12
timestamp 1621261055
transform 1 0 2304 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_20
timestamp 1621261055
transform 1 0 3072 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_279
timestamp 1621261055
transform 1 0 3840 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_29
timestamp 1621261055
transform 1 0 3936 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_37
timestamp 1621261055
transform 1 0 4704 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_45
timestamp 1621261055
transform 1 0 5472 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_53
timestamp 1621261055
transform 1 0 6240 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_61
timestamp 1621261055
transform 1 0 7008 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_280
timestamp 1621261055
transform 1 0 9120 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_69
timestamp 1621261055
transform 1 0 7776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_77
timestamp 1621261055
transform 1 0 8544 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_81
timestamp 1621261055
transform 1 0 8928 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_84
timestamp 1621261055
transform 1 0 9216 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_92
timestamp 1621261055
transform 1 0 9984 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_100
timestamp 1621261055
transform 1 0 10752 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_108
timestamp 1621261055
transform 1 0 11520 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_116
timestamp 1621261055
transform 1 0 12288 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_124
timestamp 1621261055
transform 1 0 13056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_281
timestamp 1621261055
transform 1 0 14400 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_132
timestamp 1621261055
transform 1 0 13824 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_136
timestamp 1621261055
transform 1 0 14208 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_139
timestamp 1621261055
transform 1 0 14496 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_147
timestamp 1621261055
transform 1 0 15264 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_155
timestamp 1621261055
transform 1 0 16032 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_163
timestamp 1621261055
transform 1 0 16800 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_171
timestamp 1621261055
transform 1 0 17568 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_179
timestamp 1621261055
transform 1 0 18336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_187
timestamp 1621261055
transform 1 0 19104 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_282
timestamp 1621261055
transform 1 0 19680 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_191
timestamp 1621261055
transform 1 0 19488 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_194
timestamp 1621261055
transform 1 0 19776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_202
timestamp 1621261055
transform 1 0 20544 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_210
timestamp 1621261055
transform 1 0 21312 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_218
timestamp 1621261055
transform 1 0 22080 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_226
timestamp 1621261055
transform 1 0 22848 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_283
timestamp 1621261055
transform 1 0 24960 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_234
timestamp 1621261055
transform 1 0 23616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_242
timestamp 1621261055
transform 1 0 24384 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_246
timestamp 1621261055
transform 1 0 24768 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_249
timestamp 1621261055
transform 1 0 25056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_257
timestamp 1621261055
transform 1 0 25824 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_265
timestamp 1621261055
transform 1 0 26592 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_273
timestamp 1621261055
transform 1 0 27360 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_281
timestamp 1621261055
transform 1 0 28128 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_289
timestamp 1621261055
transform 1 0 28896 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_284
timestamp 1621261055
transform 1 0 30240 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_297
timestamp 1621261055
transform 1 0 29664 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_301
timestamp 1621261055
transform 1 0 30048 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_304
timestamp 1621261055
transform 1 0 30336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_312
timestamp 1621261055
transform 1 0 31104 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_320
timestamp 1621261055
transform 1 0 31872 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_328
timestamp 1621261055
transform 1 0 32640 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_336
timestamp 1621261055
transform 1 0 33408 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_344
timestamp 1621261055
transform 1 0 34176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_352
timestamp 1621261055
transform 1 0 34944 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_356
timestamp 1621261055
transform 1 0 35328 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_285
timestamp 1621261055
transform 1 0 35520 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_359
timestamp 1621261055
transform 1 0 35616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_367
timestamp 1621261055
transform 1 0 36384 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_375
timestamp 1621261055
transform 1 0 37152 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_383
timestamp 1621261055
transform 1 0 37920 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_391
timestamp 1621261055
transform 1 0 38688 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_399
timestamp 1621261055
transform 1 0 39456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_286
timestamp 1621261055
transform 1 0 40800 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_407
timestamp 1621261055
transform 1 0 40224 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_411
timestamp 1621261055
transform 1 0 40608 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_414
timestamp 1621261055
transform 1 0 40896 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_422
timestamp 1621261055
transform 1 0 41664 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_430
timestamp 1621261055
transform 1 0 42432 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_438
timestamp 1621261055
transform 1 0 43200 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_446
timestamp 1621261055
transform 1 0 43968 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_454
timestamp 1621261055
transform 1 0 44736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_462
timestamp 1621261055
transform 1 0 45504 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _054_
timestamp 1621261055
transform 1 0 46752 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_287
timestamp 1621261055
transform 1 0 46080 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_82
timestamp 1621261055
transform 1 0 46560 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_466
timestamp 1621261055
transform 1 0 45888 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_10_469
timestamp 1621261055
transform 1 0 46176 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_478
timestamp 1621261055
transform 1 0 47040 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_486
timestamp 1621261055
transform 1 0 47808 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_494
timestamp 1621261055
transform 1 0 48576 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_502
timestamp 1621261055
transform 1 0 49344 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_288
timestamp 1621261055
transform 1 0 51360 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_510
timestamp 1621261055
transform 1 0 50112 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_518
timestamp 1621261055
transform 1 0 50880 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_522
timestamp 1621261055
transform 1 0 51264 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_524
timestamp 1621261055
transform 1 0 51456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _077_
timestamp 1621261055
transform 1 0 53568 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _156_
timestamp 1621261055
transform 1 0 52896 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_10_532
timestamp 1621261055
transform 1 0 52224 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_536
timestamp 1621261055
transform 1 0 52608 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_538
timestamp 1621261055
transform 1 0 52800 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_542
timestamp 1621261055
transform 1 0 53184 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output458
timestamp 1621261055
transform 1 0 54240 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output460
timestamp 1621261055
transform -1 0 55392 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_113
timestamp 1621261055
transform -1 0 55008 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_10_549
timestamp 1621261055
transform 1 0 53856 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_557
timestamp 1621261055
transform 1 0 54624 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_10_565
timestamp 1621261055
transform 1 0 55392 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_289
timestamp 1621261055
transform 1 0 56640 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input191
timestamp 1621261055
transform 1 0 57600 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output461
timestamp 1621261055
transform 1 0 55776 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_573
timestamp 1621261055
transform 1 0 56160 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_577
timestamp 1621261055
transform 1 0 56544 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_579
timestamp 1621261055
transform 1 0 56736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_10_587
timestamp 1621261055
transform 1 0 57504 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_21
timestamp 1621261055
transform -1 0 58848 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_592
timestamp 1621261055
transform 1 0 57984 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_596
timestamp 1621261055
transform 1 0 58368 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_22
timestamp 1621261055
transform 1 0 1152 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_4
timestamp 1621261055
transform 1 0 1536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_12
timestamp 1621261055
transform 1 0 2304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_20
timestamp 1621261055
transform 1 0 3072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_28
timestamp 1621261055
transform 1 0 3840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_36
timestamp 1621261055
transform 1 0 4608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_290
timestamp 1621261055
transform 1 0 6432 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_44
timestamp 1621261055
transform 1 0 5376 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_52
timestamp 1621261055
transform 1 0 6144 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_54
timestamp 1621261055
transform 1 0 6336 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_56
timestamp 1621261055
transform 1 0 6528 0 1 9990
box -38 -49 806 715
use INV  INV
timestamp 1624196784
transform 1 0 7680 0 1 9990
box 0 -48 576 714
use sky130_fd_sc_ls__diode_2  ANTENNA_45
timestamp 1621261055
transform 1 0 7488 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_64
timestamp 1621261055
transform 1 0 7296 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_74
timestamp 1621261055
transform 1 0 8256 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_82
timestamp 1621261055
transform 1 0 9024 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_90
timestamp 1621261055
transform 1 0 9792 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_98
timestamp 1621261055
transform 1 0 10560 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_291
timestamp 1621261055
transform 1 0 11712 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_106
timestamp 1621261055
transform 1 0 11328 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_111
timestamp 1621261055
transform 1 0 11808 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_119
timestamp 1621261055
transform 1 0 12576 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_127
timestamp 1621261055
transform 1 0 13344 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_135
timestamp 1621261055
transform 1 0 14112 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_143
timestamp 1621261055
transform 1 0 14880 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_292
timestamp 1621261055
transform 1 0 16992 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_151
timestamp 1621261055
transform 1 0 15648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_159
timestamp 1621261055
transform 1 0 16416 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_163
timestamp 1621261055
transform 1 0 16800 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_166
timestamp 1621261055
transform 1 0 17088 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _193_
timestamp 1621261055
transform 1 0 17472 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_11_173
timestamp 1621261055
transform 1 0 17760 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_181
timestamp 1621261055
transform 1 0 18528 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_189
timestamp 1621261055
transform 1 0 19296 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_197
timestamp 1621261055
transform 1 0 20064 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_205
timestamp 1621261055
transform 1 0 20832 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_293
timestamp 1621261055
transform 1 0 22272 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_213
timestamp 1621261055
transform 1 0 21600 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_217
timestamp 1621261055
transform 1 0 21984 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_219
timestamp 1621261055
transform 1 0 22176 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_221
timestamp 1621261055
transform 1 0 22368 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_229
timestamp 1621261055
transform 1 0 23136 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_237
timestamp 1621261055
transform 1 0 23904 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_245
timestamp 1621261055
transform 1 0 24672 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_253
timestamp 1621261055
transform 1 0 25440 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_261
timestamp 1621261055
transform 1 0 26208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_269
timestamp 1621261055
transform 1 0 26976 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_273
timestamp 1621261055
transform 1 0 27360 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_294
timestamp 1621261055
transform 1 0 27552 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_276
timestamp 1621261055
transform 1 0 27648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_284
timestamp 1621261055
transform 1 0 28416 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_292
timestamp 1621261055
transform 1 0 29184 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_300
timestamp 1621261055
transform 1 0 29952 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_308
timestamp 1621261055
transform 1 0 30720 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_295
timestamp 1621261055
transform 1 0 32832 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_316
timestamp 1621261055
transform 1 0 31488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_324
timestamp 1621261055
transform 1 0 32256 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_328
timestamp 1621261055
transform 1 0 32640 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_331
timestamp 1621261055
transform 1 0 32928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_339
timestamp 1621261055
transform 1 0 33696 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_347
timestamp 1621261055
transform 1 0 34464 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_355
timestamp 1621261055
transform 1 0 35232 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_363
timestamp 1621261055
transform 1 0 36000 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_371
timestamp 1621261055
transform 1 0 36768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_296
timestamp 1621261055
transform 1 0 38112 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_379
timestamp 1621261055
transform 1 0 37536 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_383
timestamp 1621261055
transform 1 0 37920 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_386
timestamp 1621261055
transform 1 0 38208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_394
timestamp 1621261055
transform 1 0 38976 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_402
timestamp 1621261055
transform 1 0 39744 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_410
timestamp 1621261055
transform 1 0 40512 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_418
timestamp 1621261055
transform 1 0 41280 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_297
timestamp 1621261055
transform 1 0 43392 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_426
timestamp 1621261055
transform 1 0 42048 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_434
timestamp 1621261055
transform 1 0 42816 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_438
timestamp 1621261055
transform 1 0 43200 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_441
timestamp 1621261055
transform 1 0 43488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_449
timestamp 1621261055
transform 1 0 44256 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_457
timestamp 1621261055
transform 1 0 45024 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_465
timestamp 1621261055
transform 1 0 45792 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_473
timestamp 1621261055
transform 1 0 46560 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_481
timestamp 1621261055
transform 1 0 47328 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_298
timestamp 1621261055
transform 1 0 48672 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_489
timestamp 1621261055
transform 1 0 48096 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_493
timestamp 1621261055
transform 1 0 48480 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_496
timestamp 1621261055
transform 1 0 48768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_504
timestamp 1621261055
transform 1 0 49536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_512
timestamp 1621261055
transform 1 0 50304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_520
timestamp 1621261055
transform 1 0 51072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_528
timestamp 1621261055
transform 1 0 51840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_536
timestamp 1621261055
transform 1 0 52608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_544
timestamp 1621261055
transform 1 0 53376 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_299
timestamp 1621261055
transform 1 0 53952 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output471
timestamp 1621261055
transform -1 0 55296 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_115
timestamp 1621261055
transform -1 0 55680 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_126
timestamp 1621261055
transform -1 0 54912 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_548
timestamp 1621261055
transform 1 0 53760 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_551
timestamp 1621261055
transform 1 0 54048 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_555
timestamp 1621261055
transform 1 0 54432 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_557
timestamp 1621261055
transform 1 0 54624 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_564
timestamp 1621261055
transform 1 0 55296 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output462
timestamp 1621261055
transform -1 0 56064 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output463
timestamp 1621261055
transform 1 0 56448 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output464
timestamp 1621261055
transform -1 0 57600 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_116
timestamp 1621261055
transform -1 0 56256 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_117
timestamp 1621261055
transform -1 0 57216 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_574
timestamp 1621261055
transform 1 0 56256 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_580
timestamp 1621261055
transform 1 0 56832 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_588
timestamp 1621261055
transform 1 0 57600 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_23
timestamp 1621261055
transform -1 0 58848 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_596
timestamp 1621261055
transform 1 0 58368 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _029_
timestamp 1621261055
transform 1 0 2976 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_24
timestamp 1621261055
transform 1 0 1152 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_12
timestamp 1621261055
transform 1 0 2784 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_4
timestamp 1621261055
transform 1 0 1536 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_12
timestamp 1621261055
transform 1 0 2304 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_12_16
timestamp 1621261055
transform 1 0 2688 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_300
timestamp 1621261055
transform 1 0 3840 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_22
timestamp 1621261055
transform 1 0 3264 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_26
timestamp 1621261055
transform 1 0 3648 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_29
timestamp 1621261055
transform 1 0 3936 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_37
timestamp 1621261055
transform 1 0 4704 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_45
timestamp 1621261055
transform 1 0 5472 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_53
timestamp 1621261055
transform 1 0 6240 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_61
timestamp 1621261055
transform 1 0 7008 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_301
timestamp 1621261055
transform 1 0 9120 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_69
timestamp 1621261055
transform 1 0 7776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_77
timestamp 1621261055
transform 1 0 8544 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_81
timestamp 1621261055
transform 1 0 8928 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_84
timestamp 1621261055
transform 1 0 9216 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_92
timestamp 1621261055
transform 1 0 9984 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_100
timestamp 1621261055
transform 1 0 10752 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_108
timestamp 1621261055
transform 1 0 11520 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_116
timestamp 1621261055
transform 1 0 12288 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_124
timestamp 1621261055
transform 1 0 13056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_302
timestamp 1621261055
transform 1 0 14400 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_132
timestamp 1621261055
transform 1 0 13824 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_136
timestamp 1621261055
transform 1 0 14208 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_139
timestamp 1621261055
transform 1 0 14496 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_147
timestamp 1621261055
transform 1 0 15264 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_155
timestamp 1621261055
transform 1 0 16032 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_163
timestamp 1621261055
transform 1 0 16800 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_171
timestamp 1621261055
transform 1 0 17568 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_179
timestamp 1621261055
transform 1 0 18336 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_187
timestamp 1621261055
transform 1 0 19104 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_303
timestamp 1621261055
transform 1 0 19680 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_191
timestamp 1621261055
transform 1 0 19488 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_194
timestamp 1621261055
transform 1 0 19776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_202
timestamp 1621261055
transform 1 0 20544 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_210
timestamp 1621261055
transform 1 0 21312 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_218
timestamp 1621261055
transform 1 0 22080 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_226
timestamp 1621261055
transform 1 0 22848 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_304
timestamp 1621261055
transform 1 0 24960 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_234
timestamp 1621261055
transform 1 0 23616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_242
timestamp 1621261055
transform 1 0 24384 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_246
timestamp 1621261055
transform 1 0 24768 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_249
timestamp 1621261055
transform 1 0 25056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_257
timestamp 1621261055
transform 1 0 25824 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_265
timestamp 1621261055
transform 1 0 26592 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_273
timestamp 1621261055
transform 1 0 27360 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_281
timestamp 1621261055
transform 1 0 28128 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_289
timestamp 1621261055
transform 1 0 28896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_305
timestamp 1621261055
transform 1 0 30240 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_297
timestamp 1621261055
transform 1 0 29664 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_301
timestamp 1621261055
transform 1 0 30048 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_304
timestamp 1621261055
transform 1 0 30336 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_312
timestamp 1621261055
transform 1 0 31104 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_320
timestamp 1621261055
transform 1 0 31872 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_328
timestamp 1621261055
transform 1 0 32640 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_336
timestamp 1621261055
transform 1 0 33408 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_344
timestamp 1621261055
transform 1 0 34176 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_352
timestamp 1621261055
transform 1 0 34944 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_356
timestamp 1621261055
transform 1 0 35328 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_306
timestamp 1621261055
transform 1 0 35520 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_359
timestamp 1621261055
transform 1 0 35616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_367
timestamp 1621261055
transform 1 0 36384 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_375
timestamp 1621261055
transform 1 0 37152 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_383
timestamp 1621261055
transform 1 0 37920 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_391
timestamp 1621261055
transform 1 0 38688 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_399
timestamp 1621261055
transform 1 0 39456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_307
timestamp 1621261055
transform 1 0 40800 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_407
timestamp 1621261055
transform 1 0 40224 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_411
timestamp 1621261055
transform 1 0 40608 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_414
timestamp 1621261055
transform 1 0 40896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _157_
timestamp 1621261055
transform 1 0 41664 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_425
timestamp 1621261055
transform 1 0 41952 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_433
timestamp 1621261055
transform 1 0 42720 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_441
timestamp 1621261055
transform 1 0 43488 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _099_
timestamp 1621261055
transform 1 0 44544 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_449
timestamp 1621261055
transform 1 0 44256 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_451
timestamp 1621261055
transform 1 0 44448 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_455
timestamp 1621261055
transform 1 0 44832 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_308
timestamp 1621261055
transform 1 0 46080 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_463
timestamp 1621261055
transform 1 0 45600 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_12_467
timestamp 1621261055
transform 1 0 45984 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_469
timestamp 1621261055
transform 1 0 46176 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_477
timestamp 1621261055
transform 1 0 46944 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_485
timestamp 1621261055
transform 1 0 47712 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_493
timestamp 1621261055
transform 1 0 48480 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_501
timestamp 1621261055
transform 1 0 49248 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_309
timestamp 1621261055
transform 1 0 51360 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_509
timestamp 1621261055
transform 1 0 50016 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_517
timestamp 1621261055
transform 1 0 50784 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_521
timestamp 1621261055
transform 1 0 51168 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_524
timestamp 1621261055
transform 1 0 51456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_532
timestamp 1621261055
transform 1 0 52224 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_540
timestamp 1621261055
transform 1 0 52992 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _135_
timestamp 1621261055
transform 1 0 54528 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_548
timestamp 1621261055
transform 1 0 53760 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_559
timestamp 1621261055
transform 1 0 54816 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_567
timestamp 1621261055
transform 1 0 55584 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_310
timestamp 1621261055
transform 1 0 56640 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output465
timestamp 1621261055
transform 1 0 57120 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output470
timestamp 1621261055
transform 1 0 55872 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_119
timestamp 1621261055
transform 1 0 56928 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_569
timestamp 1621261055
transform 1 0 55776 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_574
timestamp 1621261055
transform 1 0 56256 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_579
timestamp 1621261055
transform 1 0 56736 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_587
timestamp 1621261055
transform 1 0 57504 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_25
timestamp 1621261055
transform -1 0 58848 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_595
timestamp 1621261055
transform 1 0 58272 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _051_
timestamp 1621261055
transform 1 0 2112 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _129_
timestamp 1621261055
transform 1 0 2784 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_26
timestamp 1621261055
transform 1 0 1152 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_70
timestamp 1621261055
transform 1 0 1920 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_13_4
timestamp 1621261055
transform 1 0 1536 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_13_13
timestamp 1621261055
transform 1 0 2400 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_20
timestamp 1621261055
transform 1 0 3072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_28
timestamp 1621261055
transform 1 0 3840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_36
timestamp 1621261055
transform 1 0 4608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_311
timestamp 1621261055
transform 1 0 6432 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_44
timestamp 1621261055
transform 1 0 5376 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_52
timestamp 1621261055
transform 1 0 6144 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_54
timestamp 1621261055
transform 1 0 6336 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_56
timestamp 1621261055
transform 1 0 6528 0 1 11322
box -38 -49 806 715
use INVX1  INVX1
timestamp 1624196784
transform 1 0 7680 0 1 11322
box 0 -48 576 714
use sky130_fd_sc_ls__diode_2  ANTENNA_49
timestamp 1621261055
transform 1 0 7488 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_64
timestamp 1621261055
transform 1 0 7296 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_74
timestamp 1621261055
transform 1 0 8256 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_82
timestamp 1621261055
transform 1 0 9024 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_90
timestamp 1621261055
transform 1 0 9792 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_98
timestamp 1621261055
transform 1 0 10560 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_312
timestamp 1621261055
transform 1 0 11712 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_106
timestamp 1621261055
transform 1 0 11328 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_111
timestamp 1621261055
transform 1 0 11808 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_119
timestamp 1621261055
transform 1 0 12576 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_127
timestamp 1621261055
transform 1 0 13344 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_135
timestamp 1621261055
transform 1 0 14112 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_143
timestamp 1621261055
transform 1 0 14880 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_313
timestamp 1621261055
transform 1 0 16992 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_151
timestamp 1621261055
transform 1 0 15648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_159
timestamp 1621261055
transform 1 0 16416 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_163
timestamp 1621261055
transform 1 0 16800 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_166
timestamp 1621261055
transform 1 0 17088 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_174
timestamp 1621261055
transform 1 0 17856 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_182
timestamp 1621261055
transform 1 0 18624 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_190
timestamp 1621261055
transform 1 0 19392 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_198
timestamp 1621261055
transform 1 0 20160 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_206
timestamp 1621261055
transform 1 0 20928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_314
timestamp 1621261055
transform 1 0 22272 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_214
timestamp 1621261055
transform 1 0 21696 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_218
timestamp 1621261055
transform 1 0 22080 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_221
timestamp 1621261055
transform 1 0 22368 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_229
timestamp 1621261055
transform 1 0 23136 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_237
timestamp 1621261055
transform 1 0 23904 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_245
timestamp 1621261055
transform 1 0 24672 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_253
timestamp 1621261055
transform 1 0 25440 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_261
timestamp 1621261055
transform 1 0 26208 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_269
timestamp 1621261055
transform 1 0 26976 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_273
timestamp 1621261055
transform 1 0 27360 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_315
timestamp 1621261055
transform 1 0 27552 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_276
timestamp 1621261055
transform 1 0 27648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_284
timestamp 1621261055
transform 1 0 28416 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_292
timestamp 1621261055
transform 1 0 29184 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_300
timestamp 1621261055
transform 1 0 29952 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_308
timestamp 1621261055
transform 1 0 30720 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_316
timestamp 1621261055
transform 1 0 32832 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_316
timestamp 1621261055
transform 1 0 31488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_324
timestamp 1621261055
transform 1 0 32256 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_328
timestamp 1621261055
transform 1 0 32640 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_331
timestamp 1621261055
transform 1 0 32928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _165_
timestamp 1621261055
transform 1 0 33696 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_13_342
timestamp 1621261055
transform 1 0 33984 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_350
timestamp 1621261055
transform 1 0 34752 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_358
timestamp 1621261055
transform 1 0 35520 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_366
timestamp 1621261055
transform 1 0 36288 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_374
timestamp 1621261055
transform 1 0 37056 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_317
timestamp 1621261055
transform 1 0 38112 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_382
timestamp 1621261055
transform 1 0 37824 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_384
timestamp 1621261055
transform 1 0 38016 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_386
timestamp 1621261055
transform 1 0 38208 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_394
timestamp 1621261055
transform 1 0 38976 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_398
timestamp 1621261055
transform 1 0 39360 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _053_
timestamp 1621261055
transform 1 0 39840 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_76
timestamp 1621261055
transform 1 0 39648 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_400
timestamp 1621261055
transform 1 0 39552 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_406
timestamp 1621261055
transform 1 0 40128 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_414
timestamp 1621261055
transform 1 0 40896 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_318
timestamp 1621261055
transform 1 0 43392 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_422
timestamp 1621261055
transform 1 0 41664 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_430
timestamp 1621261055
transform 1 0 42432 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_438
timestamp 1621261055
transform 1 0 43200 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_441
timestamp 1621261055
transform 1 0 43488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_449
timestamp 1621261055
transform 1 0 44256 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_457
timestamp 1621261055
transform 1 0 45024 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_465
timestamp 1621261055
transform 1 0 45792 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_473
timestamp 1621261055
transform 1 0 46560 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_481
timestamp 1621261055
transform 1 0 47328 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_319
timestamp 1621261055
transform 1 0 48672 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_489
timestamp 1621261055
transform 1 0 48096 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_493
timestamp 1621261055
transform 1 0 48480 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_496
timestamp 1621261055
transform 1 0 48768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_504
timestamp 1621261055
transform 1 0 49536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_512
timestamp 1621261055
transform 1 0 50304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_520
timestamp 1621261055
transform 1 0 51072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_528
timestamp 1621261055
transform 1 0 51840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_536
timestamp 1621261055
transform 1 0 52608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_544
timestamp 1621261055
transform 1 0 53376 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_320
timestamp 1621261055
transform 1 0 53952 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_10
timestamp 1621261055
transform 1 0 55488 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_548
timestamp 1621261055
transform 1 0 53760 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_551
timestamp 1621261055
transform 1 0 54048 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_559
timestamp 1621261055
transform 1 0 54816 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_563
timestamp 1621261055
transform 1 0 55200 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_565
timestamp 1621261055
transform 1 0 55392 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _018_
timestamp 1621261055
transform 1 0 55680 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output467
timestamp 1621261055
transform -1 0 57504 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output474
timestamp 1621261055
transform -1 0 56736 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_121
timestamp 1621261055
transform -1 0 57120 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_128
timestamp 1621261055
transform -1 0 56352 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_129
timestamp 1621261055
transform -1 0 56928 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_571
timestamp 1621261055
transform 1 0 55968 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_587
timestamp 1621261055
transform 1 0 57504 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_27
timestamp 1621261055
transform -1 0 58848 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_595
timestamp 1621261055
transform 1 0 58272 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_28
timestamp 1621261055
transform 1 0 1152 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_14_4
timestamp 1621261055
transform 1 0 1536 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_12
timestamp 1621261055
transform 1 0 2304 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_20
timestamp 1621261055
transform 1 0 3072 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_321
timestamp 1621261055
transform 1 0 3840 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_29
timestamp 1621261055
transform 1 0 3936 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_37
timestamp 1621261055
transform 1 0 4704 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_45
timestamp 1621261055
transform 1 0 5472 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_53
timestamp 1621261055
transform 1 0 6240 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_61
timestamp 1621261055
transform 1 0 7008 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_322
timestamp 1621261055
transform 1 0 9120 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_69
timestamp 1621261055
transform 1 0 7776 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_77
timestamp 1621261055
transform 1 0 8544 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_81
timestamp 1621261055
transform 1 0 8928 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_84
timestamp 1621261055
transform 1 0 9216 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_92
timestamp 1621261055
transform 1 0 9984 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_100
timestamp 1621261055
transform 1 0 10752 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_108
timestamp 1621261055
transform 1 0 11520 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_116
timestamp 1621261055
transform 1 0 12288 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_124
timestamp 1621261055
transform 1 0 13056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_323
timestamp 1621261055
transform 1 0 14400 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_132
timestamp 1621261055
transform 1 0 13824 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_136
timestamp 1621261055
transform 1 0 14208 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_139
timestamp 1621261055
transform 1 0 14496 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_147
timestamp 1621261055
transform 1 0 15264 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_155
timestamp 1621261055
transform 1 0 16032 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_163
timestamp 1621261055
transform 1 0 16800 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_171
timestamp 1621261055
transform 1 0 17568 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_179
timestamp 1621261055
transform 1 0 18336 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_187
timestamp 1621261055
transform 1 0 19104 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _158_
timestamp 1621261055
transform 1 0 20160 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_324
timestamp 1621261055
transform 1 0 19680 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_191
timestamp 1621261055
transform 1 0 19488 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_194
timestamp 1621261055
transform 1 0 19776 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_14_201
timestamp 1621261055
transform 1 0 20448 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_209
timestamp 1621261055
transform 1 0 21216 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_217
timestamp 1621261055
transform 1 0 21984 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_225
timestamp 1621261055
transform 1 0 22752 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_325
timestamp 1621261055
transform 1 0 24960 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_233
timestamp 1621261055
transform 1 0 23520 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_241
timestamp 1621261055
transform 1 0 24288 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_245
timestamp 1621261055
transform 1 0 24672 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_14_247
timestamp 1621261055
transform 1 0 24864 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_249
timestamp 1621261055
transform 1 0 25056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_257
timestamp 1621261055
transform 1 0 25824 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_265
timestamp 1621261055
transform 1 0 26592 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_273
timestamp 1621261055
transform 1 0 27360 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_281
timestamp 1621261055
transform 1 0 28128 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_289
timestamp 1621261055
transform 1 0 28896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _059_
timestamp 1621261055
transform 1 0 30816 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_326
timestamp 1621261055
transform 1 0 30240 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_297
timestamp 1621261055
transform 1 0 29664 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_301
timestamp 1621261055
transform 1 0 30048 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_304
timestamp 1621261055
transform 1 0 30336 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_14_308
timestamp 1621261055
transform 1 0 30720 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_312
timestamp 1621261055
transform 1 0 31104 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_320
timestamp 1621261055
transform 1 0 31872 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_328
timestamp 1621261055
transform 1 0 32640 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_336
timestamp 1621261055
transform 1 0 33408 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_344
timestamp 1621261055
transform 1 0 34176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_352
timestamp 1621261055
transform 1 0 34944 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_356
timestamp 1621261055
transform 1 0 35328 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_327
timestamp 1621261055
transform 1 0 35520 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_359
timestamp 1621261055
transform 1 0 35616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_367
timestamp 1621261055
transform 1 0 36384 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_375
timestamp 1621261055
transform 1 0 37152 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_383
timestamp 1621261055
transform 1 0 37920 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_391
timestamp 1621261055
transform 1 0 38688 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_399
timestamp 1621261055
transform 1 0 39456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_328
timestamp 1621261055
transform 1 0 40800 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_407
timestamp 1621261055
transform 1 0 40224 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_411
timestamp 1621261055
transform 1 0 40608 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_414
timestamp 1621261055
transform 1 0 40896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_422
timestamp 1621261055
transform 1 0 41664 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_430
timestamp 1621261055
transform 1 0 42432 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_438
timestamp 1621261055
transform 1 0 43200 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _132_
timestamp 1621261055
transform 1 0 44352 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_14_446
timestamp 1621261055
transform 1 0 43968 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_14_453
timestamp 1621261055
transform 1 0 44640 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_461
timestamp 1621261055
transform 1 0 45408 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_329
timestamp 1621261055
transform 1 0 46080 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_465
timestamp 1621261055
transform 1 0 45792 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_14_467
timestamp 1621261055
transform 1 0 45984 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_469
timestamp 1621261055
transform 1 0 46176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_477
timestamp 1621261055
transform 1 0 46944 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_485
timestamp 1621261055
transform 1 0 47712 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_493
timestamp 1621261055
transform 1 0 48480 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_501
timestamp 1621261055
transform 1 0 49248 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_330
timestamp 1621261055
transform 1 0 51360 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_509
timestamp 1621261055
transform 1 0 50016 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_517
timestamp 1621261055
transform 1 0 50784 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_521
timestamp 1621261055
transform 1 0 51168 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_524
timestamp 1621261055
transform 1 0 51456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_532
timestamp 1621261055
transform 1 0 52224 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_540
timestamp 1621261055
transform 1 0 52992 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_548
timestamp 1621261055
transform 1 0 53760 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_556
timestamp 1621261055
transform 1 0 54528 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_564
timestamp 1621261055
transform 1 0 55296 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_331
timestamp 1621261055
transform 1 0 56640 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output468
timestamp 1621261055
transform -1 0 57888 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_123
timestamp 1621261055
transform -1 0 57504 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_572
timestamp 1621261055
transform 1 0 56064 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_576
timestamp 1621261055
transform 1 0 56448 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_579
timestamp 1621261055
transform 1 0 56736 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_583
timestamp 1621261055
transform 1 0 57120 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_29
timestamp 1621261055
transform -1 0 58848 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_124
timestamp 1621261055
transform -1 0 58080 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_593
timestamp 1621261055
transform 1 0 58080 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_4
timestamp 1621261055
transform 1 0 1536 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_4
timestamp 1621261055
transform 1 0 1536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_32
timestamp 1621261055
transform 1 0 1152 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_30
timestamp 1621261055
transform 1 0 1152 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_16
timestamp 1621261055
transform 1 0 2688 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_12
timestamp 1621261055
transform 1 0 2304 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_12
timestamp 1621261055
transform 1 0 2304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_20
timestamp 1621261055
transform 1 0 3072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_53
timestamp 1621261055
transform 1 0 2880 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _045_
timestamp 1621261055
transform 1 0 3072 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_342
timestamp 1621261055
transform 1 0 3840 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_28
timestamp 1621261055
transform 1 0 3840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_36
timestamp 1621261055
transform 1 0 4608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_23
timestamp 1621261055
transform 1 0 3360 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_16_27
timestamp 1621261055
transform 1 0 3744 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_29
timestamp 1621261055
transform 1 0 3936 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_37
timestamp 1621261055
transform 1 0 4704 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _141_
timestamp 1621261055
transform 1 0 6624 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_332
timestamp 1621261055
transform 1 0 6432 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_44
timestamp 1621261055
transform 1 0 5376 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_52
timestamp 1621261055
transform 1 0 6144 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_15_54
timestamp 1621261055
transform 1 0 6336 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_56
timestamp 1621261055
transform 1 0 6528 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_45
timestamp 1621261055
transform 1 0 5472 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_53
timestamp 1621261055
transform 1 0 6240 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_16_60
timestamp 1621261055
transform 1 0 6912 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_70
timestamp 1621261055
transform 1 0 7872 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_16_64
timestamp 1621261055
transform 1 0 7296 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_64
timestamp 1621261055
transform 1 0 7296 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_92
timestamp 1621261055
transform 1 0 7392 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_51
timestamp 1621261055
transform 1 0 7488 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _058_
timestamp 1621261055
transform 1 0 7584 0 -1 13986
box -38 -49 326 715
use INVX2  INVX2
timestamp 1624196784
transform 1 0 7680 0 1 12654
box 0 -48 576 714
use sky130_fd_sc_ls__decap_4  FILLER_16_78
timestamp 1621261055
transform 1 0 8640 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_74
timestamp 1621261055
transform 1 0 8256 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_84
timestamp 1621261055
transform 1 0 9216 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_16_82
timestamp 1621261055
transform 1 0 9024 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_82
timestamp 1621261055
transform 1 0 9024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_343
timestamp 1621261055
transform 1 0 9120 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _176_
timestamp 1621261055
transform 1 0 11232 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_15_90
timestamp 1621261055
transform 1 0 9792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_98
timestamp 1621261055
transform 1 0 10560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_92
timestamp 1621261055
transform 1 0 9984 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_100
timestamp 1621261055
transform 1 0 10752 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_16_104
timestamp 1621261055
transform 1 0 11136 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_333
timestamp 1621261055
transform 1 0 11712 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_106
timestamp 1621261055
transform 1 0 11328 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_111
timestamp 1621261055
transform 1 0 11808 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_119
timestamp 1621261055
transform 1 0 12576 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_108
timestamp 1621261055
transform 1 0 11520 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_116
timestamp 1621261055
transform 1 0 12288 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_124
timestamp 1621261055
transform 1 0 13056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_344
timestamp 1621261055
transform 1 0 14400 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_127
timestamp 1621261055
transform 1 0 13344 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_135
timestamp 1621261055
transform 1 0 14112 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_143
timestamp 1621261055
transform 1 0 14880 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_132
timestamp 1621261055
transform 1 0 13824 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_136
timestamp 1621261055
transform 1 0 14208 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_139
timestamp 1621261055
transform 1 0 14496 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_147
timestamp 1621261055
transform 1 0 15264 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_334
timestamp 1621261055
transform 1 0 16992 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_151
timestamp 1621261055
transform 1 0 15648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_159
timestamp 1621261055
transform 1 0 16416 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_163
timestamp 1621261055
transform 1 0 16800 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_166
timestamp 1621261055
transform 1 0 17088 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_155
timestamp 1621261055
transform 1 0 16032 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_163
timestamp 1621261055
transform 1 0 16800 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_174
timestamp 1621261055
transform 1 0 17856 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_182
timestamp 1621261055
transform 1 0 18624 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_171
timestamp 1621261055
transform 1 0 17568 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_179
timestamp 1621261055
transform 1 0 18336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_187
timestamp 1621261055
transform 1 0 19104 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_345
timestamp 1621261055
transform 1 0 19680 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_190
timestamp 1621261055
transform 1 0 19392 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_198
timestamp 1621261055
transform 1 0 20160 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_206
timestamp 1621261055
transform 1 0 20928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_191
timestamp 1621261055
transform 1 0 19488 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_194
timestamp 1621261055
transform 1 0 19776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_202
timestamp 1621261055
transform 1 0 20544 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_210
timestamp 1621261055
transform 1 0 21312 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_335
timestamp 1621261055
transform 1 0 22272 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_214
timestamp 1621261055
transform 1 0 21696 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_218
timestamp 1621261055
transform 1 0 22080 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_221
timestamp 1621261055
transform 1 0 22368 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_229
timestamp 1621261055
transform 1 0 23136 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_218
timestamp 1621261055
transform 1 0 22080 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_226
timestamp 1621261055
transform 1 0 22848 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_346
timestamp 1621261055
transform 1 0 24960 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_237
timestamp 1621261055
transform 1 0 23904 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_245
timestamp 1621261055
transform 1 0 24672 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_234
timestamp 1621261055
transform 1 0 23616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_242
timestamp 1621261055
transform 1 0 24384 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_246
timestamp 1621261055
transform 1 0 24768 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_249
timestamp 1621261055
transform 1 0 25056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_253
timestamp 1621261055
transform 1 0 25440 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_261
timestamp 1621261055
transform 1 0 26208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_269
timestamp 1621261055
transform 1 0 26976 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_273
timestamp 1621261055
transform 1 0 27360 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_257
timestamp 1621261055
transform 1 0 25824 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_265
timestamp 1621261055
transform 1 0 26592 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_273
timestamp 1621261055
transform 1 0 27360 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _216_
timestamp 1621261055
transform 1 0 28800 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_336
timestamp 1621261055
transform 1 0 27552 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_276
timestamp 1621261055
transform 1 0 27648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_284
timestamp 1621261055
transform 1 0 28416 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_291
timestamp 1621261055
transform 1 0 29088 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_281
timestamp 1621261055
transform 1 0 28128 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_289
timestamp 1621261055
transform 1 0 28896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_347
timestamp 1621261055
transform 1 0 30240 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_299
timestamp 1621261055
transform 1 0 29856 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_307
timestamp 1621261055
transform 1 0 30624 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_315
timestamp 1621261055
transform 1 0 31392 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_297
timestamp 1621261055
transform 1 0 29664 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_301
timestamp 1621261055
transform 1 0 30048 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_304
timestamp 1621261055
transform 1 0 30336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_312
timestamp 1621261055
transform 1 0 31104 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_337
timestamp 1621261055
transform 1 0 32832 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_323
timestamp 1621261055
transform 1 0 32160 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_327
timestamp 1621261055
transform 1 0 32544 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_15_329
timestamp 1621261055
transform 1 0 32736 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_331
timestamp 1621261055
transform 1 0 32928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_320
timestamp 1621261055
transform 1 0 31872 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_328
timestamp 1621261055
transform 1 0 32640 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_336
timestamp 1621261055
transform 1 0 33408 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_339
timestamp 1621261055
transform 1 0 33696 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_347
timestamp 1621261055
transform 1 0 34464 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_355
timestamp 1621261055
transform 1 0 35232 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_344
timestamp 1621261055
transform 1 0 34176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_352
timestamp 1621261055
transform 1 0 34944 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_356
timestamp 1621261055
transform 1 0 35328 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_348
timestamp 1621261055
transform 1 0 35520 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_363
timestamp 1621261055
transform 1 0 36000 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_371
timestamp 1621261055
transform 1 0 36768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_359
timestamp 1621261055
transform 1 0 35616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_367
timestamp 1621261055
transform 1 0 36384 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_375
timestamp 1621261055
transform 1 0 37152 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_338
timestamp 1621261055
transform 1 0 38112 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_379
timestamp 1621261055
transform 1 0 37536 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_383
timestamp 1621261055
transform 1 0 37920 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_386
timestamp 1621261055
transform 1 0 38208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_394
timestamp 1621261055
transform 1 0 38976 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_383
timestamp 1621261055
transform 1 0 37920 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_391
timestamp 1621261055
transform 1 0 38688 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_399
timestamp 1621261055
transform 1 0 39456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_349
timestamp 1621261055
transform 1 0 40800 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_402
timestamp 1621261055
transform 1 0 39744 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_410
timestamp 1621261055
transform 1 0 40512 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_418
timestamp 1621261055
transform 1 0 41280 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_407
timestamp 1621261055
transform 1 0 40224 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_411
timestamp 1621261055
transform 1 0 40608 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_414
timestamp 1621261055
transform 1 0 40896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_339
timestamp 1621261055
transform 1 0 43392 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_426
timestamp 1621261055
transform 1 0 42048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_434
timestamp 1621261055
transform 1 0 42816 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_438
timestamp 1621261055
transform 1 0 43200 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_441
timestamp 1621261055
transform 1 0 43488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_422
timestamp 1621261055
transform 1 0 41664 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_430
timestamp 1621261055
transform 1 0 42432 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_438
timestamp 1621261055
transform 1 0 43200 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_449
timestamp 1621261055
transform 1 0 44256 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_457
timestamp 1621261055
transform 1 0 45024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_446
timestamp 1621261055
transform 1 0 43968 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_454
timestamp 1621261055
transform 1 0 44736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_462
timestamp 1621261055
transform 1 0 45504 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_350
timestamp 1621261055
transform 1 0 46080 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_465
timestamp 1621261055
transform 1 0 45792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_473
timestamp 1621261055
transform 1 0 46560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_481
timestamp 1621261055
transform 1 0 47328 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_466
timestamp 1621261055
transform 1 0 45888 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_469
timestamp 1621261055
transform 1 0 46176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_477
timestamp 1621261055
transform 1 0 46944 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_340
timestamp 1621261055
transform 1 0 48672 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_489
timestamp 1621261055
transform 1 0 48096 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_493
timestamp 1621261055
transform 1 0 48480 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_496
timestamp 1621261055
transform 1 0 48768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_504
timestamp 1621261055
transform 1 0 49536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_485
timestamp 1621261055
transform 1 0 47712 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_493
timestamp 1621261055
transform 1 0 48480 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_501
timestamp 1621261055
transform 1 0 49248 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_351
timestamp 1621261055
transform 1 0 51360 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_512
timestamp 1621261055
transform 1 0 50304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_520
timestamp 1621261055
transform 1 0 51072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_509
timestamp 1621261055
transform 1 0 50016 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_517
timestamp 1621261055
transform 1 0 50784 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_521
timestamp 1621261055
transform 1 0 51168 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_524
timestamp 1621261055
transform 1 0 51456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_528
timestamp 1621261055
transform 1 0 51840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_536
timestamp 1621261055
transform 1 0 52608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_544
timestamp 1621261055
transform 1 0 53376 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_532
timestamp 1621261055
transform 1 0 52224 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_540
timestamp 1621261055
transform 1 0 52992 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_341
timestamp 1621261055
transform 1 0 53952 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_548
timestamp 1621261055
transform 1 0 53760 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_551
timestamp 1621261055
transform 1 0 54048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_559
timestamp 1621261055
transform 1 0 54816 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_567
timestamp 1621261055
transform 1 0 55584 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_548
timestamp 1621261055
transform 1 0 53760 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_556
timestamp 1621261055
transform 1 0 54528 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_564
timestamp 1621261055
transform 1 0 55296 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_352
timestamp 1621261055
transform 1 0 56640 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_575
timestamp 1621261055
transform 1 0 56352 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_583
timestamp 1621261055
transform 1 0 57120 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_587
timestamp 1621261055
transform 1 0 57504 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_572
timestamp 1621261055
transform 1 0 56064 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_576
timestamp 1621261055
transform 1 0 56448 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_579
timestamp 1621261055
transform 1 0 56736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_587
timestamp 1621261055
transform 1 0 57504 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _067_
timestamp 1621261055
transform 1 0 57696 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_31
timestamp 1621261055
transform -1 0 58848 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_33
timestamp 1621261055
transform -1 0 58848 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_15_592
timestamp 1621261055
transform 1 0 57984 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_15_596
timestamp 1621261055
transform 1 0 58368 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_595
timestamp 1621261055
transform 1 0 58272 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_34
timestamp 1621261055
transform 1 0 1152 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_4
timestamp 1621261055
transform 1 0 1536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_12
timestamp 1621261055
transform 1 0 2304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_20
timestamp 1621261055
transform 1 0 3072 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_28
timestamp 1621261055
transform 1 0 3840 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_36
timestamp 1621261055
transform 1 0 4608 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_353
timestamp 1621261055
transform 1 0 6432 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_44
timestamp 1621261055
transform 1 0 5376 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_52
timestamp 1621261055
transform 1 0 6144 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_54
timestamp 1621261055
transform 1 0 6336 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_56
timestamp 1621261055
transform 1 0 6528 0 1 13986
box -38 -49 806 715
use INVX4  INVX4
timestamp 1624196784
transform 1 0 7680 0 1 13986
box 0 -48 864 714
use sky130_fd_sc_ls__diode_2  ANTENNA_55
timestamp 1621261055
transform 1 0 7488 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_64
timestamp 1621261055
transform 1 0 7296 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_77
timestamp 1621261055
transform 1 0 8544 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_85
timestamp 1621261055
transform 1 0 9312 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_93
timestamp 1621261055
transform 1 0 10080 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_101
timestamp 1621261055
transform 1 0 10848 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_354
timestamp 1621261055
transform 1 0 11712 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_17_109
timestamp 1621261055
transform 1 0 11616 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_111
timestamp 1621261055
transform 1 0 11808 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_119
timestamp 1621261055
transform 1 0 12576 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_127
timestamp 1621261055
transform 1 0 13344 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_135
timestamp 1621261055
transform 1 0 14112 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_143
timestamp 1621261055
transform 1 0 14880 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_355
timestamp 1621261055
transform 1 0 16992 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_151
timestamp 1621261055
transform 1 0 15648 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_159
timestamp 1621261055
transform 1 0 16416 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_163
timestamp 1621261055
transform 1 0 16800 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_166
timestamp 1621261055
transform 1 0 17088 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_174
timestamp 1621261055
transform 1 0 17856 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_182
timestamp 1621261055
transform 1 0 18624 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_190
timestamp 1621261055
transform 1 0 19392 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_198
timestamp 1621261055
transform 1 0 20160 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_206
timestamp 1621261055
transform 1 0 20928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_356
timestamp 1621261055
transform 1 0 22272 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_214
timestamp 1621261055
transform 1 0 21696 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_218
timestamp 1621261055
transform 1 0 22080 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_221
timestamp 1621261055
transform 1 0 22368 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_229
timestamp 1621261055
transform 1 0 23136 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_237
timestamp 1621261055
transform 1 0 23904 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_245
timestamp 1621261055
transform 1 0 24672 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_253
timestamp 1621261055
transform 1 0 25440 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_261
timestamp 1621261055
transform 1 0 26208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_269
timestamp 1621261055
transform 1 0 26976 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_273
timestamp 1621261055
transform 1 0 27360 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_357
timestamp 1621261055
transform 1 0 27552 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_276
timestamp 1621261055
transform 1 0 27648 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_284
timestamp 1621261055
transform 1 0 28416 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_292
timestamp 1621261055
transform 1 0 29184 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_300
timestamp 1621261055
transform 1 0 29952 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_308
timestamp 1621261055
transform 1 0 30720 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_358
timestamp 1621261055
transform 1 0 32832 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_316
timestamp 1621261055
transform 1 0 31488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_324
timestamp 1621261055
transform 1 0 32256 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_328
timestamp 1621261055
transform 1 0 32640 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_331
timestamp 1621261055
transform 1 0 32928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_339
timestamp 1621261055
transform 1 0 33696 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_347
timestamp 1621261055
transform 1 0 34464 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_355
timestamp 1621261055
transform 1 0 35232 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _037_
timestamp 1621261055
transform -1 0 37056 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_97
timestamp 1621261055
transform -1 0 36768 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_17_363
timestamp 1621261055
transform 1 0 36000 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_367
timestamp 1621261055
transform 1 0 36384 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_374
timestamp 1621261055
transform 1 0 37056 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_359
timestamp 1621261055
transform 1 0 38112 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_382
timestamp 1621261055
transform 1 0 37824 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_384
timestamp 1621261055
transform 1 0 38016 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_386
timestamp 1621261055
transform 1 0 38208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_394
timestamp 1621261055
transform 1 0 38976 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_402
timestamp 1621261055
transform 1 0 39744 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_410
timestamp 1621261055
transform 1 0 40512 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_418
timestamp 1621261055
transform 1 0 41280 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_360
timestamp 1621261055
transform 1 0 43392 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_426
timestamp 1621261055
transform 1 0 42048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_434
timestamp 1621261055
transform 1 0 42816 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_438
timestamp 1621261055
transform 1 0 43200 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_441
timestamp 1621261055
transform 1 0 43488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_449
timestamp 1621261055
transform 1 0 44256 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_457
timestamp 1621261055
transform 1 0 45024 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_465
timestamp 1621261055
transform 1 0 45792 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_473
timestamp 1621261055
transform 1 0 46560 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_481
timestamp 1621261055
transform 1 0 47328 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_361
timestamp 1621261055
transform 1 0 48672 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_489
timestamp 1621261055
transform 1 0 48096 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_493
timestamp 1621261055
transform 1 0 48480 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_496
timestamp 1621261055
transform 1 0 48768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_504
timestamp 1621261055
transform 1 0 49536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_512
timestamp 1621261055
transform 1 0 50304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_520
timestamp 1621261055
transform 1 0 51072 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_528
timestamp 1621261055
transform 1 0 51840 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_536
timestamp 1621261055
transform 1 0 52608 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_544
timestamp 1621261055
transform 1 0 53376 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_362
timestamp 1621261055
transform 1 0 53952 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_548
timestamp 1621261055
transform 1 0 53760 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_551
timestamp 1621261055
transform 1 0 54048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_559
timestamp 1621261055
transform 1 0 54816 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_567
timestamp 1621261055
transform 1 0 55584 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_575
timestamp 1621261055
transform 1 0 56352 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_583
timestamp 1621261055
transform 1 0 57120 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_35
timestamp 1621261055
transform -1 0 58848 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_17_591
timestamp 1621261055
transform 1 0 57888 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_595
timestamp 1621261055
transform 1 0 58272 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_36
timestamp 1621261055
transform 1 0 1152 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_18_4
timestamp 1621261055
transform 1 0 1536 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_12
timestamp 1621261055
transform 1 0 2304 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_20
timestamp 1621261055
transform 1 0 3072 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_363
timestamp 1621261055
transform 1 0 3840 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_29
timestamp 1621261055
transform 1 0 3936 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_37
timestamp 1621261055
transform 1 0 4704 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_45
timestamp 1621261055
transform 1 0 5472 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_53
timestamp 1621261055
transform 1 0 6240 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_61
timestamp 1621261055
transform 1 0 7008 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _192_
timestamp 1621261055
transform 1 0 7680 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_364
timestamp 1621261055
transform 1 0 9120 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_65
timestamp 1621261055
transform 1 0 7392 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_18_67
timestamp 1621261055
transform 1 0 7584 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_71
timestamp 1621261055
transform 1 0 7968 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_79
timestamp 1621261055
transform 1 0 8736 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_18_84
timestamp 1621261055
transform 1 0 9216 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_92
timestamp 1621261055
transform 1 0 9984 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_100
timestamp 1621261055
transform 1 0 10752 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_108
timestamp 1621261055
transform 1 0 11520 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_116
timestamp 1621261055
transform 1 0 12288 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_124
timestamp 1621261055
transform 1 0 13056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_365
timestamp 1621261055
transform 1 0 14400 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_132
timestamp 1621261055
transform 1 0 13824 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_136
timestamp 1621261055
transform 1 0 14208 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_139
timestamp 1621261055
transform 1 0 14496 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_147
timestamp 1621261055
transform 1 0 15264 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_155
timestamp 1621261055
transform 1 0 16032 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_163
timestamp 1621261055
transform 1 0 16800 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_171
timestamp 1621261055
transform 1 0 17568 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_179
timestamp 1621261055
transform 1 0 18336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_187
timestamp 1621261055
transform 1 0 19104 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _074_
timestamp 1621261055
transform 1 0 20256 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _078_
timestamp 1621261055
transform 1 0 20928 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_366
timestamp 1621261055
transform 1 0 19680 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_191
timestamp 1621261055
transform 1 0 19488 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_18_194
timestamp 1621261055
transform 1 0 19776 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_18_198
timestamp 1621261055
transform 1 0 20160 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_202
timestamp 1621261055
transform 1 0 20544 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_18_209
timestamp 1621261055
transform 1 0 21216 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_217
timestamp 1621261055
transform 1 0 21984 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_225
timestamp 1621261055
transform 1 0 22752 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_367
timestamp 1621261055
transform 1 0 24960 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_233
timestamp 1621261055
transform 1 0 23520 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_241
timestamp 1621261055
transform 1 0 24288 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_245
timestamp 1621261055
transform 1 0 24672 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_18_247
timestamp 1621261055
transform 1 0 24864 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_249
timestamp 1621261055
transform 1 0 25056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_257
timestamp 1621261055
transform 1 0 25824 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_265
timestamp 1621261055
transform 1 0 26592 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_273
timestamp 1621261055
transform 1 0 27360 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_281
timestamp 1621261055
transform 1 0 28128 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_289
timestamp 1621261055
transform 1 0 28896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_368
timestamp 1621261055
transform 1 0 30240 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_297
timestamp 1621261055
transform 1 0 29664 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_301
timestamp 1621261055
transform 1 0 30048 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_304
timestamp 1621261055
transform 1 0 30336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_312
timestamp 1621261055
transform 1 0 31104 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_320
timestamp 1621261055
transform 1 0 31872 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_328
timestamp 1621261055
transform 1 0 32640 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_336
timestamp 1621261055
transform 1 0 33408 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_344
timestamp 1621261055
transform 1 0 34176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_352
timestamp 1621261055
transform 1 0 34944 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_356
timestamp 1621261055
transform 1 0 35328 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _008_
timestamp 1621261055
transform -1 0 37056 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_369
timestamp 1621261055
transform 1 0 35520 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_17
timestamp 1621261055
transform -1 0 36768 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_359
timestamp 1621261055
transform 1 0 35616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_367
timestamp 1621261055
transform 1 0 36384 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_374
timestamp 1621261055
transform 1 0 37056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_382
timestamp 1621261055
transform 1 0 37824 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_390
timestamp 1621261055
transform 1 0 38592 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_398
timestamp 1621261055
transform 1 0 39360 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_370
timestamp 1621261055
transform 1 0 40800 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_406
timestamp 1621261055
transform 1 0 40128 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_410
timestamp 1621261055
transform 1 0 40512 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_18_412
timestamp 1621261055
transform 1 0 40704 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_414
timestamp 1621261055
transform 1 0 40896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_422
timestamp 1621261055
transform 1 0 41664 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_430
timestamp 1621261055
transform 1 0 42432 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_438
timestamp 1621261055
transform 1 0 43200 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_446
timestamp 1621261055
transform 1 0 43968 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_454
timestamp 1621261055
transform 1 0 44736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_462
timestamp 1621261055
transform 1 0 45504 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_371
timestamp 1621261055
transform 1 0 46080 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_466
timestamp 1621261055
transform 1 0 45888 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_469
timestamp 1621261055
transform 1 0 46176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_477
timestamp 1621261055
transform 1 0 46944 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_485
timestamp 1621261055
transform 1 0 47712 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_493
timestamp 1621261055
transform 1 0 48480 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_501
timestamp 1621261055
transform 1 0 49248 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_372
timestamp 1621261055
transform 1 0 51360 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_509
timestamp 1621261055
transform 1 0 50016 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_517
timestamp 1621261055
transform 1 0 50784 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_521
timestamp 1621261055
transform 1 0 51168 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_524
timestamp 1621261055
transform 1 0 51456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _170_
timestamp 1621261055
transform 1 0 52416 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_532
timestamp 1621261055
transform 1 0 52224 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_537
timestamp 1621261055
transform 1 0 52704 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_545
timestamp 1621261055
transform 1 0 53472 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_553
timestamp 1621261055
transform 1 0 54240 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_561
timestamp 1621261055
transform 1 0 55008 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_373
timestamp 1621261055
transform 1 0 56640 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_569
timestamp 1621261055
transform 1 0 55776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_18_577
timestamp 1621261055
transform 1 0 56544 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_579
timestamp 1621261055
transform 1 0 56736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_587
timestamp 1621261055
transform 1 0 57504 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_37
timestamp 1621261055
transform -1 0 58848 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_595
timestamp 1621261055
transform 1 0 58272 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_38
timestamp 1621261055
transform 1 0 1152 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_4
timestamp 1621261055
transform 1 0 1536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_12
timestamp 1621261055
transform 1 0 2304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_20
timestamp 1621261055
transform 1 0 3072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_28
timestamp 1621261055
transform 1 0 3840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_36
timestamp 1621261055
transform 1 0 4608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_374
timestamp 1621261055
transform 1 0 6432 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_44
timestamp 1621261055
transform 1 0 5376 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_52
timestamp 1621261055
transform 1 0 6144 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_54
timestamp 1621261055
transform 1 0 6336 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_56
timestamp 1621261055
transform 1 0 6528 0 1 15318
box -38 -49 806 715
use MUX2X1  MUX2X1
timestamp 1624196784
transform 1 0 7680 0 1 15318
box 0 -48 1728 714
use sky130_fd_sc_ls__diode_2  ANTENNA_63
timestamp 1621261055
transform 1 0 7488 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_64
timestamp 1621261055
transform 1 0 7296 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_86
timestamp 1621261055
transform 1 0 9408 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_94
timestamp 1621261055
transform 1 0 10176 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_102
timestamp 1621261055
transform 1 0 10944 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_375
timestamp 1621261055
transform 1 0 11712 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_111
timestamp 1621261055
transform 1 0 11808 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_119
timestamp 1621261055
transform 1 0 12576 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_127
timestamp 1621261055
transform 1 0 13344 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_135
timestamp 1621261055
transform 1 0 14112 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_143
timestamp 1621261055
transform 1 0 14880 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_376
timestamp 1621261055
transform 1 0 16992 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_151
timestamp 1621261055
transform 1 0 15648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_159
timestamp 1621261055
transform 1 0 16416 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_163
timestamp 1621261055
transform 1 0 16800 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_166
timestamp 1621261055
transform 1 0 17088 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_174
timestamp 1621261055
transform 1 0 17856 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_182
timestamp 1621261055
transform 1 0 18624 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_190
timestamp 1621261055
transform 1 0 19392 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_198
timestamp 1621261055
transform 1 0 20160 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_206
timestamp 1621261055
transform 1 0 20928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_377
timestamp 1621261055
transform 1 0 22272 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_214
timestamp 1621261055
transform 1 0 21696 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_218
timestamp 1621261055
transform 1 0 22080 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_221
timestamp 1621261055
transform 1 0 22368 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_229
timestamp 1621261055
transform 1 0 23136 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_237
timestamp 1621261055
transform 1 0 23904 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_245
timestamp 1621261055
transform 1 0 24672 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_253
timestamp 1621261055
transform 1 0 25440 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_261
timestamp 1621261055
transform 1 0 26208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_269
timestamp 1621261055
transform 1 0 26976 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_273
timestamp 1621261055
transform 1 0 27360 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_378
timestamp 1621261055
transform 1 0 27552 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_276
timestamp 1621261055
transform 1 0 27648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_284
timestamp 1621261055
transform 1 0 28416 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_292
timestamp 1621261055
transform 1 0 29184 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_300
timestamp 1621261055
transform 1 0 29952 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_308
timestamp 1621261055
transform 1 0 30720 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_379
timestamp 1621261055
transform 1 0 32832 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_316
timestamp 1621261055
transform 1 0 31488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_324
timestamp 1621261055
transform 1 0 32256 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_328
timestamp 1621261055
transform 1 0 32640 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_331
timestamp 1621261055
transform 1 0 32928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _027_
timestamp 1621261055
transform -1 0 35520 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_8
timestamp 1621261055
transform -1 0 35232 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_339
timestamp 1621261055
transform 1 0 33696 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_347
timestamp 1621261055
transform 1 0 34464 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_351
timestamp 1621261055
transform 1 0 34848 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_358
timestamp 1621261055
transform 1 0 35520 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_366
timestamp 1621261055
transform 1 0 36288 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_374
timestamp 1621261055
transform 1 0 37056 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_380
timestamp 1621261055
transform 1 0 38112 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_382
timestamp 1621261055
transform 1 0 37824 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_384
timestamp 1621261055
transform 1 0 38016 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_386
timestamp 1621261055
transform 1 0 38208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_394
timestamp 1621261055
transform 1 0 38976 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_402
timestamp 1621261055
transform 1 0 39744 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_410
timestamp 1621261055
transform 1 0 40512 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_418
timestamp 1621261055
transform 1 0 41280 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_381
timestamp 1621261055
transform 1 0 43392 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_426
timestamp 1621261055
transform 1 0 42048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_434
timestamp 1621261055
transform 1 0 42816 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_438
timestamp 1621261055
transform 1 0 43200 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_441
timestamp 1621261055
transform 1 0 43488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_449
timestamp 1621261055
transform 1 0 44256 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_457
timestamp 1621261055
transform 1 0 45024 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_465
timestamp 1621261055
transform 1 0 45792 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_473
timestamp 1621261055
transform 1 0 46560 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_481
timestamp 1621261055
transform 1 0 47328 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_382
timestamp 1621261055
transform 1 0 48672 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_489
timestamp 1621261055
transform 1 0 48096 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_493
timestamp 1621261055
transform 1 0 48480 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_496
timestamp 1621261055
transform 1 0 48768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_504
timestamp 1621261055
transform 1 0 49536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_512
timestamp 1621261055
transform 1 0 50304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_520
timestamp 1621261055
transform 1 0 51072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_528
timestamp 1621261055
transform 1 0 51840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_536
timestamp 1621261055
transform 1 0 52608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_544
timestamp 1621261055
transform 1 0 53376 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_383
timestamp 1621261055
transform 1 0 53952 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_548
timestamp 1621261055
transform 1 0 53760 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_551
timestamp 1621261055
transform 1 0 54048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_559
timestamp 1621261055
transform 1 0 54816 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_567
timestamp 1621261055
transform 1 0 55584 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_575
timestamp 1621261055
transform 1 0 56352 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_583
timestamp 1621261055
transform 1 0 57120 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_39
timestamp 1621261055
transform -1 0 58848 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_19_591
timestamp 1621261055
transform 1 0 57888 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_595
timestamp 1621261055
transform 1 0 58272 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_40
timestamp 1621261055
transform 1 0 1152 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_20_4
timestamp 1621261055
transform 1 0 1536 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_12
timestamp 1621261055
transform 1 0 2304 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_20
timestamp 1621261055
transform 1 0 3072 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_384
timestamp 1621261055
transform 1 0 3840 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_29
timestamp 1621261055
transform 1 0 3936 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_37
timestamp 1621261055
transform 1 0 4704 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_45
timestamp 1621261055
transform 1 0 5472 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_53
timestamp 1621261055
transform 1 0 6240 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_61
timestamp 1621261055
transform 1 0 7008 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_385
timestamp 1621261055
transform 1 0 9120 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_69
timestamp 1621261055
transform 1 0 7776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_77
timestamp 1621261055
transform 1 0 8544 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_81
timestamp 1621261055
transform 1 0 8928 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_84
timestamp 1621261055
transform 1 0 9216 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_92
timestamp 1621261055
transform 1 0 9984 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_100
timestamp 1621261055
transform 1 0 10752 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_108
timestamp 1621261055
transform 1 0 11520 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_116
timestamp 1621261055
transform 1 0 12288 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_124
timestamp 1621261055
transform 1 0 13056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_386
timestamp 1621261055
transform 1 0 14400 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_132
timestamp 1621261055
transform 1 0 13824 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_136
timestamp 1621261055
transform 1 0 14208 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_139
timestamp 1621261055
transform 1 0 14496 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_147
timestamp 1621261055
transform 1 0 15264 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_155
timestamp 1621261055
transform 1 0 16032 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_163
timestamp 1621261055
transform 1 0 16800 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_171
timestamp 1621261055
transform 1 0 17568 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_179
timestamp 1621261055
transform 1 0 18336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_187
timestamp 1621261055
transform 1 0 19104 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_387
timestamp 1621261055
transform 1 0 19680 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_191
timestamp 1621261055
transform 1 0 19488 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_194
timestamp 1621261055
transform 1 0 19776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_202
timestamp 1621261055
transform 1 0 20544 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_210
timestamp 1621261055
transform 1 0 21312 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_218
timestamp 1621261055
transform 1 0 22080 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_226
timestamp 1621261055
transform 1 0 22848 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_388
timestamp 1621261055
transform 1 0 24960 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_234
timestamp 1621261055
transform 1 0 23616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_242
timestamp 1621261055
transform 1 0 24384 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_246
timestamp 1621261055
transform 1 0 24768 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_249
timestamp 1621261055
transform 1 0 25056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_257
timestamp 1621261055
transform 1 0 25824 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_265
timestamp 1621261055
transform 1 0 26592 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_273
timestamp 1621261055
transform 1 0 27360 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_281
timestamp 1621261055
transform 1 0 28128 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_289
timestamp 1621261055
transform 1 0 28896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_389
timestamp 1621261055
transform 1 0 30240 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_297
timestamp 1621261055
transform 1 0 29664 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_301
timestamp 1621261055
transform 1 0 30048 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_304
timestamp 1621261055
transform 1 0 30336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_312
timestamp 1621261055
transform 1 0 31104 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_320
timestamp 1621261055
transform 1 0 31872 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_328
timestamp 1621261055
transform 1 0 32640 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_336
timestamp 1621261055
transform 1 0 33408 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_344
timestamp 1621261055
transform 1 0 34176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_352
timestamp 1621261055
transform 1 0 34944 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_356
timestamp 1621261055
transform 1 0 35328 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_390
timestamp 1621261055
transform 1 0 35520 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_359
timestamp 1621261055
transform 1 0 35616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_367
timestamp 1621261055
transform 1 0 36384 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_375
timestamp 1621261055
transform 1 0 37152 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_383
timestamp 1621261055
transform 1 0 37920 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_391
timestamp 1621261055
transform 1 0 38688 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_399
timestamp 1621261055
transform 1 0 39456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_391
timestamp 1621261055
transform 1 0 40800 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_407
timestamp 1621261055
transform 1 0 40224 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_411
timestamp 1621261055
transform 1 0 40608 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_414
timestamp 1621261055
transform 1 0 40896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_422
timestamp 1621261055
transform 1 0 41664 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_430
timestamp 1621261055
transform 1 0 42432 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_438
timestamp 1621261055
transform 1 0 43200 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _033_
timestamp 1621261055
transform 1 0 44256 0 -1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_27
timestamp 1621261055
transform 1 0 44064 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_20_446
timestamp 1621261055
transform 1 0 43968 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_452
timestamp 1621261055
transform 1 0 44544 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_460
timestamp 1621261055
transform 1 0 45312 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_392
timestamp 1621261055
transform 1 0 46080 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_469
timestamp 1621261055
transform 1 0 46176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_477
timestamp 1621261055
transform 1 0 46944 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _111_
timestamp 1621261055
transform 1 0 49344 0 -1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_20_485
timestamp 1621261055
transform 1 0 47712 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_493
timestamp 1621261055
transform 1 0 48480 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_20_501
timestamp 1621261055
transform 1 0 49248 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_393
timestamp 1621261055
transform 1 0 51360 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_505
timestamp 1621261055
transform 1 0 49632 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_513
timestamp 1621261055
transform 1 0 50400 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_521
timestamp 1621261055
transform 1 0 51168 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_524
timestamp 1621261055
transform 1 0 51456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_532
timestamp 1621261055
transform 1 0 52224 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_540
timestamp 1621261055
transform 1 0 52992 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_548
timestamp 1621261055
transform 1 0 53760 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_556
timestamp 1621261055
transform 1 0 54528 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_564
timestamp 1621261055
transform 1 0 55296 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_394
timestamp 1621261055
transform 1 0 56640 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_572
timestamp 1621261055
transform 1 0 56064 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_576
timestamp 1621261055
transform 1 0 56448 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_579
timestamp 1621261055
transform 1 0 56736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_587
timestamp 1621261055
transform 1 0 57504 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_41
timestamp 1621261055
transform -1 0 58848 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_595
timestamp 1621261055
transform 1 0 58272 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_42
timestamp 1621261055
transform 1 0 1152 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_21_4
timestamp 1621261055
transform 1 0 1536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_12
timestamp 1621261055
transform 1 0 2304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_20
timestamp 1621261055
transform 1 0 3072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_28
timestamp 1621261055
transform 1 0 3840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_36
timestamp 1621261055
transform 1 0 4608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_395
timestamp 1621261055
transform 1 0 6432 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_44
timestamp 1621261055
transform 1 0 5376 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_52
timestamp 1621261055
transform 1 0 6144 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_21_54
timestamp 1621261055
transform 1 0 6336 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_56
timestamp 1621261055
transform 1 0 6528 0 1 16650
box -38 -49 806 715
use NAND2X1  NAND2X1
timestamp 1624196784
transform 1 0 7680 0 1 16650
box 0 -48 864 714
use sky130_fd_sc_ls__diode_2  ANTENNA_68
timestamp 1621261055
transform 1 0 7488 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_64
timestamp 1621261055
transform 1 0 7296 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_77
timestamp 1621261055
transform 1 0 8544 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_85
timestamp 1621261055
transform 1 0 9312 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_93
timestamp 1621261055
transform 1 0 10080 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_101
timestamp 1621261055
transform 1 0 10848 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_396
timestamp 1621261055
transform 1 0 11712 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_21_109
timestamp 1621261055
transform 1 0 11616 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_111
timestamp 1621261055
transform 1 0 11808 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_119
timestamp 1621261055
transform 1 0 12576 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_127
timestamp 1621261055
transform 1 0 13344 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_135
timestamp 1621261055
transform 1 0 14112 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_143
timestamp 1621261055
transform 1 0 14880 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_397
timestamp 1621261055
transform 1 0 16992 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_151
timestamp 1621261055
transform 1 0 15648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_159
timestamp 1621261055
transform 1 0 16416 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_163
timestamp 1621261055
transform 1 0 16800 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_166
timestamp 1621261055
transform 1 0 17088 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _116_
timestamp 1621261055
transform 1 0 19200 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_21_174
timestamp 1621261055
transform 1 0 17856 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_182
timestamp 1621261055
transform 1 0 18624 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_186
timestamp 1621261055
transform 1 0 19008 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_191
timestamp 1621261055
transform 1 0 19488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_199
timestamp 1621261055
transform 1 0 20256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_207
timestamp 1621261055
transform 1 0 21024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_398
timestamp 1621261055
transform 1 0 22272 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_215
timestamp 1621261055
transform 1 0 21792 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_21_219
timestamp 1621261055
transform 1 0 22176 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_221
timestamp 1621261055
transform 1 0 22368 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_229
timestamp 1621261055
transform 1 0 23136 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_237
timestamp 1621261055
transform 1 0 23904 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_245
timestamp 1621261055
transform 1 0 24672 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_253
timestamp 1621261055
transform 1 0 25440 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_261
timestamp 1621261055
transform 1 0 26208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_269
timestamp 1621261055
transform 1 0 26976 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_273
timestamp 1621261055
transform 1 0 27360 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_399
timestamp 1621261055
transform 1 0 27552 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_276
timestamp 1621261055
transform 1 0 27648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_284
timestamp 1621261055
transform 1 0 28416 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_292
timestamp 1621261055
transform 1 0 29184 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_300
timestamp 1621261055
transform 1 0 29952 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_308
timestamp 1621261055
transform 1 0 30720 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_400
timestamp 1621261055
transform 1 0 32832 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_316
timestamp 1621261055
transform 1 0 31488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_324
timestamp 1621261055
transform 1 0 32256 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_328
timestamp 1621261055
transform 1 0 32640 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_331
timestamp 1621261055
transform 1 0 32928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_101
timestamp 1621261055
transform -1 0 35520 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_339
timestamp 1621261055
transform 1 0 33696 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_347
timestamp 1621261055
transform 1 0 34464 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_21_355
timestamp 1621261055
transform 1 0 35232 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _038_
timestamp 1621261055
transform -1 0 35808 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_21_361
timestamp 1621261055
transform 1 0 35808 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_369
timestamp 1621261055
transform 1 0 36576 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_377
timestamp 1621261055
transform 1 0 37344 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_401
timestamp 1621261055
transform 1 0 38112 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_386
timestamp 1621261055
transform 1 0 38208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_394
timestamp 1621261055
transform 1 0 38976 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_402
timestamp 1621261055
transform 1 0 39744 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_410
timestamp 1621261055
transform 1 0 40512 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_418
timestamp 1621261055
transform 1 0 41280 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_402
timestamp 1621261055
transform 1 0 43392 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_426
timestamp 1621261055
transform 1 0 42048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_434
timestamp 1621261055
transform 1 0 42816 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_438
timestamp 1621261055
transform 1 0 43200 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_441
timestamp 1621261055
transform 1 0 43488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_449
timestamp 1621261055
transform 1 0 44256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_457
timestamp 1621261055
transform 1 0 45024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_465
timestamp 1621261055
transform 1 0 45792 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_473
timestamp 1621261055
transform 1 0 46560 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_481
timestamp 1621261055
transform 1 0 47328 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_403
timestamp 1621261055
transform 1 0 48672 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_489
timestamp 1621261055
transform 1 0 48096 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_493
timestamp 1621261055
transform 1 0 48480 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_496
timestamp 1621261055
transform 1 0 48768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_504
timestamp 1621261055
transform 1 0 49536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_512
timestamp 1621261055
transform 1 0 50304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_520
timestamp 1621261055
transform 1 0 51072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_528
timestamp 1621261055
transform 1 0 51840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_536
timestamp 1621261055
transform 1 0 52608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_544
timestamp 1621261055
transform 1 0 53376 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_404
timestamp 1621261055
transform 1 0 53952 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_548
timestamp 1621261055
transform 1 0 53760 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_551
timestamp 1621261055
transform 1 0 54048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_559
timestamp 1621261055
transform 1 0 54816 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_567
timestamp 1621261055
transform 1 0 55584 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_575
timestamp 1621261055
transform 1 0 56352 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_583
timestamp 1621261055
transform 1 0 57120 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_43
timestamp 1621261055
transform -1 0 58848 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_21_591
timestamp 1621261055
transform 1 0 57888 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_595
timestamp 1621261055
transform 1 0 58272 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_44
timestamp 1621261055
transform 1 0 1152 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_22_4
timestamp 1621261055
transform 1 0 1536 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_12
timestamp 1621261055
transform 1 0 2304 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_20
timestamp 1621261055
transform 1 0 3072 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_405
timestamp 1621261055
transform 1 0 3840 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_29
timestamp 1621261055
transform 1 0 3936 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_37
timestamp 1621261055
transform 1 0 4704 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_45
timestamp 1621261055
transform 1 0 5472 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_53
timestamp 1621261055
transform 1 0 6240 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_61
timestamp 1621261055
transform 1 0 7008 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_406
timestamp 1621261055
transform 1 0 9120 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_69
timestamp 1621261055
transform 1 0 7776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_77
timestamp 1621261055
transform 1 0 8544 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_81
timestamp 1621261055
transform 1 0 8928 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_84
timestamp 1621261055
transform 1 0 9216 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_92
timestamp 1621261055
transform 1 0 9984 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_100
timestamp 1621261055
transform 1 0 10752 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_108
timestamp 1621261055
transform 1 0 11520 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_116
timestamp 1621261055
transform 1 0 12288 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_124
timestamp 1621261055
transform 1 0 13056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_407
timestamp 1621261055
transform 1 0 14400 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_132
timestamp 1621261055
transform 1 0 13824 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_136
timestamp 1621261055
transform 1 0 14208 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_139
timestamp 1621261055
transform 1 0 14496 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_147
timestamp 1621261055
transform 1 0 15264 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_155
timestamp 1621261055
transform 1 0 16032 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_163
timestamp 1621261055
transform 1 0 16800 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_171
timestamp 1621261055
transform 1 0 17568 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_179
timestamp 1621261055
transform 1 0 18336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_187
timestamp 1621261055
transform 1 0 19104 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_408
timestamp 1621261055
transform 1 0 19680 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_191
timestamp 1621261055
transform 1 0 19488 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_194
timestamp 1621261055
transform 1 0 19776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_202
timestamp 1621261055
transform 1 0 20544 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_210
timestamp 1621261055
transform 1 0 21312 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _019_
timestamp 1621261055
transform 1 0 22464 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _213_
timestamp 1621261055
transform 1 0 23136 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_31
timestamp 1621261055
transform 1 0 22272 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_218
timestamp 1621261055
transform 1 0 22080 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_22_225
timestamp 1621261055
transform 1 0 22752 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_409
timestamp 1621261055
transform 1 0 24960 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_232
timestamp 1621261055
transform 1 0 23424 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_240
timestamp 1621261055
transform 1 0 24192 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_249
timestamp 1621261055
transform 1 0 25056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_257
timestamp 1621261055
transform 1 0 25824 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_265
timestamp 1621261055
transform 1 0 26592 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_273
timestamp 1621261055
transform 1 0 27360 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_281
timestamp 1621261055
transform 1 0 28128 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_289
timestamp 1621261055
transform 1 0 28896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_410
timestamp 1621261055
transform 1 0 30240 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_297
timestamp 1621261055
transform 1 0 29664 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_301
timestamp 1621261055
transform 1 0 30048 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_304
timestamp 1621261055
transform 1 0 30336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_312
timestamp 1621261055
transform 1 0 31104 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_320
timestamp 1621261055
transform 1 0 31872 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_328
timestamp 1621261055
transform 1 0 32640 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_336
timestamp 1621261055
transform 1 0 33408 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_344
timestamp 1621261055
transform 1 0 34176 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_352
timestamp 1621261055
transform 1 0 34944 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_356
timestamp 1621261055
transform 1 0 35328 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_411
timestamp 1621261055
transform 1 0 35520 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_359
timestamp 1621261055
transform 1 0 35616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_367
timestamp 1621261055
transform 1 0 36384 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_375
timestamp 1621261055
transform 1 0 37152 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_383
timestamp 1621261055
transform 1 0 37920 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_391
timestamp 1621261055
transform 1 0 38688 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_399
timestamp 1621261055
transform 1 0 39456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_412
timestamp 1621261055
transform 1 0 40800 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_407
timestamp 1621261055
transform 1 0 40224 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_411
timestamp 1621261055
transform 1 0 40608 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_414
timestamp 1621261055
transform 1 0 40896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_422
timestamp 1621261055
transform 1 0 41664 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_430
timestamp 1621261055
transform 1 0 42432 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_438
timestamp 1621261055
transform 1 0 43200 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_446
timestamp 1621261055
transform 1 0 43968 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_454
timestamp 1621261055
transform 1 0 44736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_462
timestamp 1621261055
transform 1 0 45504 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_413
timestamp 1621261055
transform 1 0 46080 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_466
timestamp 1621261055
transform 1 0 45888 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_469
timestamp 1621261055
transform 1 0 46176 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_477
timestamp 1621261055
transform 1 0 46944 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_485
timestamp 1621261055
transform 1 0 47712 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_493
timestamp 1621261055
transform 1 0 48480 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_501
timestamp 1621261055
transform 1 0 49248 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_414
timestamp 1621261055
transform 1 0 51360 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_509
timestamp 1621261055
transform 1 0 50016 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_517
timestamp 1621261055
transform 1 0 50784 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_521
timestamp 1621261055
transform 1 0 51168 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_524
timestamp 1621261055
transform 1 0 51456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_532
timestamp 1621261055
transform 1 0 52224 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_540
timestamp 1621261055
transform 1 0 52992 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_548
timestamp 1621261055
transform 1 0 53760 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_556
timestamp 1621261055
transform 1 0 54528 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_564
timestamp 1621261055
transform 1 0 55296 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_415
timestamp 1621261055
transform 1 0 56640 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_572
timestamp 1621261055
transform 1 0 56064 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_576
timestamp 1621261055
transform 1 0 56448 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_579
timestamp 1621261055
transform 1 0 56736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_587
timestamp 1621261055
transform 1 0 57504 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_45
timestamp 1621261055
transform -1 0 58848 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_595
timestamp 1621261055
transform 1 0 58272 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_46
timestamp 1621261055
transform 1 0 1152 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_48
timestamp 1621261055
transform 1 0 1152 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_4
timestamp 1621261055
transform 1 0 1536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_12
timestamp 1621261055
transform 1 0 2304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_20
timestamp 1621261055
transform 1 0 3072 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_4
timestamp 1621261055
transform 1 0 1536 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_12
timestamp 1621261055
transform 1 0 2304 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_20
timestamp 1621261055
transform 1 0 3072 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_426
timestamp 1621261055
transform 1 0 3840 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_28
timestamp 1621261055
transform 1 0 3840 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_36
timestamp 1621261055
transform 1 0 4608 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_29
timestamp 1621261055
transform 1 0 3936 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_37
timestamp 1621261055
transform 1 0 4704 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_416
timestamp 1621261055
transform 1 0 6432 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_44
timestamp 1621261055
transform 1 0 5376 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_52
timestamp 1621261055
transform 1 0 6144 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_23_54
timestamp 1621261055
transform 1 0 6336 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_56
timestamp 1621261055
transform 1 0 6528 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_45
timestamp 1621261055
transform 1 0 5472 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_53
timestamp 1621261055
transform 1 0 6240 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_61
timestamp 1621261055
transform 1 0 7008 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_69
timestamp 1621261055
transform 1 0 7776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_24_65
timestamp 1621261055
transform 1 0 7392 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_64
timestamp 1621261055
transform 1 0 7296 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_80
timestamp 1621261055
transform 1 0 7488 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _113_
timestamp 1621261055
transform 1 0 7488 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_84
timestamp 1621261055
transform 1 0 9216 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_81
timestamp 1621261055
transform 1 0 8928 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_77
timestamp 1621261055
transform 1 0 8544 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_80
timestamp 1621261055
transform 1 0 8832 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_427
timestamp 1621261055
transform 1 0 9120 0 -1 19314
box -38 -49 134 715
use NAND3X1  NAND3X1
timestamp 1624196784
transform 1 0 7680 0 1 17982
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_8  FILLER_23_88
timestamp 1621261055
transform 1 0 9600 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_96
timestamp 1621261055
transform 1 0 10368 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_104
timestamp 1621261055
transform 1 0 11136 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_92
timestamp 1621261055
transform 1 0 9984 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_100
timestamp 1621261055
transform 1 0 10752 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_417
timestamp 1621261055
transform 1 0 11712 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_108
timestamp 1621261055
transform 1 0 11520 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_111
timestamp 1621261055
transform 1 0 11808 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_119
timestamp 1621261055
transform 1 0 12576 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_108
timestamp 1621261055
transform 1 0 11520 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_116
timestamp 1621261055
transform 1 0 12288 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_124
timestamp 1621261055
transform 1 0 13056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_428
timestamp 1621261055
transform 1 0 14400 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_127
timestamp 1621261055
transform 1 0 13344 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_135
timestamp 1621261055
transform 1 0 14112 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_143
timestamp 1621261055
transform 1 0 14880 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_132
timestamp 1621261055
transform 1 0 13824 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_136
timestamp 1621261055
transform 1 0 14208 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_139
timestamp 1621261055
transform 1 0 14496 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_147
timestamp 1621261055
transform 1 0 15264 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_418
timestamp 1621261055
transform 1 0 16992 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_151
timestamp 1621261055
transform 1 0 15648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_159
timestamp 1621261055
transform 1 0 16416 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_163
timestamp 1621261055
transform 1 0 16800 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_166
timestamp 1621261055
transform 1 0 17088 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_155
timestamp 1621261055
transform 1 0 16032 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_163
timestamp 1621261055
transform 1 0 16800 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _069_
timestamp 1621261055
transform 1 0 18048 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_174
timestamp 1621261055
transform 1 0 17856 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_179
timestamp 1621261055
transform 1 0 18336 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_187
timestamp 1621261055
transform 1 0 19104 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_171
timestamp 1621261055
transform 1 0 17568 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_179
timestamp 1621261055
transform 1 0 18336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_187
timestamp 1621261055
transform 1 0 19104 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_429
timestamp 1621261055
transform 1 0 19680 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_195
timestamp 1621261055
transform 1 0 19872 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_203
timestamp 1621261055
transform 1 0 20640 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_191
timestamp 1621261055
transform 1 0 19488 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_194
timestamp 1621261055
transform 1 0 19776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_202
timestamp 1621261055
transform 1 0 20544 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_210
timestamp 1621261055
transform 1 0 21312 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_419
timestamp 1621261055
transform 1 0 22272 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_211
timestamp 1621261055
transform 1 0 21408 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_219
timestamp 1621261055
transform 1 0 22176 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_221
timestamp 1621261055
transform 1 0 22368 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_229
timestamp 1621261055
transform 1 0 23136 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_218
timestamp 1621261055
transform 1 0 22080 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_226
timestamp 1621261055
transform 1 0 22848 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_430
timestamp 1621261055
transform 1 0 24960 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_237
timestamp 1621261055
transform 1 0 23904 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_245
timestamp 1621261055
transform 1 0 24672 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_234
timestamp 1621261055
transform 1 0 23616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_242
timestamp 1621261055
transform 1 0 24384 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_246
timestamp 1621261055
transform 1 0 24768 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_249
timestamp 1621261055
transform 1 0 25056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_253
timestamp 1621261055
transform 1 0 25440 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_261
timestamp 1621261055
transform 1 0 26208 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_269
timestamp 1621261055
transform 1 0 26976 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_273
timestamp 1621261055
transform 1 0 27360 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_257
timestamp 1621261055
transform 1 0 25824 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_265
timestamp 1621261055
transform 1 0 26592 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_273
timestamp 1621261055
transform 1 0 27360 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_420
timestamp 1621261055
transform 1 0 27552 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_276
timestamp 1621261055
transform 1 0 27648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_284
timestamp 1621261055
transform 1 0 28416 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_292
timestamp 1621261055
transform 1 0 29184 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_281
timestamp 1621261055
transform 1 0 28128 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_289
timestamp 1621261055
transform 1 0 28896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_301
timestamp 1621261055
transform 1 0 30048 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_297
timestamp 1621261055
transform 1 0 29664 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_23_300
timestamp 1621261055
transform 1 0 29952 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_304
timestamp 1621261055
transform 1 0 30336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_310
timestamp 1621261055
transform 1 0 30912 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_306
timestamp 1621261055
transform 1 0 30528 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_304
timestamp 1621261055
transform 1 0 30336 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_431
timestamp 1621261055
transform 1 0 30240 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _133_
timestamp 1621261055
transform 1 0 30624 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_312
timestamp 1621261055
transform 1 0 31104 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_421
timestamp 1621261055
transform 1 0 32832 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_318
timestamp 1621261055
transform 1 0 31680 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_326
timestamp 1621261055
transform 1 0 32448 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_331
timestamp 1621261055
transform 1 0 32928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_320
timestamp 1621261055
transform 1 0 31872 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_328
timestamp 1621261055
transform 1 0 32640 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_336
timestamp 1621261055
transform 1 0 33408 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_339
timestamp 1621261055
transform 1 0 33696 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_347
timestamp 1621261055
transform 1 0 34464 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_355
timestamp 1621261055
transform 1 0 35232 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_344
timestamp 1621261055
transform 1 0 34176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_352
timestamp 1621261055
transform 1 0 34944 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_356
timestamp 1621261055
transform 1 0 35328 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_432
timestamp 1621261055
transform 1 0 35520 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_363
timestamp 1621261055
transform 1 0 36000 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_371
timestamp 1621261055
transform 1 0 36768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_359
timestamp 1621261055
transform 1 0 35616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_367
timestamp 1621261055
transform 1 0 36384 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_375
timestamp 1621261055
transform 1 0 37152 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_422
timestamp 1621261055
transform 1 0 38112 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_23_379
timestamp 1621261055
transform 1 0 37536 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_383
timestamp 1621261055
transform 1 0 37920 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_386
timestamp 1621261055
transform 1 0 38208 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_394
timestamp 1621261055
transform 1 0 38976 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_383
timestamp 1621261055
transform 1 0 37920 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_391
timestamp 1621261055
transform 1 0 38688 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_399
timestamp 1621261055
transform 1 0 39456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_433
timestamp 1621261055
transform 1 0 40800 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_402
timestamp 1621261055
transform 1 0 39744 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_410
timestamp 1621261055
transform 1 0 40512 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_418
timestamp 1621261055
transform 1 0 41280 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_407
timestamp 1621261055
transform 1 0 40224 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_411
timestamp 1621261055
transform 1 0 40608 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_414
timestamp 1621261055
transform 1 0 40896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_422
timestamp 1621261055
transform 1 0 41664 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_426
timestamp 1621261055
transform 1 0 42048 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_430
timestamp 1621261055
transform 1 0 42432 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_435
timestamp 1621261055
transform 1 0 42912 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_430
timestamp 1621261055
transform 1 0 42432 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _205_
timestamp 1621261055
transform 1 0 42624 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_438
timestamp 1621261055
transform 1 0 43200 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_441
timestamp 1621261055
transform 1 0 43488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_439
timestamp 1621261055
transform 1 0 43296 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_423
timestamp 1621261055
transform 1 0 43392 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _181_
timestamp 1621261055
transform 1 0 44736 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_23_449
timestamp 1621261055
transform 1 0 44256 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_457
timestamp 1621261055
transform 1 0 45024 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_446
timestamp 1621261055
transform 1 0 43968 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_457
timestamp 1621261055
transform 1 0 45024 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _220_
timestamp 1621261055
transform -1 0 46272 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_434
timestamp 1621261055
transform 1 0 46080 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_33
timestamp 1621261055
transform -1 0 45984 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_470
timestamp 1621261055
transform 1 0 46272 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_478
timestamp 1621261055
transform 1 0 47040 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_465
timestamp 1621261055
transform 1 0 45792 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_24_467
timestamp 1621261055
transform 1 0 45984 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_469
timestamp 1621261055
transform 1 0 46176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_477
timestamp 1621261055
transform 1 0 46944 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_424
timestamp 1621261055
transform 1 0 48672 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_486
timestamp 1621261055
transform 1 0 47808 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_494
timestamp 1621261055
transform 1 0 48576 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_496
timestamp 1621261055
transform 1 0 48768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_504
timestamp 1621261055
transform 1 0 49536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_485
timestamp 1621261055
transform 1 0 47712 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_493
timestamp 1621261055
transform 1 0 48480 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_501
timestamp 1621261055
transform 1 0 49248 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_435
timestamp 1621261055
transform 1 0 51360 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_512
timestamp 1621261055
transform 1 0 50304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_520
timestamp 1621261055
transform 1 0 51072 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_509
timestamp 1621261055
transform 1 0 50016 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_517
timestamp 1621261055
transform 1 0 50784 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_521
timestamp 1621261055
transform 1 0 51168 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_524
timestamp 1621261055
transform 1 0 51456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_528
timestamp 1621261055
transform 1 0 51840 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_536
timestamp 1621261055
transform 1 0 52608 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_544
timestamp 1621261055
transform 1 0 53376 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_532
timestamp 1621261055
transform 1 0 52224 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_540
timestamp 1621261055
transform 1 0 52992 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_425
timestamp 1621261055
transform 1 0 53952 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_548
timestamp 1621261055
transform 1 0 53760 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_551
timestamp 1621261055
transform 1 0 54048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_559
timestamp 1621261055
transform 1 0 54816 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_567
timestamp 1621261055
transform 1 0 55584 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_548
timestamp 1621261055
transform 1 0 53760 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_556
timestamp 1621261055
transform 1 0 54528 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_564
timestamp 1621261055
transform 1 0 55296 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_436
timestamp 1621261055
transform 1 0 56640 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_575
timestamp 1621261055
transform 1 0 56352 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_583
timestamp 1621261055
transform 1 0 57120 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_572
timestamp 1621261055
transform 1 0 56064 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_576
timestamp 1621261055
transform 1 0 56448 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_579
timestamp 1621261055
transform 1 0 56736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_587
timestamp 1621261055
transform 1 0 57504 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_47
timestamp 1621261055
transform -1 0 58848 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_49
timestamp 1621261055
transform -1 0 58848 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_23_591
timestamp 1621261055
transform 1 0 57888 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_595
timestamp 1621261055
transform 1 0 58272 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_595
timestamp 1621261055
transform 1 0 58272 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_50
timestamp 1621261055
transform 1 0 1152 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_4
timestamp 1621261055
transform 1 0 1536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_12
timestamp 1621261055
transform 1 0 2304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_20
timestamp 1621261055
transform 1 0 3072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_28
timestamp 1621261055
transform 1 0 3840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_36
timestamp 1621261055
transform 1 0 4608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_437
timestamp 1621261055
transform 1 0 6432 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_44
timestamp 1621261055
transform 1 0 5376 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_52
timestamp 1621261055
transform 1 0 6144 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_54
timestamp 1621261055
transform 1 0 6336 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_56
timestamp 1621261055
transform 1 0 6528 0 1 19314
box -38 -49 806 715
use OR2X1  OR2X1
timestamp 1624196784
transform 1 0 7680 0 1 19314
box 0 -48 1152 714
use sky130_fd_sc_ls__diode_2  ANTENNA_84
timestamp 1621261055
transform 1 0 7488 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_64
timestamp 1621261055
transform 1 0 7296 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_80
timestamp 1621261055
transform 1 0 8832 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_88
timestamp 1621261055
transform 1 0 9600 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_96
timestamp 1621261055
transform 1 0 10368 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_104
timestamp 1621261055
transform 1 0 11136 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _052_
timestamp 1621261055
transform 1 0 12192 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_438
timestamp 1621261055
transform 1 0 11712 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_73
timestamp 1621261055
transform 1 0 12000 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_108
timestamp 1621261055
transform 1 0 11520 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_111
timestamp 1621261055
transform 1 0 11808 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_118
timestamp 1621261055
transform 1 0 12480 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_126
timestamp 1621261055
transform 1 0 13248 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_134
timestamp 1621261055
transform 1 0 14016 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_142
timestamp 1621261055
transform 1 0 14784 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_439
timestamp 1621261055
transform 1 0 16992 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_150
timestamp 1621261055
transform 1 0 15552 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_158
timestamp 1621261055
transform 1 0 16320 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_162
timestamp 1621261055
transform 1 0 16704 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_164
timestamp 1621261055
transform 1 0 16896 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_166
timestamp 1621261055
transform 1 0 17088 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _210_
timestamp 1621261055
transform 1 0 18720 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_25_174
timestamp 1621261055
transform 1 0 17856 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_25_182
timestamp 1621261055
transform 1 0 18624 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_186
timestamp 1621261055
transform 1 0 19008 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_194
timestamp 1621261055
transform 1 0 19776 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_202
timestamp 1621261055
transform 1 0 20544 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_210
timestamp 1621261055
transform 1 0 21312 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_440
timestamp 1621261055
transform 1 0 22272 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_218
timestamp 1621261055
transform 1 0 22080 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_221
timestamp 1621261055
transform 1 0 22368 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_229
timestamp 1621261055
transform 1 0 23136 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_237
timestamp 1621261055
transform 1 0 23904 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_245
timestamp 1621261055
transform 1 0 24672 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_253
timestamp 1621261055
transform 1 0 25440 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_261
timestamp 1621261055
transform 1 0 26208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_269
timestamp 1621261055
transform 1 0 26976 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_273
timestamp 1621261055
transform 1 0 27360 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_441
timestamp 1621261055
transform 1 0 27552 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_276
timestamp 1621261055
transform 1 0 27648 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_284
timestamp 1621261055
transform 1 0 28416 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_292
timestamp 1621261055
transform 1 0 29184 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _066_
timestamp 1621261055
transform 1 0 30336 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_25_300
timestamp 1621261055
transform 1 0 29952 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_307
timestamp 1621261055
transform 1 0 30624 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_315
timestamp 1621261055
transform 1 0 31392 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_442
timestamp 1621261055
transform 1 0 32832 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_323
timestamp 1621261055
transform 1 0 32160 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_327
timestamp 1621261055
transform 1 0 32544 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_329
timestamp 1621261055
transform 1 0 32736 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_331
timestamp 1621261055
transform 1 0 32928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_339
timestamp 1621261055
transform 1 0 33696 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_347
timestamp 1621261055
transform 1 0 34464 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_355
timestamp 1621261055
transform 1 0 35232 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_363
timestamp 1621261055
transform 1 0 36000 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_371
timestamp 1621261055
transform 1 0 36768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_443
timestamp 1621261055
transform 1 0 38112 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_379
timestamp 1621261055
transform 1 0 37536 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_383
timestamp 1621261055
transform 1 0 37920 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_386
timestamp 1621261055
transform 1 0 38208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_394
timestamp 1621261055
transform 1 0 38976 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_402
timestamp 1621261055
transform 1 0 39744 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_410
timestamp 1621261055
transform 1 0 40512 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_418
timestamp 1621261055
transform 1 0 41280 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_444
timestamp 1621261055
transform 1 0 43392 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_426
timestamp 1621261055
transform 1 0 42048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_434
timestamp 1621261055
transform 1 0 42816 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_438
timestamp 1621261055
transform 1 0 43200 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_441
timestamp 1621261055
transform 1 0 43488 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_449
timestamp 1621261055
transform 1 0 44256 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_457
timestamp 1621261055
transform 1 0 45024 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_465
timestamp 1621261055
transform 1 0 45792 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_473
timestamp 1621261055
transform 1 0 46560 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_481
timestamp 1621261055
transform 1 0 47328 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_445
timestamp 1621261055
transform 1 0 48672 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_489
timestamp 1621261055
transform 1 0 48096 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_493
timestamp 1621261055
transform 1 0 48480 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_496
timestamp 1621261055
transform 1 0 48768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_504
timestamp 1621261055
transform 1 0 49536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_512
timestamp 1621261055
transform 1 0 50304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_520
timestamp 1621261055
transform 1 0 51072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_528
timestamp 1621261055
transform 1 0 51840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_536
timestamp 1621261055
transform 1 0 52608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_544
timestamp 1621261055
transform 1 0 53376 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_446
timestamp 1621261055
transform 1 0 53952 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_548
timestamp 1621261055
transform 1 0 53760 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_551
timestamp 1621261055
transform 1 0 54048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_559
timestamp 1621261055
transform 1 0 54816 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_567
timestamp 1621261055
transform 1 0 55584 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_575
timestamp 1621261055
transform 1 0 56352 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_583
timestamp 1621261055
transform 1 0 57120 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_51
timestamp 1621261055
transform -1 0 58848 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_25_591
timestamp 1621261055
transform 1 0 57888 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_595
timestamp 1621261055
transform 1 0 58272 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_52
timestamp 1621261055
transform 1 0 1152 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_26_4
timestamp 1621261055
transform 1 0 1536 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_12
timestamp 1621261055
transform 1 0 2304 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_20
timestamp 1621261055
transform 1 0 3072 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_447
timestamp 1621261055
transform 1 0 3840 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_29
timestamp 1621261055
transform 1 0 3936 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_37
timestamp 1621261055
transform 1 0 4704 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_45
timestamp 1621261055
transform 1 0 5472 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_53
timestamp 1621261055
transform 1 0 6240 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_61
timestamp 1621261055
transform 1 0 7008 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_448
timestamp 1621261055
transform 1 0 9120 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_69
timestamp 1621261055
transform 1 0 7776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_77
timestamp 1621261055
transform 1 0 8544 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_81
timestamp 1621261055
transform 1 0 8928 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_26_84
timestamp 1621261055
transform 1 0 9216 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _155_
timestamp 1621261055
transform 1 0 9600 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_91
timestamp 1621261055
transform 1 0 9888 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_99
timestamp 1621261055
transform 1 0 10656 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_107
timestamp 1621261055
transform 1 0 11424 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_115
timestamp 1621261055
transform 1 0 12192 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_123
timestamp 1621261055
transform 1 0 12960 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_449
timestamp 1621261055
transform 1 0 14400 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_131
timestamp 1621261055
transform 1 0 13728 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_135
timestamp 1621261055
transform 1 0 14112 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_137
timestamp 1621261055
transform 1 0 14304 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_139
timestamp 1621261055
transform 1 0 14496 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_147
timestamp 1621261055
transform 1 0 15264 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_155
timestamp 1621261055
transform 1 0 16032 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_163
timestamp 1621261055
transform 1 0 16800 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_171
timestamp 1621261055
transform 1 0 17568 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_179
timestamp 1621261055
transform 1 0 18336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_187
timestamp 1621261055
transform 1 0 19104 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_450
timestamp 1621261055
transform 1 0 19680 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_191
timestamp 1621261055
transform 1 0 19488 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_194
timestamp 1621261055
transform 1 0 19776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_202
timestamp 1621261055
transform 1 0 20544 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_210
timestamp 1621261055
transform 1 0 21312 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _000_
timestamp 1621261055
transform 1 0 22176 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_4
timestamp 1621261055
transform 1 0 21984 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_214
timestamp 1621261055
transform 1 0 21696 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_216
timestamp 1621261055
transform 1 0 21888 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_222
timestamp 1621261055
transform 1 0 22464 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_230
timestamp 1621261055
transform 1 0 23232 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_451
timestamp 1621261055
transform 1 0 24960 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_238
timestamp 1621261055
transform 1 0 24000 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_246
timestamp 1621261055
transform 1 0 24768 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_249
timestamp 1621261055
transform 1 0 25056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_257
timestamp 1621261055
transform 1 0 25824 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_265
timestamp 1621261055
transform 1 0 26592 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_273
timestamp 1621261055
transform 1 0 27360 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_281
timestamp 1621261055
transform 1 0 28128 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_289
timestamp 1621261055
transform 1 0 28896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_452
timestamp 1621261055
transform 1 0 30240 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_297
timestamp 1621261055
transform 1 0 29664 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_301
timestamp 1621261055
transform 1 0 30048 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_304
timestamp 1621261055
transform 1 0 30336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_312
timestamp 1621261055
transform 1 0 31104 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_320
timestamp 1621261055
transform 1 0 31872 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_328
timestamp 1621261055
transform 1 0 32640 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_336
timestamp 1621261055
transform 1 0 33408 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_344
timestamp 1621261055
transform 1 0 34176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_352
timestamp 1621261055
transform 1 0 34944 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_356
timestamp 1621261055
transform 1 0 35328 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_453
timestamp 1621261055
transform 1 0 35520 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_359
timestamp 1621261055
transform 1 0 35616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_367
timestamp 1621261055
transform 1 0 36384 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_375
timestamp 1621261055
transform 1 0 37152 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_383
timestamp 1621261055
transform 1 0 37920 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_391
timestamp 1621261055
transform 1 0 38688 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_399
timestamp 1621261055
transform 1 0 39456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_454
timestamp 1621261055
transform 1 0 40800 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_407
timestamp 1621261055
transform 1 0 40224 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_411
timestamp 1621261055
transform 1 0 40608 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_414
timestamp 1621261055
transform 1 0 40896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_422
timestamp 1621261055
transform 1 0 41664 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_430
timestamp 1621261055
transform 1 0 42432 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_438
timestamp 1621261055
transform 1 0 43200 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _126_
timestamp 1621261055
transform 1 0 44928 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_446
timestamp 1621261055
transform 1 0 43968 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_454
timestamp 1621261055
transform 1 0 44736 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_459
timestamp 1621261055
transform 1 0 45216 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_455
timestamp 1621261055
transform 1 0 46080 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_26_467
timestamp 1621261055
transform 1 0 45984 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_469
timestamp 1621261055
transform 1 0 46176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_477
timestamp 1621261055
transform 1 0 46944 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _173_
timestamp 1621261055
transform 1 0 49440 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_485
timestamp 1621261055
transform 1 0 47712 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_493
timestamp 1621261055
transform 1 0 48480 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_501
timestamp 1621261055
transform 1 0 49248 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_456
timestamp 1621261055
transform 1 0 51360 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_506
timestamp 1621261055
transform 1 0 49728 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_514
timestamp 1621261055
transform 1 0 50496 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_26_522
timestamp 1621261055
transform 1 0 51264 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_524
timestamp 1621261055
transform 1 0 51456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_532
timestamp 1621261055
transform 1 0 52224 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_540
timestamp 1621261055
transform 1 0 52992 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_548
timestamp 1621261055
transform 1 0 53760 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_556
timestamp 1621261055
transform 1 0 54528 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_564
timestamp 1621261055
transform 1 0 55296 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_457
timestamp 1621261055
transform 1 0 56640 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_572
timestamp 1621261055
transform 1 0 56064 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_576
timestamp 1621261055
transform 1 0 56448 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_579
timestamp 1621261055
transform 1 0 56736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_587
timestamp 1621261055
transform 1 0 57504 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_53
timestamp 1621261055
transform -1 0 58848 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_595
timestamp 1621261055
transform 1 0 58272 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_54
timestamp 1621261055
transform 1 0 1152 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_4
timestamp 1621261055
transform 1 0 1536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_12
timestamp 1621261055
transform 1 0 2304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_20
timestamp 1621261055
transform 1 0 3072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_28
timestamp 1621261055
transform 1 0 3840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_36
timestamp 1621261055
transform 1 0 4608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_458
timestamp 1621261055
transform 1 0 6432 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_44
timestamp 1621261055
transform 1 0 5376 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_52
timestamp 1621261055
transform 1 0 6144 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_54
timestamp 1621261055
transform 1 0 6336 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_56
timestamp 1621261055
transform 1 0 6528 0 1 20646
box -38 -49 806 715
use OR2X2  OR2X2
timestamp 1624196784
transform 1 0 7680 0 1 20646
box 0 -48 1152 714
use sky130_fd_sc_ls__diode_2  ANTENNA_89
timestamp 1621261055
transform 1 0 7488 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_64
timestamp 1621261055
transform 1 0 7296 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_80
timestamp 1621261055
transform 1 0 8832 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_88
timestamp 1621261055
transform 1 0 9600 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_96
timestamp 1621261055
transform 1 0 10368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_104
timestamp 1621261055
transform 1 0 11136 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_459
timestamp 1621261055
transform 1 0 11712 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_108
timestamp 1621261055
transform 1 0 11520 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_111
timestamp 1621261055
transform 1 0 11808 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_119
timestamp 1621261055
transform 1 0 12576 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_127
timestamp 1621261055
transform 1 0 13344 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_135
timestamp 1621261055
transform 1 0 14112 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_143
timestamp 1621261055
transform 1 0 14880 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_460
timestamp 1621261055
transform 1 0 16992 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_151
timestamp 1621261055
transform 1 0 15648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_159
timestamp 1621261055
transform 1 0 16416 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_163
timestamp 1621261055
transform 1 0 16800 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_166
timestamp 1621261055
transform 1 0 17088 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_174
timestamp 1621261055
transform 1 0 17856 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_182
timestamp 1621261055
transform 1 0 18624 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_190
timestamp 1621261055
transform 1 0 19392 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_198
timestamp 1621261055
transform 1 0 20160 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_206
timestamp 1621261055
transform 1 0 20928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_461
timestamp 1621261055
transform 1 0 22272 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_214
timestamp 1621261055
transform 1 0 21696 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_218
timestamp 1621261055
transform 1 0 22080 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_221
timestamp 1621261055
transform 1 0 22368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_229
timestamp 1621261055
transform 1 0 23136 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_237
timestamp 1621261055
transform 1 0 23904 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_245
timestamp 1621261055
transform 1 0 24672 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_253
timestamp 1621261055
transform 1 0 25440 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_261
timestamp 1621261055
transform 1 0 26208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_269
timestamp 1621261055
transform 1 0 26976 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_273
timestamp 1621261055
transform 1 0 27360 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_462
timestamp 1621261055
transform 1 0 27552 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_276
timestamp 1621261055
transform 1 0 27648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_284
timestamp 1621261055
transform 1 0 28416 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_292
timestamp 1621261055
transform 1 0 29184 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_300
timestamp 1621261055
transform 1 0 29952 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_308
timestamp 1621261055
transform 1 0 30720 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _140_
timestamp 1621261055
transform 1 0 33312 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_463
timestamp 1621261055
transform 1 0 32832 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_316
timestamp 1621261055
transform 1 0 31488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_324
timestamp 1621261055
transform 1 0 32256 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_328
timestamp 1621261055
transform 1 0 32640 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_27_331
timestamp 1621261055
transform 1 0 32928 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_338
timestamp 1621261055
transform 1 0 33600 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_346
timestamp 1621261055
transform 1 0 34368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_354
timestamp 1621261055
transform 1 0 35136 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_362
timestamp 1621261055
transform 1 0 35904 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_370
timestamp 1621261055
transform 1 0 36672 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_378
timestamp 1621261055
transform 1 0 37440 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_464
timestamp 1621261055
transform 1 0 38112 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_382
timestamp 1621261055
transform 1 0 37824 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_384
timestamp 1621261055
transform 1 0 38016 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_386
timestamp 1621261055
transform 1 0 38208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_394
timestamp 1621261055
transform 1 0 38976 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_402
timestamp 1621261055
transform 1 0 39744 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_410
timestamp 1621261055
transform 1 0 40512 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_418
timestamp 1621261055
transform 1 0 41280 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_465
timestamp 1621261055
transform 1 0 43392 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_426
timestamp 1621261055
transform 1 0 42048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_434
timestamp 1621261055
transform 1 0 42816 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_438
timestamp 1621261055
transform 1 0 43200 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_441
timestamp 1621261055
transform 1 0 43488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_449
timestamp 1621261055
transform 1 0 44256 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_457
timestamp 1621261055
transform 1 0 45024 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_465
timestamp 1621261055
transform 1 0 45792 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_473
timestamp 1621261055
transform 1 0 46560 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_481
timestamp 1621261055
transform 1 0 47328 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_466
timestamp 1621261055
transform 1 0 48672 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_489
timestamp 1621261055
transform 1 0 48096 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_493
timestamp 1621261055
transform 1 0 48480 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_496
timestamp 1621261055
transform 1 0 48768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_504
timestamp 1621261055
transform 1 0 49536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _222_
timestamp 1621261055
transform -1 0 51168 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_2
timestamp 1621261055
transform -1 0 50880 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_27_512
timestamp 1621261055
transform 1 0 50304 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_521
timestamp 1621261055
transform 1 0 51168 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_529
timestamp 1621261055
transform 1 0 51936 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_537
timestamp 1621261055
transform 1 0 52704 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_545
timestamp 1621261055
transform 1 0 53472 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_467
timestamp 1621261055
transform 1 0 53952 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_27_549
timestamp 1621261055
transform 1 0 53856 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_551
timestamp 1621261055
transform 1 0 54048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_559
timestamp 1621261055
transform 1 0 54816 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_567
timestamp 1621261055
transform 1 0 55584 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_575
timestamp 1621261055
transform 1 0 56352 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_583
timestamp 1621261055
transform 1 0 57120 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_55
timestamp 1621261055
transform -1 0 58848 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_27_591
timestamp 1621261055
transform 1 0 57888 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_595
timestamp 1621261055
transform 1 0 58272 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_56
timestamp 1621261055
transform 1 0 1152 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_28_4
timestamp 1621261055
transform 1 0 1536 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_12
timestamp 1621261055
transform 1 0 2304 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_20
timestamp 1621261055
transform 1 0 3072 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_468
timestamp 1621261055
transform 1 0 3840 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_29
timestamp 1621261055
transform 1 0 3936 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_37
timestamp 1621261055
transform 1 0 4704 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_45
timestamp 1621261055
transform 1 0 5472 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_53
timestamp 1621261055
transform 1 0 6240 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_61
timestamp 1621261055
transform 1 0 7008 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_469
timestamp 1621261055
transform 1 0 9120 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_69
timestamp 1621261055
transform 1 0 7776 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_77
timestamp 1621261055
transform 1 0 8544 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_81
timestamp 1621261055
transform 1 0 8928 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_84
timestamp 1621261055
transform 1 0 9216 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_92
timestamp 1621261055
transform 1 0 9984 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_100
timestamp 1621261055
transform 1 0 10752 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_108
timestamp 1621261055
transform 1 0 11520 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_116
timestamp 1621261055
transform 1 0 12288 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_124
timestamp 1621261055
transform 1 0 13056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_470
timestamp 1621261055
transform 1 0 14400 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_132
timestamp 1621261055
transform 1 0 13824 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_136
timestamp 1621261055
transform 1 0 14208 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_139
timestamp 1621261055
transform 1 0 14496 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_147
timestamp 1621261055
transform 1 0 15264 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_155
timestamp 1621261055
transform 1 0 16032 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_163
timestamp 1621261055
transform 1 0 16800 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_171
timestamp 1621261055
transform 1 0 17568 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_179
timestamp 1621261055
transform 1 0 18336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_187
timestamp 1621261055
transform 1 0 19104 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_471
timestamp 1621261055
transform 1 0 19680 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_191
timestamp 1621261055
transform 1 0 19488 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_194
timestamp 1621261055
transform 1 0 19776 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_202
timestamp 1621261055
transform 1 0 20544 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_210
timestamp 1621261055
transform 1 0 21312 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_218
timestamp 1621261055
transform 1 0 22080 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_226
timestamp 1621261055
transform 1 0 22848 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_472
timestamp 1621261055
transform 1 0 24960 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_234
timestamp 1621261055
transform 1 0 23616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_242
timestamp 1621261055
transform 1 0 24384 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_246
timestamp 1621261055
transform 1 0 24768 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_249
timestamp 1621261055
transform 1 0 25056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_257
timestamp 1621261055
transform 1 0 25824 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_265
timestamp 1621261055
transform 1 0 26592 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_273
timestamp 1621261055
transform 1 0 27360 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_281
timestamp 1621261055
transform 1 0 28128 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_289
timestamp 1621261055
transform 1 0 28896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_473
timestamp 1621261055
transform 1 0 30240 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_297
timestamp 1621261055
transform 1 0 29664 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_301
timestamp 1621261055
transform 1 0 30048 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_304
timestamp 1621261055
transform 1 0 30336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_312
timestamp 1621261055
transform 1 0 31104 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_320
timestamp 1621261055
transform 1 0 31872 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_328
timestamp 1621261055
transform 1 0 32640 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_336
timestamp 1621261055
transform 1 0 33408 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_344
timestamp 1621261055
transform 1 0 34176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_352
timestamp 1621261055
transform 1 0 34944 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_356
timestamp 1621261055
transform 1 0 35328 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_474
timestamp 1621261055
transform 1 0 35520 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_359
timestamp 1621261055
transform 1 0 35616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_367
timestamp 1621261055
transform 1 0 36384 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_375
timestamp 1621261055
transform 1 0 37152 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_383
timestamp 1621261055
transform 1 0 37920 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_391
timestamp 1621261055
transform 1 0 38688 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_399
timestamp 1621261055
transform 1 0 39456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_475
timestamp 1621261055
transform 1 0 40800 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_407
timestamp 1621261055
transform 1 0 40224 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_411
timestamp 1621261055
transform 1 0 40608 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_414
timestamp 1621261055
transform 1 0 40896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_422
timestamp 1621261055
transform 1 0 41664 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_430
timestamp 1621261055
transform 1 0 42432 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_438
timestamp 1621261055
transform 1 0 43200 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_446
timestamp 1621261055
transform 1 0 43968 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_454
timestamp 1621261055
transform 1 0 44736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_462
timestamp 1621261055
transform 1 0 45504 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_476
timestamp 1621261055
transform 1 0 46080 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_466
timestamp 1621261055
transform 1 0 45888 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_469
timestamp 1621261055
transform 1 0 46176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_477
timestamp 1621261055
transform 1 0 46944 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_485
timestamp 1621261055
transform 1 0 47712 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_493
timestamp 1621261055
transform 1 0 48480 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_501
timestamp 1621261055
transform 1 0 49248 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_477
timestamp 1621261055
transform 1 0 51360 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_509
timestamp 1621261055
transform 1 0 50016 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_517
timestamp 1621261055
transform 1 0 50784 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_521
timestamp 1621261055
transform 1 0 51168 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_524
timestamp 1621261055
transform 1 0 51456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_532
timestamp 1621261055
transform 1 0 52224 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_540
timestamp 1621261055
transform 1 0 52992 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_548
timestamp 1621261055
transform 1 0 53760 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_556
timestamp 1621261055
transform 1 0 54528 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_564
timestamp 1621261055
transform 1 0 55296 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_478
timestamp 1621261055
transform 1 0 56640 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_572
timestamp 1621261055
transform 1 0 56064 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_576
timestamp 1621261055
transform 1 0 56448 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_579
timestamp 1621261055
transform 1 0 56736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_587
timestamp 1621261055
transform 1 0 57504 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_57
timestamp 1621261055
transform -1 0 58848 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_595
timestamp 1621261055
transform 1 0 58272 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_58
timestamp 1621261055
transform 1 0 1152 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_29_4
timestamp 1621261055
transform 1 0 1536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_12
timestamp 1621261055
transform 1 0 2304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_20
timestamp 1621261055
transform 1 0 3072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_28
timestamp 1621261055
transform 1 0 3840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_36
timestamp 1621261055
transform 1 0 4608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_479
timestamp 1621261055
transform 1 0 6432 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_44
timestamp 1621261055
transform 1 0 5376 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_52
timestamp 1621261055
transform 1 0 6144 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_54
timestamp 1621261055
transform 1 0 6336 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_56
timestamp 1621261055
transform 1 0 6528 0 1 21978
box -38 -49 806 715
use XOR2X1  XOR2X1
timestamp 1624196784
transform 1 0 7680 0 1 21978
box 0 -48 2016 714
use sky130_fd_sc_ls__decap_4  FILLER_29_64
timestamp 1621261055
transform 1 0 7296 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_29_89
timestamp 1621261055
transform 1 0 9696 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_97
timestamp 1621261055
transform 1 0 10464 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_105
timestamp 1621261055
transform 1 0 11232 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_480
timestamp 1621261055
transform 1 0 11712 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_29_109
timestamp 1621261055
transform 1 0 11616 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_111
timestamp 1621261055
transform 1 0 11808 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_119
timestamp 1621261055
transform 1 0 12576 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_127
timestamp 1621261055
transform 1 0 13344 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_135
timestamp 1621261055
transform 1 0 14112 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_143
timestamp 1621261055
transform 1 0 14880 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_29_147
timestamp 1621261055
transform 1 0 15264 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _118_
timestamp 1621261055
transform 1 0 15360 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_481
timestamp 1621261055
transform 1 0 16992 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_151
timestamp 1621261055
transform 1 0 15648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_159
timestamp 1621261055
transform 1 0 16416 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_163
timestamp 1621261055
transform 1 0 16800 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_166
timestamp 1621261055
transform 1 0 17088 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_174
timestamp 1621261055
transform 1 0 17856 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_182
timestamp 1621261055
transform 1 0 18624 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_190
timestamp 1621261055
transform 1 0 19392 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_198
timestamp 1621261055
transform 1 0 20160 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_206
timestamp 1621261055
transform 1 0 20928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_482
timestamp 1621261055
transform 1 0 22272 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_214
timestamp 1621261055
transform 1 0 21696 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_218
timestamp 1621261055
transform 1 0 22080 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_221
timestamp 1621261055
transform 1 0 22368 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_229
timestamp 1621261055
transform 1 0 23136 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_237
timestamp 1621261055
transform 1 0 23904 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_245
timestamp 1621261055
transform 1 0 24672 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _048_
timestamp 1621261055
transform 1 0 26880 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_61
timestamp 1621261055
transform 1 0 26688 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_253
timestamp 1621261055
transform 1 0 25440 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_261
timestamp 1621261055
transform 1 0 26208 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_29_265
timestamp 1621261055
transform 1 0 26592 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_271
timestamp 1621261055
transform 1 0 27168 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_483
timestamp 1621261055
transform 1 0 27552 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_276
timestamp 1621261055
transform 1 0 27648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_284
timestamp 1621261055
transform 1 0 28416 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_292
timestamp 1621261055
transform 1 0 29184 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_300
timestamp 1621261055
transform 1 0 29952 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_308
timestamp 1621261055
transform 1 0 30720 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_484
timestamp 1621261055
transform 1 0 32832 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_316
timestamp 1621261055
transform 1 0 31488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_324
timestamp 1621261055
transform 1 0 32256 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_328
timestamp 1621261055
transform 1 0 32640 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_331
timestamp 1621261055
transform 1 0 32928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_339
timestamp 1621261055
transform 1 0 33696 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_347
timestamp 1621261055
transform 1 0 34464 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_355
timestamp 1621261055
transform 1 0 35232 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_363
timestamp 1621261055
transform 1 0 36000 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_371
timestamp 1621261055
transform 1 0 36768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_485
timestamp 1621261055
transform 1 0 38112 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_379
timestamp 1621261055
transform 1 0 37536 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_383
timestamp 1621261055
transform 1 0 37920 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_386
timestamp 1621261055
transform 1 0 38208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_394
timestamp 1621261055
transform 1 0 38976 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_402
timestamp 1621261055
transform 1 0 39744 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_410
timestamp 1621261055
transform 1 0 40512 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_418
timestamp 1621261055
transform 1 0 41280 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_486
timestamp 1621261055
transform 1 0 43392 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_426
timestamp 1621261055
transform 1 0 42048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_434
timestamp 1621261055
transform 1 0 42816 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_438
timestamp 1621261055
transform 1 0 43200 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_441
timestamp 1621261055
transform 1 0 43488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_449
timestamp 1621261055
transform 1 0 44256 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_457
timestamp 1621261055
transform 1 0 45024 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_465
timestamp 1621261055
transform 1 0 45792 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_473
timestamp 1621261055
transform 1 0 46560 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_481
timestamp 1621261055
transform 1 0 47328 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_487
timestamp 1621261055
transform 1 0 48672 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_489
timestamp 1621261055
transform 1 0 48096 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_493
timestamp 1621261055
transform 1 0 48480 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_496
timestamp 1621261055
transform 1 0 48768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_504
timestamp 1621261055
transform 1 0 49536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_512
timestamp 1621261055
transform 1 0 50304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_520
timestamp 1621261055
transform 1 0 51072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_528
timestamp 1621261055
transform 1 0 51840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_536
timestamp 1621261055
transform 1 0 52608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_544
timestamp 1621261055
transform 1 0 53376 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_488
timestamp 1621261055
transform 1 0 53952 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_548
timestamp 1621261055
transform 1 0 53760 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_551
timestamp 1621261055
transform 1 0 54048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_559
timestamp 1621261055
transform 1 0 54816 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_567
timestamp 1621261055
transform 1 0 55584 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_575
timestamp 1621261055
transform 1 0 56352 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_583
timestamp 1621261055
transform 1 0 57120 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_59
timestamp 1621261055
transform -1 0 58848 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_29_591
timestamp 1621261055
transform 1 0 57888 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_595
timestamp 1621261055
transform 1 0 58272 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_60
timestamp 1621261055
transform 1 0 1152 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_62
timestamp 1621261055
transform 1 0 1152 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_4
timestamp 1621261055
transform 1 0 1536 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_12
timestamp 1621261055
transform 1 0 2304 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_20
timestamp 1621261055
transform 1 0 3072 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_4
timestamp 1621261055
transform 1 0 1536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_12
timestamp 1621261055
transform 1 0 2304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_20
timestamp 1621261055
transform 1 0 3072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_489
timestamp 1621261055
transform 1 0 3840 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_29
timestamp 1621261055
transform 1 0 3936 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_37
timestamp 1621261055
transform 1 0 4704 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_28
timestamp 1621261055
transform 1 0 3840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_36
timestamp 1621261055
transform 1 0 4608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_500
timestamp 1621261055
transform 1 0 6432 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_45
timestamp 1621261055
transform 1 0 5472 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_53
timestamp 1621261055
transform 1 0 6240 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_61
timestamp 1621261055
transform 1 0 7008 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_44
timestamp 1621261055
transform 1 0 5376 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_52
timestamp 1621261055
transform 1 0 6144 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_31_54
timestamp 1621261055
transform 1 0 6336 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_56
timestamp 1621261055
transform 1 0 6528 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_490
timestamp 1621261055
transform 1 0 9120 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_69
timestamp 1621261055
transform 1 0 7776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_77
timestamp 1621261055
transform 1 0 8544 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_81
timestamp 1621261055
transform 1 0 8928 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_84
timestamp 1621261055
transform 1 0 9216 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_64
timestamp 1621261055
transform 1 0 7296 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_72
timestamp 1621261055
transform 1 0 8064 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_80
timestamp 1621261055
transform 1 0 8832 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_92
timestamp 1621261055
transform 1 0 9984 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_100
timestamp 1621261055
transform 1 0 10752 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_88
timestamp 1621261055
transform 1 0 9600 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_96
timestamp 1621261055
transform 1 0 10368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_104
timestamp 1621261055
transform 1 0 11136 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_501
timestamp 1621261055
transform 1 0 11712 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_108
timestamp 1621261055
transform 1 0 11520 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_116
timestamp 1621261055
transform 1 0 12288 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_124
timestamp 1621261055
transform 1 0 13056 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_30_126
timestamp 1621261055
transform 1 0 13248 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_108
timestamp 1621261055
transform 1 0 11520 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_111
timestamp 1621261055
transform 1 0 11808 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_119
timestamp 1621261055
transform 1 0 12576 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _112_
timestamp 1621261055
transform 1 0 13344 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_491
timestamp 1621261055
transform 1 0 14400 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_130
timestamp 1621261055
transform 1 0 13632 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_139
timestamp 1621261055
transform 1 0 14496 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_147
timestamp 1621261055
transform 1 0 15264 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_127
timestamp 1621261055
transform 1 0 13344 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_135
timestamp 1621261055
transform 1 0 14112 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_143
timestamp 1621261055
transform 1 0 14880 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_502
timestamp 1621261055
transform 1 0 16992 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_155
timestamp 1621261055
transform 1 0 16032 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_163
timestamp 1621261055
transform 1 0 16800 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_151
timestamp 1621261055
transform 1 0 15648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_159
timestamp 1621261055
transform 1 0 16416 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_163
timestamp 1621261055
transform 1 0 16800 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_166
timestamp 1621261055
transform 1 0 17088 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _142_
timestamp 1621261055
transform 1 0 17568 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_30_174
timestamp 1621261055
transform 1 0 17856 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_182
timestamp 1621261055
transform 1 0 18624 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_174
timestamp 1621261055
transform 1 0 17856 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_182
timestamp 1621261055
transform 1 0 18624 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_492
timestamp 1621261055
transform 1 0 19680 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_190
timestamp 1621261055
transform 1 0 19392 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_30_192
timestamp 1621261055
transform 1 0 19584 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_194
timestamp 1621261055
transform 1 0 19776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_202
timestamp 1621261055
transform 1 0 20544 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_210
timestamp 1621261055
transform 1 0 21312 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_190
timestamp 1621261055
transform 1 0 19392 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_198
timestamp 1621261055
transform 1 0 20160 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_206
timestamp 1621261055
transform 1 0 20928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_503
timestamp 1621261055
transform 1 0 22272 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_218
timestamp 1621261055
transform 1 0 22080 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_226
timestamp 1621261055
transform 1 0 22848 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_214
timestamp 1621261055
transform 1 0 21696 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_218
timestamp 1621261055
transform 1 0 22080 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_221
timestamp 1621261055
transform 1 0 22368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_229
timestamp 1621261055
transform 1 0 23136 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_493
timestamp 1621261055
transform 1 0 24960 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_234
timestamp 1621261055
transform 1 0 23616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_242
timestamp 1621261055
transform 1 0 24384 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_246
timestamp 1621261055
transform 1 0 24768 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_249
timestamp 1621261055
transform 1 0 25056 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_237
timestamp 1621261055
transform 1 0 23904 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_245
timestamp 1621261055
transform 1 0 24672 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _187_
timestamp 1621261055
transform 1 0 26688 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_30_257
timestamp 1621261055
transform 1 0 25824 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_265
timestamp 1621261055
transform 1 0 26592 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_269
timestamp 1621261055
transform 1 0 26976 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_253
timestamp 1621261055
transform 1 0 25440 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_261
timestamp 1621261055
transform 1 0 26208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_269
timestamp 1621261055
transform 1 0 26976 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_273
timestamp 1621261055
transform 1 0 27360 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_504
timestamp 1621261055
transform 1 0 27552 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_277
timestamp 1621261055
transform 1 0 27744 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_285
timestamp 1621261055
transform 1 0 28512 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_293
timestamp 1621261055
transform 1 0 29280 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_276
timestamp 1621261055
transform 1 0 27648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_284
timestamp 1621261055
transform 1 0 28416 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_292
timestamp 1621261055
transform 1 0 29184 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _169_
timestamp 1621261055
transform 1 0 30720 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_494
timestamp 1621261055
transform 1 0 30240 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_301
timestamp 1621261055
transform 1 0 30048 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_304
timestamp 1621261055
transform 1 0 30336 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_311
timestamp 1621261055
transform 1 0 31008 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_300
timestamp 1621261055
transform 1 0 29952 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_308
timestamp 1621261055
transform 1 0 30720 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_505
timestamp 1621261055
transform 1 0 32832 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_319
timestamp 1621261055
transform 1 0 31776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_327
timestamp 1621261055
transform 1 0 32544 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_335
timestamp 1621261055
transform 1 0 33312 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_316
timestamp 1621261055
transform 1 0 31488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_324
timestamp 1621261055
transform 1 0 32256 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_328
timestamp 1621261055
transform 1 0 32640 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_331
timestamp 1621261055
transform 1 0 32928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_343
timestamp 1621261055
transform 1 0 34080 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_351
timestamp 1621261055
transform 1 0 34848 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_355
timestamp 1621261055
transform 1 0 35232 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_30_357
timestamp 1621261055
transform 1 0 35424 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_339
timestamp 1621261055
transform 1 0 33696 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_347
timestamp 1621261055
transform 1 0 34464 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_355
timestamp 1621261055
transform 1 0 35232 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_495
timestamp 1621261055
transform 1 0 35520 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_359
timestamp 1621261055
transform 1 0 35616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_367
timestamp 1621261055
transform 1 0 36384 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_375
timestamp 1621261055
transform 1 0 37152 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_363
timestamp 1621261055
transform 1 0 36000 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_371
timestamp 1621261055
transform 1 0 36768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_386
timestamp 1621261055
transform 1 0 38208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_383
timestamp 1621261055
transform 1 0 37920 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_379
timestamp 1621261055
transform 1 0 37536 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_30_383
timestamp 1621261055
transform 1 0 37920 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_506
timestamp 1621261055
transform 1 0 38112 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_394
timestamp 1621261055
transform 1 0 38976 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_393
timestamp 1621261055
transform 1 0 38880 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_389
timestamp 1621261055
transform 1 0 38496 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_387
timestamp 1621261055
transform 1 0 38304 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _164_
timestamp 1621261055
transform 1 0 38592 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _034_
timestamp 1621261055
transform -1 0 41568 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_496
timestamp 1621261055
transform 1 0 40800 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_37
timestamp 1621261055
transform -1 0 41280 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_401
timestamp 1621261055
transform 1 0 39648 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_409
timestamp 1621261055
transform 1 0 40416 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_414
timestamp 1621261055
transform 1 0 40896 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_402
timestamp 1621261055
transform 1 0 39744 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_410
timestamp 1621261055
transform 1 0 40512 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_418
timestamp 1621261055
transform 1 0 41280 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_507
timestamp 1621261055
transform 1 0 43392 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_421
timestamp 1621261055
transform 1 0 41568 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_429
timestamp 1621261055
transform 1 0 42336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_437
timestamp 1621261055
transform 1 0 43104 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_426
timestamp 1621261055
transform 1 0 42048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_434
timestamp 1621261055
transform 1 0 42816 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_438
timestamp 1621261055
transform 1 0 43200 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_441
timestamp 1621261055
transform 1 0 43488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_445
timestamp 1621261055
transform 1 0 43872 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_453
timestamp 1621261055
transform 1 0 44640 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_461
timestamp 1621261055
transform 1 0 45408 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_449
timestamp 1621261055
transform 1 0 44256 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_457
timestamp 1621261055
transform 1 0 45024 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_497
timestamp 1621261055
transform 1 0 46080 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_465
timestamp 1621261055
transform 1 0 45792 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_30_467
timestamp 1621261055
transform 1 0 45984 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_469
timestamp 1621261055
transform 1 0 46176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_477
timestamp 1621261055
transform 1 0 46944 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_465
timestamp 1621261055
transform 1 0 45792 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_473
timestamp 1621261055
transform 1 0 46560 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_481
timestamp 1621261055
transform 1 0 47328 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_508
timestamp 1621261055
transform 1 0 48672 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_485
timestamp 1621261055
transform 1 0 47712 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_493
timestamp 1621261055
transform 1 0 48480 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_501
timestamp 1621261055
transform 1 0 49248 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_489
timestamp 1621261055
transform 1 0 48096 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_493
timestamp 1621261055
transform 1 0 48480 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_496
timestamp 1621261055
transform 1 0 48768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_504
timestamp 1621261055
transform 1 0 49536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_498
timestamp 1621261055
transform 1 0 51360 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_509
timestamp 1621261055
transform 1 0 50016 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_517
timestamp 1621261055
transform 1 0 50784 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_521
timestamp 1621261055
transform 1 0 51168 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_524
timestamp 1621261055
transform 1 0 51456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_512
timestamp 1621261055
transform 1 0 50304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_520
timestamp 1621261055
transform 1 0 51072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_532
timestamp 1621261055
transform 1 0 52224 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_540
timestamp 1621261055
transform 1 0 52992 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_528
timestamp 1621261055
transform 1 0 51840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_536
timestamp 1621261055
transform 1 0 52608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_544
timestamp 1621261055
transform 1 0 53376 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_509
timestamp 1621261055
transform 1 0 53952 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_548
timestamp 1621261055
transform 1 0 53760 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_556
timestamp 1621261055
transform 1 0 54528 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_564
timestamp 1621261055
transform 1 0 55296 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_548
timestamp 1621261055
transform 1 0 53760 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_551
timestamp 1621261055
transform 1 0 54048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_559
timestamp 1621261055
transform 1 0 54816 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_567
timestamp 1621261055
transform 1 0 55584 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_499
timestamp 1621261055
transform 1 0 56640 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_572
timestamp 1621261055
transform 1 0 56064 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_576
timestamp 1621261055
transform 1 0 56448 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_579
timestamp 1621261055
transform 1 0 56736 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_587
timestamp 1621261055
transform 1 0 57504 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_575
timestamp 1621261055
transform 1 0 56352 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_583
timestamp 1621261055
transform 1 0 57120 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_61
timestamp 1621261055
transform -1 0 58848 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_63
timestamp 1621261055
transform -1 0 58848 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_595
timestamp 1621261055
transform 1 0 58272 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_591
timestamp 1621261055
transform 1 0 57888 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_595
timestamp 1621261055
transform 1 0 58272 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_64
timestamp 1621261055
transform 1 0 1152 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_32_4
timestamp 1621261055
transform 1 0 1536 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_12
timestamp 1621261055
transform 1 0 2304 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_20
timestamp 1621261055
transform 1 0 3072 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_510
timestamp 1621261055
transform 1 0 3840 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_29
timestamp 1621261055
transform 1 0 3936 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_37
timestamp 1621261055
transform 1 0 4704 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_45
timestamp 1621261055
transform 1 0 5472 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_53
timestamp 1621261055
transform 1 0 6240 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_61
timestamp 1621261055
transform 1 0 7008 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_511
timestamp 1621261055
transform 1 0 9120 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_69
timestamp 1621261055
transform 1 0 7776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_77
timestamp 1621261055
transform 1 0 8544 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_81
timestamp 1621261055
transform 1 0 8928 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_84
timestamp 1621261055
transform 1 0 9216 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_92
timestamp 1621261055
transform 1 0 9984 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_100
timestamp 1621261055
transform 1 0 10752 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_108
timestamp 1621261055
transform 1 0 11520 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_116
timestamp 1621261055
transform 1 0 12288 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_124
timestamp 1621261055
transform 1 0 13056 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_512
timestamp 1621261055
transform 1 0 14400 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_132
timestamp 1621261055
transform 1 0 13824 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_136
timestamp 1621261055
transform 1 0 14208 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_139
timestamp 1621261055
transform 1 0 14496 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_147
timestamp 1621261055
transform 1 0 15264 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_155
timestamp 1621261055
transform 1 0 16032 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_163
timestamp 1621261055
transform 1 0 16800 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_171
timestamp 1621261055
transform 1 0 17568 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_179
timestamp 1621261055
transform 1 0 18336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_187
timestamp 1621261055
transform 1 0 19104 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_513
timestamp 1621261055
transform 1 0 19680 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_191
timestamp 1621261055
transform 1 0 19488 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_194
timestamp 1621261055
transform 1 0 19776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_202
timestamp 1621261055
transform 1 0 20544 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_210
timestamp 1621261055
transform 1 0 21312 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_218
timestamp 1621261055
transform 1 0 22080 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_226
timestamp 1621261055
transform 1 0 22848 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_514
timestamp 1621261055
transform 1 0 24960 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_234
timestamp 1621261055
transform 1 0 23616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_242
timestamp 1621261055
transform 1 0 24384 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_246
timestamp 1621261055
transform 1 0 24768 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_249
timestamp 1621261055
transform 1 0 25056 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_257
timestamp 1621261055
transform 1 0 25824 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_265
timestamp 1621261055
transform 1 0 26592 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_273
timestamp 1621261055
transform 1 0 27360 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_281
timestamp 1621261055
transform 1 0 28128 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_289
timestamp 1621261055
transform 1 0 28896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_515
timestamp 1621261055
transform 1 0 30240 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_297
timestamp 1621261055
transform 1 0 29664 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_301
timestamp 1621261055
transform 1 0 30048 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_304
timestamp 1621261055
transform 1 0 30336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_312
timestamp 1621261055
transform 1 0 31104 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_320
timestamp 1621261055
transform 1 0 31872 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_328
timestamp 1621261055
transform 1 0 32640 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_336
timestamp 1621261055
transform 1 0 33408 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_344
timestamp 1621261055
transform 1 0 34176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_352
timestamp 1621261055
transform 1 0 34944 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_356
timestamp 1621261055
transform 1 0 35328 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_516
timestamp 1621261055
transform 1 0 35520 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_359
timestamp 1621261055
transform 1 0 35616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_367
timestamp 1621261055
transform 1 0 36384 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_375
timestamp 1621261055
transform 1 0 37152 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_383
timestamp 1621261055
transform 1 0 37920 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_391
timestamp 1621261055
transform 1 0 38688 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_399
timestamp 1621261055
transform 1 0 39456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_517
timestamp 1621261055
transform 1 0 40800 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_407
timestamp 1621261055
transform 1 0 40224 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_411
timestamp 1621261055
transform 1 0 40608 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_414
timestamp 1621261055
transform 1 0 40896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _025_
timestamp 1621261055
transform -1 0 43104 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_6
timestamp 1621261055
transform -1 0 42816 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_422
timestamp 1621261055
transform 1 0 41664 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_430
timestamp 1621261055
transform 1 0 42432 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_437
timestamp 1621261055
transform 1 0 43104 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_445
timestamp 1621261055
transform 1 0 43872 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_453
timestamp 1621261055
transform 1 0 44640 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_461
timestamp 1621261055
transform 1 0 45408 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_518
timestamp 1621261055
transform 1 0 46080 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_465
timestamp 1621261055
transform 1 0 45792 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_32_467
timestamp 1621261055
transform 1 0 45984 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_469
timestamp 1621261055
transform 1 0 46176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_477
timestamp 1621261055
transform 1 0 46944 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_485
timestamp 1621261055
transform 1 0 47712 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_493
timestamp 1621261055
transform 1 0 48480 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_501
timestamp 1621261055
transform 1 0 49248 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_519
timestamp 1621261055
transform 1 0 51360 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_509
timestamp 1621261055
transform 1 0 50016 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_517
timestamp 1621261055
transform 1 0 50784 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_521
timestamp 1621261055
transform 1 0 51168 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_524
timestamp 1621261055
transform 1 0 51456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_532
timestamp 1621261055
transform 1 0 52224 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_540
timestamp 1621261055
transform 1 0 52992 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_548
timestamp 1621261055
transform 1 0 53760 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_556
timestamp 1621261055
transform 1 0 54528 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_564
timestamp 1621261055
transform 1 0 55296 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_520
timestamp 1621261055
transform 1 0 56640 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_572
timestamp 1621261055
transform 1 0 56064 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_576
timestamp 1621261055
transform 1 0 56448 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_579
timestamp 1621261055
transform 1 0 56736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_587
timestamp 1621261055
transform 1 0 57504 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_65
timestamp 1621261055
transform -1 0 58848 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_595
timestamp 1621261055
transform 1 0 58272 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_66
timestamp 1621261055
transform 1 0 1152 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_4
timestamp 1621261055
transform 1 0 1536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_12
timestamp 1621261055
transform 1 0 2304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_20
timestamp 1621261055
transform 1 0 3072 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_28
timestamp 1621261055
transform 1 0 3840 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_36
timestamp 1621261055
transform 1 0 4608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_521
timestamp 1621261055
transform 1 0 6432 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_44
timestamp 1621261055
transform 1 0 5376 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_52
timestamp 1621261055
transform 1 0 6144 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_54
timestamp 1621261055
transform 1 0 6336 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_56
timestamp 1621261055
transform 1 0 6528 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_64
timestamp 1621261055
transform 1 0 7296 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_72
timestamp 1621261055
transform 1 0 8064 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_80
timestamp 1621261055
transform 1 0 8832 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_88
timestamp 1621261055
transform 1 0 9600 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_96
timestamp 1621261055
transform 1 0 10368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_104
timestamp 1621261055
transform 1 0 11136 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_522
timestamp 1621261055
transform 1 0 11712 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_108
timestamp 1621261055
transform 1 0 11520 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_111
timestamp 1621261055
transform 1 0 11808 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_119
timestamp 1621261055
transform 1 0 12576 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_127
timestamp 1621261055
transform 1 0 13344 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_135
timestamp 1621261055
transform 1 0 14112 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_143
timestamp 1621261055
transform 1 0 14880 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_523
timestamp 1621261055
transform 1 0 16992 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_151
timestamp 1621261055
transform 1 0 15648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_159
timestamp 1621261055
transform 1 0 16416 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_163
timestamp 1621261055
transform 1 0 16800 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_166
timestamp 1621261055
transform 1 0 17088 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_174
timestamp 1621261055
transform 1 0 17856 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_182
timestamp 1621261055
transform 1 0 18624 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_190
timestamp 1621261055
transform 1 0 19392 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_198
timestamp 1621261055
transform 1 0 20160 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_206
timestamp 1621261055
transform 1 0 20928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_524
timestamp 1621261055
transform 1 0 22272 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_214
timestamp 1621261055
transform 1 0 21696 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_218
timestamp 1621261055
transform 1 0 22080 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_221
timestamp 1621261055
transform 1 0 22368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_229
timestamp 1621261055
transform 1 0 23136 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _095_
timestamp 1621261055
transform 1 0 25248 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_33_237
timestamp 1621261055
transform 1 0 23904 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_245
timestamp 1621261055
transform 1 0 24672 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_249
timestamp 1621261055
transform 1 0 25056 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_254
timestamp 1621261055
transform 1 0 25536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_262
timestamp 1621261055
transform 1 0 26304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_270
timestamp 1621261055
transform 1 0 27072 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_525
timestamp 1621261055
transform 1 0 27552 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_33_274
timestamp 1621261055
transform 1 0 27456 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_276
timestamp 1621261055
transform 1 0 27648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_284
timestamp 1621261055
transform 1 0 28416 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_292
timestamp 1621261055
transform 1 0 29184 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_300
timestamp 1621261055
transform 1 0 29952 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_308
timestamp 1621261055
transform 1 0 30720 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_526
timestamp 1621261055
transform 1 0 32832 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_316
timestamp 1621261055
transform 1 0 31488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_324
timestamp 1621261055
transform 1 0 32256 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_328
timestamp 1621261055
transform 1 0 32640 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_331
timestamp 1621261055
transform 1 0 32928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_339
timestamp 1621261055
transform 1 0 33696 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_347
timestamp 1621261055
transform 1 0 34464 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_355
timestamp 1621261055
transform 1 0 35232 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_363
timestamp 1621261055
transform 1 0 36000 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_371
timestamp 1621261055
transform 1 0 36768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_527
timestamp 1621261055
transform 1 0 38112 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_379
timestamp 1621261055
transform 1 0 37536 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_383
timestamp 1621261055
transform 1 0 37920 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_386
timestamp 1621261055
transform 1 0 38208 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_394
timestamp 1621261055
transform 1 0 38976 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_402
timestamp 1621261055
transform 1 0 39744 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_410
timestamp 1621261055
transform 1 0 40512 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_418
timestamp 1621261055
transform 1 0 41280 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_528
timestamp 1621261055
transform 1 0 43392 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_426
timestamp 1621261055
transform 1 0 42048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_434
timestamp 1621261055
transform 1 0 42816 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_438
timestamp 1621261055
transform 1 0 43200 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_441
timestamp 1621261055
transform 1 0 43488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_449
timestamp 1621261055
transform 1 0 44256 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_457
timestamp 1621261055
transform 1 0 45024 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _030_
timestamp 1621261055
transform -1 0 47232 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_19
timestamp 1621261055
transform -1 0 46944 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_465
timestamp 1621261055
transform 1 0 45792 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_473
timestamp 1621261055
transform 1 0 46560 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_480
timestamp 1621261055
transform 1 0 47232 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_529
timestamp 1621261055
transform 1 0 48672 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_488
timestamp 1621261055
transform 1 0 48000 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_492
timestamp 1621261055
transform 1 0 48384 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_494
timestamp 1621261055
transform 1 0 48576 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_496
timestamp 1621261055
transform 1 0 48768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_504
timestamp 1621261055
transform 1 0 49536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _194_
timestamp 1621261055
transform 1 0 50304 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_33_515
timestamp 1621261055
transform 1 0 50592 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_523
timestamp 1621261055
transform 1 0 51360 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_531
timestamp 1621261055
transform 1 0 52128 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_539
timestamp 1621261055
transform 1 0 52896 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _047_
timestamp 1621261055
transform -1 0 54720 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _108_
timestamp 1621261055
transform 1 0 55104 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_530
timestamp 1621261055
transform 1 0 53952 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_59
timestamp 1621261055
transform -1 0 54432 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_547
timestamp 1621261055
transform 1 0 53664 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_549
timestamp 1621261055
transform 1 0 53856 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_551
timestamp 1621261055
transform 1 0 54048 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_33_558
timestamp 1621261055
transform 1 0 54720 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_565
timestamp 1621261055
transform 1 0 55392 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_573
timestamp 1621261055
transform 1 0 56160 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_581
timestamp 1621261055
transform 1 0 56928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_67
timestamp 1621261055
transform -1 0 58848 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_589
timestamp 1621261055
transform 1 0 57696 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_68
timestamp 1621261055
transform 1 0 1152 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_4
timestamp 1621261055
transform 1 0 1536 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_12
timestamp 1621261055
transform 1 0 2304 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_20
timestamp 1621261055
transform 1 0 3072 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_531
timestamp 1621261055
transform 1 0 3840 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_29
timestamp 1621261055
transform 1 0 3936 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_37
timestamp 1621261055
transform 1 0 4704 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_45
timestamp 1621261055
transform 1 0 5472 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_53
timestamp 1621261055
transform 1 0 6240 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_61
timestamp 1621261055
transform 1 0 7008 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_532
timestamp 1621261055
transform 1 0 9120 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_69
timestamp 1621261055
transform 1 0 7776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_77
timestamp 1621261055
transform 1 0 8544 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_81
timestamp 1621261055
transform 1 0 8928 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_84
timestamp 1621261055
transform 1 0 9216 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_92
timestamp 1621261055
transform 1 0 9984 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_100
timestamp 1621261055
transform 1 0 10752 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_108
timestamp 1621261055
transform 1 0 11520 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_116
timestamp 1621261055
transform 1 0 12288 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_124
timestamp 1621261055
transform 1 0 13056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_533
timestamp 1621261055
transform 1 0 14400 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_132
timestamp 1621261055
transform 1 0 13824 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_136
timestamp 1621261055
transform 1 0 14208 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_139
timestamp 1621261055
transform 1 0 14496 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_147
timestamp 1621261055
transform 1 0 15264 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_155
timestamp 1621261055
transform 1 0 16032 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_163
timestamp 1621261055
transform 1 0 16800 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_171
timestamp 1621261055
transform 1 0 17568 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_179
timestamp 1621261055
transform 1 0 18336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_187
timestamp 1621261055
transform 1 0 19104 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_534
timestamp 1621261055
transform 1 0 19680 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_191
timestamp 1621261055
transform 1 0 19488 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_194
timestamp 1621261055
transform 1 0 19776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_202
timestamp 1621261055
transform 1 0 20544 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_210
timestamp 1621261055
transform 1 0 21312 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_218
timestamp 1621261055
transform 1 0 22080 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_226
timestamp 1621261055
transform 1 0 22848 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_535
timestamp 1621261055
transform 1 0 24960 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_234
timestamp 1621261055
transform 1 0 23616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_242
timestamp 1621261055
transform 1 0 24384 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_246
timestamp 1621261055
transform 1 0 24768 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_249
timestamp 1621261055
transform 1 0 25056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_257
timestamp 1621261055
transform 1 0 25824 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_265
timestamp 1621261055
transform 1 0 26592 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_273
timestamp 1621261055
transform 1 0 27360 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_281
timestamp 1621261055
transform 1 0 28128 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_289
timestamp 1621261055
transform 1 0 28896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_536
timestamp 1621261055
transform 1 0 30240 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_297
timestamp 1621261055
transform 1 0 29664 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_301
timestamp 1621261055
transform 1 0 30048 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_304
timestamp 1621261055
transform 1 0 30336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_312
timestamp 1621261055
transform 1 0 31104 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_320
timestamp 1621261055
transform 1 0 31872 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_328
timestamp 1621261055
transform 1 0 32640 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_336
timestamp 1621261055
transform 1 0 33408 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_344
timestamp 1621261055
transform 1 0 34176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_352
timestamp 1621261055
transform 1 0 34944 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_356
timestamp 1621261055
transform 1 0 35328 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_537
timestamp 1621261055
transform 1 0 35520 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_359
timestamp 1621261055
transform 1 0 35616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_367
timestamp 1621261055
transform 1 0 36384 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_375
timestamp 1621261055
transform 1 0 37152 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_383
timestamp 1621261055
transform 1 0 37920 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_391
timestamp 1621261055
transform 1 0 38688 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_399
timestamp 1621261055
transform 1 0 39456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_538
timestamp 1621261055
transform 1 0 40800 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_407
timestamp 1621261055
transform 1 0 40224 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_411
timestamp 1621261055
transform 1 0 40608 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_414
timestamp 1621261055
transform 1 0 40896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_422
timestamp 1621261055
transform 1 0 41664 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_430
timestamp 1621261055
transform 1 0 42432 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_438
timestamp 1621261055
transform 1 0 43200 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_446
timestamp 1621261055
transform 1 0 43968 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_454
timestamp 1621261055
transform 1 0 44736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_462
timestamp 1621261055
transform 1 0 45504 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_539
timestamp 1621261055
transform 1 0 46080 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_466
timestamp 1621261055
transform 1 0 45888 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_469
timestamp 1621261055
transform 1 0 46176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_477
timestamp 1621261055
transform 1 0 46944 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_485
timestamp 1621261055
transform 1 0 47712 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_493
timestamp 1621261055
transform 1 0 48480 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_501
timestamp 1621261055
transform 1 0 49248 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_540
timestamp 1621261055
transform 1 0 51360 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_509
timestamp 1621261055
transform 1 0 50016 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_517
timestamp 1621261055
transform 1 0 50784 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_521
timestamp 1621261055
transform 1 0 51168 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_524
timestamp 1621261055
transform 1 0 51456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_532
timestamp 1621261055
transform 1 0 52224 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_540
timestamp 1621261055
transform 1 0 52992 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_548
timestamp 1621261055
transform 1 0 53760 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_556
timestamp 1621261055
transform 1 0 54528 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_564
timestamp 1621261055
transform 1 0 55296 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _114_
timestamp 1621261055
transform 1 0 57120 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_541
timestamp 1621261055
transform 1 0 56640 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_572
timestamp 1621261055
transform 1 0 56064 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_576
timestamp 1621261055
transform 1 0 56448 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_34_579
timestamp 1621261055
transform 1 0 56736 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_586
timestamp 1621261055
transform 1 0 57408 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_69
timestamp 1621261055
transform -1 0 58848 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_594
timestamp 1621261055
transform 1 0 58176 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_34_596
timestamp 1621261055
transform 1 0 58368 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_70
timestamp 1621261055
transform 1 0 1152 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_4
timestamp 1621261055
transform 1 0 1536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_12
timestamp 1621261055
transform 1 0 2304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_20
timestamp 1621261055
transform 1 0 3072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_28
timestamp 1621261055
transform 1 0 3840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_36
timestamp 1621261055
transform 1 0 4608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_542
timestamp 1621261055
transform 1 0 6432 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_44
timestamp 1621261055
transform 1 0 5376 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_52
timestamp 1621261055
transform 1 0 6144 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_35_54
timestamp 1621261055
transform 1 0 6336 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_56
timestamp 1621261055
transform 1 0 6528 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_64
timestamp 1621261055
transform 1 0 7296 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_72
timestamp 1621261055
transform 1 0 8064 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_80
timestamp 1621261055
transform 1 0 8832 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_88
timestamp 1621261055
transform 1 0 9600 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_96
timestamp 1621261055
transform 1 0 10368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_104
timestamp 1621261055
transform 1 0 11136 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_543
timestamp 1621261055
transform 1 0 11712 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_108
timestamp 1621261055
transform 1 0 11520 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_111
timestamp 1621261055
transform 1 0 11808 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_119
timestamp 1621261055
transform 1 0 12576 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_127
timestamp 1621261055
transform 1 0 13344 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_135
timestamp 1621261055
transform 1 0 14112 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_143
timestamp 1621261055
transform 1 0 14880 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_544
timestamp 1621261055
transform 1 0 16992 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_151
timestamp 1621261055
transform 1 0 15648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_159
timestamp 1621261055
transform 1 0 16416 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_163
timestamp 1621261055
transform 1 0 16800 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_166
timestamp 1621261055
transform 1 0 17088 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_174
timestamp 1621261055
transform 1 0 17856 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_182
timestamp 1621261055
transform 1 0 18624 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_190
timestamp 1621261055
transform 1 0 19392 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_198
timestamp 1621261055
transform 1 0 20160 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_206
timestamp 1621261055
transform 1 0 20928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_545
timestamp 1621261055
transform 1 0 22272 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_214
timestamp 1621261055
transform 1 0 21696 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_218
timestamp 1621261055
transform 1 0 22080 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_221
timestamp 1621261055
transform 1 0 22368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_229
timestamp 1621261055
transform 1 0 23136 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_237
timestamp 1621261055
transform 1 0 23904 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_245
timestamp 1621261055
transform 1 0 24672 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_253
timestamp 1621261055
transform 1 0 25440 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_261
timestamp 1621261055
transform 1 0 26208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_269
timestamp 1621261055
transform 1 0 26976 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_273
timestamp 1621261055
transform 1 0 27360 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_546
timestamp 1621261055
transform 1 0 27552 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_276
timestamp 1621261055
transform 1 0 27648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_284
timestamp 1621261055
transform 1 0 28416 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_292
timestamp 1621261055
transform 1 0 29184 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_300
timestamp 1621261055
transform 1 0 29952 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_308
timestamp 1621261055
transform 1 0 30720 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_547
timestamp 1621261055
transform 1 0 32832 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_316
timestamp 1621261055
transform 1 0 31488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_324
timestamp 1621261055
transform 1 0 32256 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_328
timestamp 1621261055
transform 1 0 32640 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_331
timestamp 1621261055
transform 1 0 32928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_339
timestamp 1621261055
transform 1 0 33696 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_347
timestamp 1621261055
transform 1 0 34464 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_355
timestamp 1621261055
transform 1 0 35232 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_363
timestamp 1621261055
transform 1 0 36000 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_371
timestamp 1621261055
transform 1 0 36768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_548
timestamp 1621261055
transform 1 0 38112 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_379
timestamp 1621261055
transform 1 0 37536 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_383
timestamp 1621261055
transform 1 0 37920 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_386
timestamp 1621261055
transform 1 0 38208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_394
timestamp 1621261055
transform 1 0 38976 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_402
timestamp 1621261055
transform 1 0 39744 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_410
timestamp 1621261055
transform 1 0 40512 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_418
timestamp 1621261055
transform 1 0 41280 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_549
timestamp 1621261055
transform 1 0 43392 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_426
timestamp 1621261055
transform 1 0 42048 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_434
timestamp 1621261055
transform 1 0 42816 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_438
timestamp 1621261055
transform 1 0 43200 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_441
timestamp 1621261055
transform 1 0 43488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_449
timestamp 1621261055
transform 1 0 44256 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_457
timestamp 1621261055
transform 1 0 45024 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_465
timestamp 1621261055
transform 1 0 45792 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_473
timestamp 1621261055
transform 1 0 46560 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_481
timestamp 1621261055
transform 1 0 47328 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_550
timestamp 1621261055
transform 1 0 48672 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_489
timestamp 1621261055
transform 1 0 48096 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_493
timestamp 1621261055
transform 1 0 48480 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_496
timestamp 1621261055
transform 1 0 48768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_504
timestamp 1621261055
transform 1 0 49536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_512
timestamp 1621261055
transform 1 0 50304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_520
timestamp 1621261055
transform 1 0 51072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_528
timestamp 1621261055
transform 1 0 51840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_536
timestamp 1621261055
transform 1 0 52608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_544
timestamp 1621261055
transform 1 0 53376 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_551
timestamp 1621261055
transform 1 0 53952 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_548
timestamp 1621261055
transform 1 0 53760 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_551
timestamp 1621261055
transform 1 0 54048 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_559
timestamp 1621261055
transform 1 0 54816 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_567
timestamp 1621261055
transform 1 0 55584 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_575
timestamp 1621261055
transform 1 0 56352 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_583
timestamp 1621261055
transform 1 0 57120 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_71
timestamp 1621261055
transform -1 0 58848 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_35_591
timestamp 1621261055
transform 1 0 57888 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_595
timestamp 1621261055
transform 1 0 58272 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_72
timestamp 1621261055
transform 1 0 1152 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_4
timestamp 1621261055
transform 1 0 1536 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_12
timestamp 1621261055
transform 1 0 2304 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_20
timestamp 1621261055
transform 1 0 3072 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_552
timestamp 1621261055
transform 1 0 3840 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_29
timestamp 1621261055
transform 1 0 3936 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_37
timestamp 1621261055
transform 1 0 4704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_45
timestamp 1621261055
transform 1 0 5472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_53
timestamp 1621261055
transform 1 0 6240 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_61
timestamp 1621261055
transform 1 0 7008 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_553
timestamp 1621261055
transform 1 0 9120 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_69
timestamp 1621261055
transform 1 0 7776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_77
timestamp 1621261055
transform 1 0 8544 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_81
timestamp 1621261055
transform 1 0 8928 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_84
timestamp 1621261055
transform 1 0 9216 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_92
timestamp 1621261055
transform 1 0 9984 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_100
timestamp 1621261055
transform 1 0 10752 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_108
timestamp 1621261055
transform 1 0 11520 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_116
timestamp 1621261055
transform 1 0 12288 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_124
timestamp 1621261055
transform 1 0 13056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _208_
timestamp 1621261055
transform 1 0 14880 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_554
timestamp 1621261055
transform 1 0 14400 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_132
timestamp 1621261055
transform 1 0 13824 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_136
timestamp 1621261055
transform 1 0 14208 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_36_139
timestamp 1621261055
transform 1 0 14496 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_146
timestamp 1621261055
transform 1 0 15168 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _064_
timestamp 1621261055
transform 1 0 16416 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_36_154
timestamp 1621261055
transform 1 0 15936 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_36_158
timestamp 1621261055
transform 1 0 16320 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_162
timestamp 1621261055
transform 1 0 16704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _036_
timestamp 1621261055
transform -1 0 19200 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_95
timestamp 1621261055
transform -1 0 18912 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_170
timestamp 1621261055
transform 1 0 17472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_178
timestamp 1621261055
transform 1 0 18240 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_36_182
timestamp 1621261055
transform 1 0 18624 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_188
timestamp 1621261055
transform 1 0 19200 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_555
timestamp 1621261055
transform 1 0 19680 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_36_192
timestamp 1621261055
transform 1 0 19584 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_194
timestamp 1621261055
transform 1 0 19776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_202
timestamp 1621261055
transform 1 0 20544 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_210
timestamp 1621261055
transform 1 0 21312 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_218
timestamp 1621261055
transform 1 0 22080 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_226
timestamp 1621261055
transform 1 0 22848 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_556
timestamp 1621261055
transform 1 0 24960 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_234
timestamp 1621261055
transform 1 0 23616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_242
timestamp 1621261055
transform 1 0 24384 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_246
timestamp 1621261055
transform 1 0 24768 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_249
timestamp 1621261055
transform 1 0 25056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_257
timestamp 1621261055
transform 1 0 25824 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_265
timestamp 1621261055
transform 1 0 26592 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_273
timestamp 1621261055
transform 1 0 27360 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_281
timestamp 1621261055
transform 1 0 28128 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_289
timestamp 1621261055
transform 1 0 28896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_557
timestamp 1621261055
transform 1 0 30240 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_297
timestamp 1621261055
transform 1 0 29664 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_301
timestamp 1621261055
transform 1 0 30048 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_304
timestamp 1621261055
transform 1 0 30336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_312
timestamp 1621261055
transform 1 0 31104 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_320
timestamp 1621261055
transform 1 0 31872 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_328
timestamp 1621261055
transform 1 0 32640 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_336
timestamp 1621261055
transform 1 0 33408 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_344
timestamp 1621261055
transform 1 0 34176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_352
timestamp 1621261055
transform 1 0 34944 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_356
timestamp 1621261055
transform 1 0 35328 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_558
timestamp 1621261055
transform 1 0 35520 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_359
timestamp 1621261055
transform 1 0 35616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_367
timestamp 1621261055
transform 1 0 36384 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_375
timestamp 1621261055
transform 1 0 37152 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_383
timestamp 1621261055
transform 1 0 37920 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_391
timestamp 1621261055
transform 1 0 38688 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_399
timestamp 1621261055
transform 1 0 39456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_559
timestamp 1621261055
transform 1 0 40800 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_407
timestamp 1621261055
transform 1 0 40224 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_411
timestamp 1621261055
transform 1 0 40608 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_414
timestamp 1621261055
transform 1 0 40896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_422
timestamp 1621261055
transform 1 0 41664 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_430
timestamp 1621261055
transform 1 0 42432 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_438
timestamp 1621261055
transform 1 0 43200 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_446
timestamp 1621261055
transform 1 0 43968 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_454
timestamp 1621261055
transform 1 0 44736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_462
timestamp 1621261055
transform 1 0 45504 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_560
timestamp 1621261055
transform 1 0 46080 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_466
timestamp 1621261055
transform 1 0 45888 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_469
timestamp 1621261055
transform 1 0 46176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_477
timestamp 1621261055
transform 1 0 46944 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_485
timestamp 1621261055
transform 1 0 47712 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_493
timestamp 1621261055
transform 1 0 48480 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_501
timestamp 1621261055
transform 1 0 49248 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_561
timestamp 1621261055
transform 1 0 51360 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_509
timestamp 1621261055
transform 1 0 50016 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_517
timestamp 1621261055
transform 1 0 50784 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_521
timestamp 1621261055
transform 1 0 51168 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_524
timestamp 1621261055
transform 1 0 51456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_532
timestamp 1621261055
transform 1 0 52224 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_540
timestamp 1621261055
transform 1 0 52992 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_548
timestamp 1621261055
transform 1 0 53760 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_556
timestamp 1621261055
transform 1 0 54528 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_564
timestamp 1621261055
transform 1 0 55296 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_562
timestamp 1621261055
transform 1 0 56640 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_572
timestamp 1621261055
transform 1 0 56064 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_576
timestamp 1621261055
transform 1 0 56448 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_579
timestamp 1621261055
transform 1 0 56736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_587
timestamp 1621261055
transform 1 0 57504 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_73
timestamp 1621261055
transform -1 0 58848 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_595
timestamp 1621261055
transform 1 0 58272 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_74
timestamp 1621261055
transform 1 0 1152 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_4
timestamp 1621261055
transform 1 0 1536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_12
timestamp 1621261055
transform 1 0 2304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_20
timestamp 1621261055
transform 1 0 3072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_28
timestamp 1621261055
transform 1 0 3840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_36
timestamp 1621261055
transform 1 0 4608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_563
timestamp 1621261055
transform 1 0 6432 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_44
timestamp 1621261055
transform 1 0 5376 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_52
timestamp 1621261055
transform 1 0 6144 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_54
timestamp 1621261055
transform 1 0 6336 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_56
timestamp 1621261055
transform 1 0 6528 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_64
timestamp 1621261055
transform 1 0 7296 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_72
timestamp 1621261055
transform 1 0 8064 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_80
timestamp 1621261055
transform 1 0 8832 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_88
timestamp 1621261055
transform 1 0 9600 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_96
timestamp 1621261055
transform 1 0 10368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_104
timestamp 1621261055
transform 1 0 11136 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_564
timestamp 1621261055
transform 1 0 11712 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_108
timestamp 1621261055
transform 1 0 11520 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_111
timestamp 1621261055
transform 1 0 11808 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_119
timestamp 1621261055
transform 1 0 12576 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_127
timestamp 1621261055
transform 1 0 13344 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_135
timestamp 1621261055
transform 1 0 14112 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_143
timestamp 1621261055
transform 1 0 14880 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_565
timestamp 1621261055
transform 1 0 16992 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_151
timestamp 1621261055
transform 1 0 15648 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_159
timestamp 1621261055
transform 1 0 16416 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_163
timestamp 1621261055
transform 1 0 16800 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_166
timestamp 1621261055
transform 1 0 17088 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _120_
timestamp 1621261055
transform 1 0 18048 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_174
timestamp 1621261055
transform 1 0 17856 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_179
timestamp 1621261055
transform 1 0 18336 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_187
timestamp 1621261055
transform 1 0 19104 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_195
timestamp 1621261055
transform 1 0 19872 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_203
timestamp 1621261055
transform 1 0 20640 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_566
timestamp 1621261055
transform 1 0 22272 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_211
timestamp 1621261055
transform 1 0 21408 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_37_219
timestamp 1621261055
transform 1 0 22176 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_221
timestamp 1621261055
transform 1 0 22368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_229
timestamp 1621261055
transform 1 0 23136 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _043_
timestamp 1621261055
transform -1 0 24576 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_47
timestamp 1621261055
transform -1 0 24288 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_237
timestamp 1621261055
transform 1 0 23904 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_244
timestamp 1621261055
transform 1 0 24576 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_252
timestamp 1621261055
transform 1 0 25344 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_260
timestamp 1621261055
transform 1 0 26112 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_268
timestamp 1621261055
transform 1 0 26880 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_272
timestamp 1621261055
transform 1 0 27264 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _023_
timestamp 1621261055
transform 1 0 28032 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_567
timestamp 1621261055
transform 1 0 27552 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_35
timestamp 1621261055
transform 1 0 27840 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_274
timestamp 1621261055
transform 1 0 27456 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_276
timestamp 1621261055
transform 1 0 27648 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_283
timestamp 1621261055
transform 1 0 28320 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_291
timestamp 1621261055
transform 1 0 29088 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_299
timestamp 1621261055
transform 1 0 29856 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_307
timestamp 1621261055
transform 1 0 30624 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_315
timestamp 1621261055
transform 1 0 31392 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_568
timestamp 1621261055
transform 1 0 32832 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_323
timestamp 1621261055
transform 1 0 32160 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_327
timestamp 1621261055
transform 1 0 32544 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_329
timestamp 1621261055
transform 1 0 32736 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_331
timestamp 1621261055
transform 1 0 32928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_339
timestamp 1621261055
transform 1 0 33696 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_347
timestamp 1621261055
transform 1 0 34464 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_355
timestamp 1621261055
transform 1 0 35232 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_363
timestamp 1621261055
transform 1 0 36000 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_371
timestamp 1621261055
transform 1 0 36768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_569
timestamp 1621261055
transform 1 0 38112 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_379
timestamp 1621261055
transform 1 0 37536 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_383
timestamp 1621261055
transform 1 0 37920 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_386
timestamp 1621261055
transform 1 0 38208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_394
timestamp 1621261055
transform 1 0 38976 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_402
timestamp 1621261055
transform 1 0 39744 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_410
timestamp 1621261055
transform 1 0 40512 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_418
timestamp 1621261055
transform 1 0 41280 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_570
timestamp 1621261055
transform 1 0 43392 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_426
timestamp 1621261055
transform 1 0 42048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_434
timestamp 1621261055
transform 1 0 42816 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_438
timestamp 1621261055
transform 1 0 43200 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_441
timestamp 1621261055
transform 1 0 43488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_449
timestamp 1621261055
transform 1 0 44256 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_457
timestamp 1621261055
transform 1 0 45024 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_465
timestamp 1621261055
transform 1 0 45792 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_473
timestamp 1621261055
transform 1 0 46560 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_481
timestamp 1621261055
transform 1 0 47328 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_571
timestamp 1621261055
transform 1 0 48672 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_489
timestamp 1621261055
transform 1 0 48096 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_493
timestamp 1621261055
transform 1 0 48480 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_496
timestamp 1621261055
transform 1 0 48768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_504
timestamp 1621261055
transform 1 0 49536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_512
timestamp 1621261055
transform 1 0 50304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_520
timestamp 1621261055
transform 1 0 51072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_528
timestamp 1621261055
transform 1 0 51840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_536
timestamp 1621261055
transform 1 0 52608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_544
timestamp 1621261055
transform 1 0 53376 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_572
timestamp 1621261055
transform 1 0 53952 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_548
timestamp 1621261055
transform 1 0 53760 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_551
timestamp 1621261055
transform 1 0 54048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_559
timestamp 1621261055
transform 1 0 54816 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_567
timestamp 1621261055
transform 1 0 55584 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _138_
timestamp 1621261055
transform 1 0 56832 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _183_
timestamp 1621261055
transform 1 0 56160 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_571
timestamp 1621261055
transform 1 0 55968 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_37_576
timestamp 1621261055
transform 1 0 56448 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_583
timestamp 1621261055
transform 1 0 57120 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_75
timestamp 1621261055
transform -1 0 58848 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_37_591
timestamp 1621261055
transform 1 0 57888 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_595
timestamp 1621261055
transform 1 0 58272 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_76
timestamp 1621261055
transform 1 0 1152 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_78
timestamp 1621261055
transform 1 0 1152 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_4
timestamp 1621261055
transform 1 0 1536 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_12
timestamp 1621261055
transform 1 0 2304 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_20
timestamp 1621261055
transform 1 0 3072 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_4
timestamp 1621261055
transform 1 0 1536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_12
timestamp 1621261055
transform 1 0 2304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_20
timestamp 1621261055
transform 1 0 3072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_573
timestamp 1621261055
transform 1 0 3840 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_29
timestamp 1621261055
transform 1 0 3936 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_37
timestamp 1621261055
transform 1 0 4704 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_28
timestamp 1621261055
transform 1 0 3840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_36
timestamp 1621261055
transform 1 0 4608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_584
timestamp 1621261055
transform 1 0 6432 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_45
timestamp 1621261055
transform 1 0 5472 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_53
timestamp 1621261055
transform 1 0 6240 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_61
timestamp 1621261055
transform 1 0 7008 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_44
timestamp 1621261055
transform 1 0 5376 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_52
timestamp 1621261055
transform 1 0 6144 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_39_54
timestamp 1621261055
transform 1 0 6336 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_56
timestamp 1621261055
transform 1 0 6528 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_574
timestamp 1621261055
transform 1 0 9120 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_69
timestamp 1621261055
transform 1 0 7776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_77
timestamp 1621261055
transform 1 0 8544 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_81
timestamp 1621261055
transform 1 0 8928 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_84
timestamp 1621261055
transform 1 0 9216 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_64
timestamp 1621261055
transform 1 0 7296 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_72
timestamp 1621261055
transform 1 0 8064 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_80
timestamp 1621261055
transform 1 0 8832 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _035_
timestamp 1621261055
transform -1 0 11424 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_57
timestamp 1621261055
transform -1 0 11136 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_92
timestamp 1621261055
transform 1 0 9984 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_100
timestamp 1621261055
transform 1 0 10752 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_88
timestamp 1621261055
transform 1 0 9600 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_96
timestamp 1621261055
transform 1 0 10368 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_104
timestamp 1621261055
transform 1 0 11136 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_585
timestamp 1621261055
transform 1 0 11712 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_107
timestamp 1621261055
transform 1 0 11424 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_115
timestamp 1621261055
transform 1 0 12192 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_123
timestamp 1621261055
transform 1 0 12960 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_108
timestamp 1621261055
transform 1 0 11520 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_111
timestamp 1621261055
transform 1 0 11808 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_119
timestamp 1621261055
transform 1 0 12576 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_575
timestamp 1621261055
transform 1 0 14400 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_131
timestamp 1621261055
transform 1 0 13728 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_135
timestamp 1621261055
transform 1 0 14112 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_38_137
timestamp 1621261055
transform 1 0 14304 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_139
timestamp 1621261055
transform 1 0 14496 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_147
timestamp 1621261055
transform 1 0 15264 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_127
timestamp 1621261055
transform 1 0 13344 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_135
timestamp 1621261055
transform 1 0 14112 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_143
timestamp 1621261055
transform 1 0 14880 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_586
timestamp 1621261055
transform 1 0 16992 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_155
timestamp 1621261055
transform 1 0 16032 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_163
timestamp 1621261055
transform 1 0 16800 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_151
timestamp 1621261055
transform 1 0 15648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_159
timestamp 1621261055
transform 1 0 16416 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_163
timestamp 1621261055
transform 1 0 16800 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_166
timestamp 1621261055
transform 1 0 17088 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _203_
timestamp 1621261055
transform 1 0 18240 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_38_171
timestamp 1621261055
transform 1 0 17568 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_179
timestamp 1621261055
transform 1 0 18336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_187
timestamp 1621261055
transform 1 0 19104 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_39_174
timestamp 1621261055
transform 1 0 17856 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_181
timestamp 1621261055
transform 1 0 18528 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_189
timestamp 1621261055
transform 1 0 19296 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_576
timestamp 1621261055
transform 1 0 19680 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_191
timestamp 1621261055
transform 1 0 19488 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_194
timestamp 1621261055
transform 1 0 19776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_202
timestamp 1621261055
transform 1 0 20544 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_210
timestamp 1621261055
transform 1 0 21312 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_197
timestamp 1621261055
transform 1 0 20064 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_205
timestamp 1621261055
transform 1 0 20832 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_587
timestamp 1621261055
transform 1 0 22272 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_218
timestamp 1621261055
transform 1 0 22080 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_226
timestamp 1621261055
transform 1 0 22848 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_213
timestamp 1621261055
transform 1 0 21600 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_217
timestamp 1621261055
transform 1 0 21984 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_39_219
timestamp 1621261055
transform 1 0 22176 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_221
timestamp 1621261055
transform 1 0 22368 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_229
timestamp 1621261055
transform 1 0 23136 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_577
timestamp 1621261055
transform 1 0 24960 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_234
timestamp 1621261055
transform 1 0 23616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_242
timestamp 1621261055
transform 1 0 24384 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_246
timestamp 1621261055
transform 1 0 24768 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_249
timestamp 1621261055
transform 1 0 25056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_237
timestamp 1621261055
transform 1 0 23904 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_245
timestamp 1621261055
transform 1 0 24672 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_257
timestamp 1621261055
transform 1 0 25824 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_265
timestamp 1621261055
transform 1 0 26592 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_273
timestamp 1621261055
transform 1 0 27360 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_253
timestamp 1621261055
transform 1 0 25440 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_261
timestamp 1621261055
transform 1 0 26208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_269
timestamp 1621261055
transform 1 0 26976 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_273
timestamp 1621261055
transform 1 0 27360 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_588
timestamp 1621261055
transform 1 0 27552 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_281
timestamp 1621261055
transform 1 0 28128 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_289
timestamp 1621261055
transform 1 0 28896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_276
timestamp 1621261055
transform 1 0 27648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_284
timestamp 1621261055
transform 1 0 28416 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_292
timestamp 1621261055
transform 1 0 29184 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_578
timestamp 1621261055
transform 1 0 30240 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_297
timestamp 1621261055
transform 1 0 29664 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_301
timestamp 1621261055
transform 1 0 30048 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_304
timestamp 1621261055
transform 1 0 30336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_312
timestamp 1621261055
transform 1 0 31104 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_300
timestamp 1621261055
transform 1 0 29952 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_308
timestamp 1621261055
transform 1 0 30720 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_589
timestamp 1621261055
transform 1 0 32832 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_320
timestamp 1621261055
transform 1 0 31872 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_328
timestamp 1621261055
transform 1 0 32640 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_336
timestamp 1621261055
transform 1 0 33408 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_316
timestamp 1621261055
transform 1 0 31488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_324
timestamp 1621261055
transform 1 0 32256 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_328
timestamp 1621261055
transform 1 0 32640 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_331
timestamp 1621261055
transform 1 0 32928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_344
timestamp 1621261055
transform 1 0 34176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_352
timestamp 1621261055
transform 1 0 34944 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_356
timestamp 1621261055
transform 1 0 35328 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_339
timestamp 1621261055
transform 1 0 33696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_347
timestamp 1621261055
transform 1 0 34464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_355
timestamp 1621261055
transform 1 0 35232 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _137_
timestamp 1621261055
transform 1 0 37344 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _145_
timestamp 1621261055
transform 1 0 36000 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_579
timestamp 1621261055
transform 1 0 35520 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_359
timestamp 1621261055
transform 1 0 35616 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_366
timestamp 1621261055
transform 1 0 36288 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_374
timestamp 1621261055
transform 1 0 37056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_363
timestamp 1621261055
transform 1 0 36000 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_371
timestamp 1621261055
transform 1 0 36768 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_375
timestamp 1621261055
transform 1 0 37152 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_590
timestamp 1621261055
transform 1 0 38112 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_382
timestamp 1621261055
transform 1 0 37824 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_390
timestamp 1621261055
transform 1 0 38592 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_398
timestamp 1621261055
transform 1 0 39360 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_380
timestamp 1621261055
transform 1 0 37632 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_39_384
timestamp 1621261055
transform 1 0 38016 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_386
timestamp 1621261055
transform 1 0 38208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_394
timestamp 1621261055
transform 1 0 38976 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_580
timestamp 1621261055
transform 1 0 40800 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_406
timestamp 1621261055
transform 1 0 40128 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_410
timestamp 1621261055
transform 1 0 40512 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_38_412
timestamp 1621261055
transform 1 0 40704 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_414
timestamp 1621261055
transform 1 0 40896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_402
timestamp 1621261055
transform 1 0 39744 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_410
timestamp 1621261055
transform 1 0 40512 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_418
timestamp 1621261055
transform 1 0 41280 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_591
timestamp 1621261055
transform 1 0 43392 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_422
timestamp 1621261055
transform 1 0 41664 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_430
timestamp 1621261055
transform 1 0 42432 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_438
timestamp 1621261055
transform 1 0 43200 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_426
timestamp 1621261055
transform 1 0 42048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_434
timestamp 1621261055
transform 1 0 42816 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_438
timestamp 1621261055
transform 1 0 43200 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_441
timestamp 1621261055
transform 1 0 43488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_446
timestamp 1621261055
transform 1 0 43968 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_454
timestamp 1621261055
transform 1 0 44736 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_462
timestamp 1621261055
transform 1 0 45504 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_449
timestamp 1621261055
transform 1 0 44256 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_457
timestamp 1621261055
transform 1 0 45024 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_581
timestamp 1621261055
transform 1 0 46080 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_466
timestamp 1621261055
transform 1 0 45888 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_469
timestamp 1621261055
transform 1 0 46176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_477
timestamp 1621261055
transform 1 0 46944 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_465
timestamp 1621261055
transform 1 0 45792 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_473
timestamp 1621261055
transform 1 0 46560 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_481
timestamp 1621261055
transform 1 0 47328 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_592
timestamp 1621261055
transform 1 0 48672 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_485
timestamp 1621261055
transform 1 0 47712 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_493
timestamp 1621261055
transform 1 0 48480 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_501
timestamp 1621261055
transform 1 0 49248 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_489
timestamp 1621261055
transform 1 0 48096 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_493
timestamp 1621261055
transform 1 0 48480 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_496
timestamp 1621261055
transform 1 0 48768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_504
timestamp 1621261055
transform 1 0 49536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_582
timestamp 1621261055
transform 1 0 51360 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_509
timestamp 1621261055
transform 1 0 50016 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_517
timestamp 1621261055
transform 1 0 50784 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_521
timestamp 1621261055
transform 1 0 51168 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_524
timestamp 1621261055
transform 1 0 51456 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_512
timestamp 1621261055
transform 1 0 50304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_520
timestamp 1621261055
transform 1 0 51072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_532
timestamp 1621261055
transform 1 0 52224 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_540
timestamp 1621261055
transform 1 0 52992 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_528
timestamp 1621261055
transform 1 0 51840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_536
timestamp 1621261055
transform 1 0 52608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_544
timestamp 1621261055
transform 1 0 53376 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_593
timestamp 1621261055
transform 1 0 53952 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_548
timestamp 1621261055
transform 1 0 53760 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_556
timestamp 1621261055
transform 1 0 54528 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_564
timestamp 1621261055
transform 1 0 55296 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_548
timestamp 1621261055
transform 1 0 53760 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_551
timestamp 1621261055
transform 1 0 54048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_559
timestamp 1621261055
transform 1 0 54816 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_567
timestamp 1621261055
transform 1 0 55584 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_583
timestamp 1621261055
transform 1 0 56640 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_572
timestamp 1621261055
transform 1 0 56064 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_576
timestamp 1621261055
transform 1 0 56448 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_579
timestamp 1621261055
transform 1 0 56736 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_587
timestamp 1621261055
transform 1 0 57504 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_575
timestamp 1621261055
transform 1 0 56352 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_583
timestamp 1621261055
transform 1 0 57120 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_77
timestamp 1621261055
transform -1 0 58848 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_79
timestamp 1621261055
transform -1 0 58848 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_595
timestamp 1621261055
transform 1 0 58272 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_591
timestamp 1621261055
transform 1 0 57888 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_595
timestamp 1621261055
transform 1 0 58272 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_80
timestamp 1621261055
transform 1 0 1152 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_40_4
timestamp 1621261055
transform 1 0 1536 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_12
timestamp 1621261055
transform 1 0 2304 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_20
timestamp 1621261055
transform 1 0 3072 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_594
timestamp 1621261055
transform 1 0 3840 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_29
timestamp 1621261055
transform 1 0 3936 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_37
timestamp 1621261055
transform 1 0 4704 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _060_
timestamp 1621261055
transform 1 0 6048 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_40_45
timestamp 1621261055
transform 1 0 5472 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_49
timestamp 1621261055
transform 1 0 5856 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_54
timestamp 1621261055
transform 1 0 6336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_62
timestamp 1621261055
transform 1 0 7104 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_595
timestamp 1621261055
transform 1 0 9120 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_70
timestamp 1621261055
transform 1 0 7872 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_78
timestamp 1621261055
transform 1 0 8640 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_40_82
timestamp 1621261055
transform 1 0 9024 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_84
timestamp 1621261055
transform 1 0 9216 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_92
timestamp 1621261055
transform 1 0 9984 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_100
timestamp 1621261055
transform 1 0 10752 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_108
timestamp 1621261055
transform 1 0 11520 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_116
timestamp 1621261055
transform 1 0 12288 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_124
timestamp 1621261055
transform 1 0 13056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_596
timestamp 1621261055
transform 1 0 14400 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_132
timestamp 1621261055
transform 1 0 13824 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_136
timestamp 1621261055
transform 1 0 14208 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_139
timestamp 1621261055
transform 1 0 14496 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_147
timestamp 1621261055
transform 1 0 15264 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_155
timestamp 1621261055
transform 1 0 16032 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_163
timestamp 1621261055
transform 1 0 16800 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_171
timestamp 1621261055
transform 1 0 17568 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_179
timestamp 1621261055
transform 1 0 18336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_187
timestamp 1621261055
transform 1 0 19104 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_597
timestamp 1621261055
transform 1 0 19680 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_191
timestamp 1621261055
transform 1 0 19488 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_194
timestamp 1621261055
transform 1 0 19776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_202
timestamp 1621261055
transform 1 0 20544 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_210
timestamp 1621261055
transform 1 0 21312 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_218
timestamp 1621261055
transform 1 0 22080 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_226
timestamp 1621261055
transform 1 0 22848 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_598
timestamp 1621261055
transform 1 0 24960 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_234
timestamp 1621261055
transform 1 0 23616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_242
timestamp 1621261055
transform 1 0 24384 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_246
timestamp 1621261055
transform 1 0 24768 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_249
timestamp 1621261055
transform 1 0 25056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_257
timestamp 1621261055
transform 1 0 25824 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_265
timestamp 1621261055
transform 1 0 26592 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_273
timestamp 1621261055
transform 1 0 27360 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_281
timestamp 1621261055
transform 1 0 28128 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_289
timestamp 1621261055
transform 1 0 28896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_599
timestamp 1621261055
transform 1 0 30240 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_297
timestamp 1621261055
transform 1 0 29664 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_301
timestamp 1621261055
transform 1 0 30048 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_304
timestamp 1621261055
transform 1 0 30336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_312
timestamp 1621261055
transform 1 0 31104 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_320
timestamp 1621261055
transform 1 0 31872 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_328
timestamp 1621261055
transform 1 0 32640 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_336
timestamp 1621261055
transform 1 0 33408 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_344
timestamp 1621261055
transform 1 0 34176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_352
timestamp 1621261055
transform 1 0 34944 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_356
timestamp 1621261055
transform 1 0 35328 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _152_
timestamp 1621261055
transform 1 0 36192 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _154_
timestamp 1621261055
transform 1 0 36864 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_600
timestamp 1621261055
transform 1 0 35520 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_359
timestamp 1621261055
transform 1 0 35616 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_363
timestamp 1621261055
transform 1 0 36000 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_40_368
timestamp 1621261055
transform 1 0 36480 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_40_375
timestamp 1621261055
transform 1 0 37152 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_383
timestamp 1621261055
transform 1 0 37920 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_391
timestamp 1621261055
transform 1 0 38688 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_399
timestamp 1621261055
transform 1 0 39456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_601
timestamp 1621261055
transform 1 0 40800 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_407
timestamp 1621261055
transform 1 0 40224 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_411
timestamp 1621261055
transform 1 0 40608 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_414
timestamp 1621261055
transform 1 0 40896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_422
timestamp 1621261055
transform 1 0 41664 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_430
timestamp 1621261055
transform 1 0 42432 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_438
timestamp 1621261055
transform 1 0 43200 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_446
timestamp 1621261055
transform 1 0 43968 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_454
timestamp 1621261055
transform 1 0 44736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_462
timestamp 1621261055
transform 1 0 45504 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_602
timestamp 1621261055
transform 1 0 46080 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_466
timestamp 1621261055
transform 1 0 45888 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_469
timestamp 1621261055
transform 1 0 46176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_477
timestamp 1621261055
transform 1 0 46944 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_485
timestamp 1621261055
transform 1 0 47712 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_493
timestamp 1621261055
transform 1 0 48480 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_501
timestamp 1621261055
transform 1 0 49248 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_603
timestamp 1621261055
transform 1 0 51360 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_509
timestamp 1621261055
transform 1 0 50016 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_517
timestamp 1621261055
transform 1 0 50784 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_521
timestamp 1621261055
transform 1 0 51168 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_524
timestamp 1621261055
transform 1 0 51456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_532
timestamp 1621261055
transform 1 0 52224 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_540
timestamp 1621261055
transform 1 0 52992 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_548
timestamp 1621261055
transform 1 0 53760 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_556
timestamp 1621261055
transform 1 0 54528 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_564
timestamp 1621261055
transform 1 0 55296 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_604
timestamp 1621261055
transform 1 0 56640 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_572
timestamp 1621261055
transform 1 0 56064 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_576
timestamp 1621261055
transform 1 0 56448 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_579
timestamp 1621261055
transform 1 0 56736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_587
timestamp 1621261055
transform 1 0 57504 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_81
timestamp 1621261055
transform -1 0 58848 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_595
timestamp 1621261055
transform 1 0 58272 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_82
timestamp 1621261055
transform 1 0 1152 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_41_4
timestamp 1621261055
transform 1 0 1536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_12
timestamp 1621261055
transform 1 0 2304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_20
timestamp 1621261055
transform 1 0 3072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _160_
timestamp 1621261055
transform 1 0 4416 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_106
timestamp 1621261055
transform 1 0 4224 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_41_28
timestamp 1621261055
transform 1 0 3840 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_41_37
timestamp 1621261055
transform 1 0 4704 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_605
timestamp 1621261055
transform 1 0 6432 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_45
timestamp 1621261055
transform 1 0 5472 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_53
timestamp 1621261055
transform 1 0 6240 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_56
timestamp 1621261055
transform 1 0 6528 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_64
timestamp 1621261055
transform 1 0 7296 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_72
timestamp 1621261055
transform 1 0 8064 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_80
timestamp 1621261055
transform 1 0 8832 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_88
timestamp 1621261055
transform 1 0 9600 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_96
timestamp 1621261055
transform 1 0 10368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_104
timestamp 1621261055
transform 1 0 11136 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_606
timestamp 1621261055
transform 1 0 11712 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_108
timestamp 1621261055
transform 1 0 11520 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_111
timestamp 1621261055
transform 1 0 11808 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_119
timestamp 1621261055
transform 1 0 12576 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_127
timestamp 1621261055
transform 1 0 13344 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_135
timestamp 1621261055
transform 1 0 14112 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_143
timestamp 1621261055
transform 1 0 14880 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_607
timestamp 1621261055
transform 1 0 16992 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_151
timestamp 1621261055
transform 1 0 15648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_159
timestamp 1621261055
transform 1 0 16416 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_163
timestamp 1621261055
transform 1 0 16800 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_166
timestamp 1621261055
transform 1 0 17088 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_174
timestamp 1621261055
transform 1 0 17856 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_182
timestamp 1621261055
transform 1 0 18624 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_190
timestamp 1621261055
transform 1 0 19392 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_198
timestamp 1621261055
transform 1 0 20160 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_206
timestamp 1621261055
transform 1 0 20928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_608
timestamp 1621261055
transform 1 0 22272 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_214
timestamp 1621261055
transform 1 0 21696 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_218
timestamp 1621261055
transform 1 0 22080 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_221
timestamp 1621261055
transform 1 0 22368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_229
timestamp 1621261055
transform 1 0 23136 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_237
timestamp 1621261055
transform 1 0 23904 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_245
timestamp 1621261055
transform 1 0 24672 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_253
timestamp 1621261055
transform 1 0 25440 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_261
timestamp 1621261055
transform 1 0 26208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_269
timestamp 1621261055
transform 1 0 26976 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_273
timestamp 1621261055
transform 1 0 27360 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_609
timestamp 1621261055
transform 1 0 27552 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_276
timestamp 1621261055
transform 1 0 27648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_284
timestamp 1621261055
transform 1 0 28416 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_292
timestamp 1621261055
transform 1 0 29184 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_300
timestamp 1621261055
transform 1 0 29952 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_308
timestamp 1621261055
transform 1 0 30720 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_610
timestamp 1621261055
transform 1 0 32832 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_316
timestamp 1621261055
transform 1 0 31488 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_324
timestamp 1621261055
transform 1 0 32256 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_328
timestamp 1621261055
transform 1 0 32640 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_331
timestamp 1621261055
transform 1 0 32928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_339
timestamp 1621261055
transform 1 0 33696 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_347
timestamp 1621261055
transform 1 0 34464 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_355
timestamp 1621261055
transform 1 0 35232 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_363
timestamp 1621261055
transform 1 0 36000 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_371
timestamp 1621261055
transform 1 0 36768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _162_
timestamp 1621261055
transform 1 0 38688 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_611
timestamp 1621261055
transform 1 0 38112 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_379
timestamp 1621261055
transform 1 0 37536 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_383
timestamp 1621261055
transform 1 0 37920 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_41_386
timestamp 1621261055
transform 1 0 38208 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_41_390
timestamp 1621261055
transform 1 0 38592 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_394
timestamp 1621261055
transform 1 0 38976 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_402
timestamp 1621261055
transform 1 0 39744 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_410
timestamp 1621261055
transform 1 0 40512 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_418
timestamp 1621261055
transform 1 0 41280 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_612
timestamp 1621261055
transform 1 0 43392 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_426
timestamp 1621261055
transform 1 0 42048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_434
timestamp 1621261055
transform 1 0 42816 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_438
timestamp 1621261055
transform 1 0 43200 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_441
timestamp 1621261055
transform 1 0 43488 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_449
timestamp 1621261055
transform 1 0 44256 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_457
timestamp 1621261055
transform 1 0 45024 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_465
timestamp 1621261055
transform 1 0 45792 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_473
timestamp 1621261055
transform 1 0 46560 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_481
timestamp 1621261055
transform 1 0 47328 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_613
timestamp 1621261055
transform 1 0 48672 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_489
timestamp 1621261055
transform 1 0 48096 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_493
timestamp 1621261055
transform 1 0 48480 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_496
timestamp 1621261055
transform 1 0 48768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_504
timestamp 1621261055
transform 1 0 49536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_512
timestamp 1621261055
transform 1 0 50304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_520
timestamp 1621261055
transform 1 0 51072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_528
timestamp 1621261055
transform 1 0 51840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_536
timestamp 1621261055
transform 1 0 52608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_544
timestamp 1621261055
transform 1 0 53376 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_614
timestamp 1621261055
transform 1 0 53952 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_548
timestamp 1621261055
transform 1 0 53760 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_551
timestamp 1621261055
transform 1 0 54048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_559
timestamp 1621261055
transform 1 0 54816 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_567
timestamp 1621261055
transform 1 0 55584 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_575
timestamp 1621261055
transform 1 0 56352 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_583
timestamp 1621261055
transform 1 0 57120 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_83
timestamp 1621261055
transform -1 0 58848 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_41_591
timestamp 1621261055
transform 1 0 57888 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_595
timestamp 1621261055
transform 1 0 58272 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_84
timestamp 1621261055
transform 1 0 1152 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_42_4
timestamp 1621261055
transform 1 0 1536 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_12
timestamp 1621261055
transform 1 0 2304 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_20
timestamp 1621261055
transform 1 0 3072 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_615
timestamp 1621261055
transform 1 0 3840 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_29
timestamp 1621261055
transform 1 0 3936 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_37
timestamp 1621261055
transform 1 0 4704 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _073_
timestamp 1621261055
transform 1 0 6720 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_45
timestamp 1621261055
transform 1 0 5472 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_53
timestamp 1621261055
transform 1 0 6240 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_42_57
timestamp 1621261055
transform 1 0 6624 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_61
timestamp 1621261055
transform 1 0 7008 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_616
timestamp 1621261055
transform 1 0 9120 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_69
timestamp 1621261055
transform 1 0 7776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_77
timestamp 1621261055
transform 1 0 8544 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_81
timestamp 1621261055
transform 1 0 8928 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_84
timestamp 1621261055
transform 1 0 9216 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_92
timestamp 1621261055
transform 1 0 9984 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_100
timestamp 1621261055
transform 1 0 10752 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_108
timestamp 1621261055
transform 1 0 11520 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_116
timestamp 1621261055
transform 1 0 12288 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_124
timestamp 1621261055
transform 1 0 13056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_617
timestamp 1621261055
transform 1 0 14400 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_132
timestamp 1621261055
transform 1 0 13824 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_136
timestamp 1621261055
transform 1 0 14208 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_139
timestamp 1621261055
transform 1 0 14496 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_147
timestamp 1621261055
transform 1 0 15264 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_155
timestamp 1621261055
transform 1 0 16032 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_163
timestamp 1621261055
transform 1 0 16800 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _144_
timestamp 1621261055
transform 1 0 18816 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_171
timestamp 1621261055
transform 1 0 17568 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_179
timestamp 1621261055
transform 1 0 18336 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_42_183
timestamp 1621261055
transform 1 0 18720 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_187
timestamp 1621261055
transform 1 0 19104 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _005_
timestamp 1621261055
transform 1 0 20544 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_618
timestamp 1621261055
transform 1 0 19680 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_191
timestamp 1621261055
transform 1 0 19488 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_194
timestamp 1621261055
transform 1 0 19776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_205
timestamp 1621261055
transform 1 0 20832 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_213
timestamp 1621261055
transform 1 0 21600 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_221
timestamp 1621261055
transform 1 0 22368 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_229
timestamp 1621261055
transform 1 0 23136 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_619
timestamp 1621261055
transform 1 0 24960 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_237
timestamp 1621261055
transform 1 0 23904 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_245
timestamp 1621261055
transform 1 0 24672 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_42_247
timestamp 1621261055
transform 1 0 24864 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_249
timestamp 1621261055
transform 1 0 25056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_257
timestamp 1621261055
transform 1 0 25824 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_265
timestamp 1621261055
transform 1 0 26592 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_273
timestamp 1621261055
transform 1 0 27360 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_281
timestamp 1621261055
transform 1 0 28128 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_289
timestamp 1621261055
transform 1 0 28896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_620
timestamp 1621261055
transform 1 0 30240 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_297
timestamp 1621261055
transform 1 0 29664 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_301
timestamp 1621261055
transform 1 0 30048 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_304
timestamp 1621261055
transform 1 0 30336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_312
timestamp 1621261055
transform 1 0 31104 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_320
timestamp 1621261055
transform 1 0 31872 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_328
timestamp 1621261055
transform 1 0 32640 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_336
timestamp 1621261055
transform 1 0 33408 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_344
timestamp 1621261055
transform 1 0 34176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_352
timestamp 1621261055
transform 1 0 34944 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_356
timestamp 1621261055
transform 1 0 35328 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_621
timestamp 1621261055
transform 1 0 35520 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_359
timestamp 1621261055
transform 1 0 35616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_367
timestamp 1621261055
transform 1 0 36384 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_375
timestamp 1621261055
transform 1 0 37152 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_383
timestamp 1621261055
transform 1 0 37920 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_391
timestamp 1621261055
transform 1 0 38688 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_399
timestamp 1621261055
transform 1 0 39456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_622
timestamp 1621261055
transform 1 0 40800 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_407
timestamp 1621261055
transform 1 0 40224 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_411
timestamp 1621261055
transform 1 0 40608 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_414
timestamp 1621261055
transform 1 0 40896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_422
timestamp 1621261055
transform 1 0 41664 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_430
timestamp 1621261055
transform 1 0 42432 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_438
timestamp 1621261055
transform 1 0 43200 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_446
timestamp 1621261055
transform 1 0 43968 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_454
timestamp 1621261055
transform 1 0 44736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_462
timestamp 1621261055
transform 1 0 45504 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_623
timestamp 1621261055
transform 1 0 46080 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_466
timestamp 1621261055
transform 1 0 45888 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_469
timestamp 1621261055
transform 1 0 46176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_477
timestamp 1621261055
transform 1 0 46944 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_485
timestamp 1621261055
transform 1 0 47712 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_493
timestamp 1621261055
transform 1 0 48480 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_501
timestamp 1621261055
transform 1 0 49248 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_624
timestamp 1621261055
transform 1 0 51360 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_509
timestamp 1621261055
transform 1 0 50016 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_517
timestamp 1621261055
transform 1 0 50784 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_521
timestamp 1621261055
transform 1 0 51168 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_42_524
timestamp 1621261055
transform 1 0 51456 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _081_
timestamp 1621261055
transform 1 0 53184 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _123_
timestamp 1621261055
transform 1 0 51840 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_531
timestamp 1621261055
transform 1 0 52128 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_539
timestamp 1621261055
transform 1 0 52896 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_42_541
timestamp 1621261055
transform 1 0 53088 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_545
timestamp 1621261055
transform 1 0 53472 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _100_
timestamp 1621261055
transform 1 0 55104 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_553
timestamp 1621261055
transform 1 0 54240 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_42_561
timestamp 1621261055
transform 1 0 55008 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_565
timestamp 1621261055
transform 1 0 55392 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_625
timestamp 1621261055
transform 1 0 56640 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_573
timestamp 1621261055
transform 1 0 56160 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_42_577
timestamp 1621261055
transform 1 0 56544 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_579
timestamp 1621261055
transform 1 0 56736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_587
timestamp 1621261055
transform 1 0 57504 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_85
timestamp 1621261055
transform -1 0 58848 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_595
timestamp 1621261055
transform 1 0 58272 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_86
timestamp 1621261055
transform 1 0 1152 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_43_4
timestamp 1621261055
transform 1 0 1536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_12
timestamp 1621261055
transform 1 0 2304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_20
timestamp 1621261055
transform 1 0 3072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_28
timestamp 1621261055
transform 1 0 3840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_36
timestamp 1621261055
transform 1 0 4608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_626
timestamp 1621261055
transform 1 0 6432 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_44
timestamp 1621261055
transform 1 0 5376 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_52
timestamp 1621261055
transform 1 0 6144 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_43_54
timestamp 1621261055
transform 1 0 6336 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_56
timestamp 1621261055
transform 1 0 6528 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_64
timestamp 1621261055
transform 1 0 7296 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_72
timestamp 1621261055
transform 1 0 8064 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_80
timestamp 1621261055
transform 1 0 8832 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_88
timestamp 1621261055
transform 1 0 9600 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_96
timestamp 1621261055
transform 1 0 10368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_104
timestamp 1621261055
transform 1 0 11136 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_627
timestamp 1621261055
transform 1 0 11712 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_108
timestamp 1621261055
transform 1 0 11520 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_111
timestamp 1621261055
transform 1 0 11808 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_119
timestamp 1621261055
transform 1 0 12576 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_127
timestamp 1621261055
transform 1 0 13344 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_135
timestamp 1621261055
transform 1 0 14112 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_143
timestamp 1621261055
transform 1 0 14880 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_628
timestamp 1621261055
transform 1 0 16992 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_151
timestamp 1621261055
transform 1 0 15648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_159
timestamp 1621261055
transform 1 0 16416 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_163
timestamp 1621261055
transform 1 0 16800 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_166
timestamp 1621261055
transform 1 0 17088 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_174
timestamp 1621261055
transform 1 0 17856 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_182
timestamp 1621261055
transform 1 0 18624 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_190
timestamp 1621261055
transform 1 0 19392 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_198
timestamp 1621261055
transform 1 0 20160 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_206
timestamp 1621261055
transform 1 0 20928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_629
timestamp 1621261055
transform 1 0 22272 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_214
timestamp 1621261055
transform 1 0 21696 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_218
timestamp 1621261055
transform 1 0 22080 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_221
timestamp 1621261055
transform 1 0 22368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_229
timestamp 1621261055
transform 1 0 23136 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_237
timestamp 1621261055
transform 1 0 23904 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_245
timestamp 1621261055
transform 1 0 24672 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_253
timestamp 1621261055
transform 1 0 25440 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_261
timestamp 1621261055
transform 1 0 26208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_269
timestamp 1621261055
transform 1 0 26976 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_273
timestamp 1621261055
transform 1 0 27360 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_630
timestamp 1621261055
transform 1 0 27552 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_276
timestamp 1621261055
transform 1 0 27648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_284
timestamp 1621261055
transform 1 0 28416 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_292
timestamp 1621261055
transform 1 0 29184 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_300
timestamp 1621261055
transform 1 0 29952 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_308
timestamp 1621261055
transform 1 0 30720 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_631
timestamp 1621261055
transform 1 0 32832 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_316
timestamp 1621261055
transform 1 0 31488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_324
timestamp 1621261055
transform 1 0 32256 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_328
timestamp 1621261055
transform 1 0 32640 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_331
timestamp 1621261055
transform 1 0 32928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_339
timestamp 1621261055
transform 1 0 33696 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_347
timestamp 1621261055
transform 1 0 34464 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_355
timestamp 1621261055
transform 1 0 35232 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_363
timestamp 1621261055
transform 1 0 36000 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_371
timestamp 1621261055
transform 1 0 36768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_632
timestamp 1621261055
transform 1 0 38112 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_379
timestamp 1621261055
transform 1 0 37536 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_383
timestamp 1621261055
transform 1 0 37920 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_386
timestamp 1621261055
transform 1 0 38208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_394
timestamp 1621261055
transform 1 0 38976 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_402
timestamp 1621261055
transform 1 0 39744 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_410
timestamp 1621261055
transform 1 0 40512 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_418
timestamp 1621261055
transform 1 0 41280 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_633
timestamp 1621261055
transform 1 0 43392 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_426
timestamp 1621261055
transform 1 0 42048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_434
timestamp 1621261055
transform 1 0 42816 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_438
timestamp 1621261055
transform 1 0 43200 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_441
timestamp 1621261055
transform 1 0 43488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_449
timestamp 1621261055
transform 1 0 44256 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_457
timestamp 1621261055
transform 1 0 45024 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_465
timestamp 1621261055
transform 1 0 45792 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_473
timestamp 1621261055
transform 1 0 46560 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_481
timestamp 1621261055
transform 1 0 47328 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_634
timestamp 1621261055
transform 1 0 48672 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_489
timestamp 1621261055
transform 1 0 48096 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_493
timestamp 1621261055
transform 1 0 48480 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_496
timestamp 1621261055
transform 1 0 48768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_504
timestamp 1621261055
transform 1 0 49536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_512
timestamp 1621261055
transform 1 0 50304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_520
timestamp 1621261055
transform 1 0 51072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _117_
timestamp 1621261055
transform 1 0 52608 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_43_528
timestamp 1621261055
transform 1 0 51840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_539
timestamp 1621261055
transform 1 0 52896 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_635
timestamp 1621261055
transform 1 0 53952 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_547
timestamp 1621261055
transform 1 0 53664 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_43_549
timestamp 1621261055
transform 1 0 53856 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_551
timestamp 1621261055
transform 1 0 54048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_559
timestamp 1621261055
transform 1 0 54816 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_567
timestamp 1621261055
transform 1 0 55584 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_575
timestamp 1621261055
transform 1 0 56352 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_583
timestamp 1621261055
transform 1 0 57120 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_87
timestamp 1621261055
transform -1 0 58848 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_43_591
timestamp 1621261055
transform 1 0 57888 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_595
timestamp 1621261055
transform 1 0 58272 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_88
timestamp 1621261055
transform 1 0 1152 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_44_4
timestamp 1621261055
transform 1 0 1536 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_12
timestamp 1621261055
transform 1 0 2304 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_20
timestamp 1621261055
transform 1 0 3072 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_636
timestamp 1621261055
transform 1 0 3840 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_29
timestamp 1621261055
transform 1 0 3936 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_37
timestamp 1621261055
transform 1 0 4704 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _167_
timestamp 1621261055
transform 1 0 5664 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_45
timestamp 1621261055
transform 1 0 5472 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_50
timestamp 1621261055
transform 1 0 5952 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_58
timestamp 1621261055
transform 1 0 6720 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_637
timestamp 1621261055
transform 1 0 9120 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_66
timestamp 1621261055
transform 1 0 7488 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_74
timestamp 1621261055
transform 1 0 8256 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_44_82
timestamp 1621261055
transform 1 0 9024 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_84
timestamp 1621261055
transform 1 0 9216 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_92
timestamp 1621261055
transform 1 0 9984 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_100
timestamp 1621261055
transform 1 0 10752 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_108
timestamp 1621261055
transform 1 0 11520 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_116
timestamp 1621261055
transform 1 0 12288 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_124
timestamp 1621261055
transform 1 0 13056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_638
timestamp 1621261055
transform 1 0 14400 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_132
timestamp 1621261055
transform 1 0 13824 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_136
timestamp 1621261055
transform 1 0 14208 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_139
timestamp 1621261055
transform 1 0 14496 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_147
timestamp 1621261055
transform 1 0 15264 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_155
timestamp 1621261055
transform 1 0 16032 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_163
timestamp 1621261055
transform 1 0 16800 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_171
timestamp 1621261055
transform 1 0 17568 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_179
timestamp 1621261055
transform 1 0 18336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_187
timestamp 1621261055
transform 1 0 19104 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_639
timestamp 1621261055
transform 1 0 19680 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_191
timestamp 1621261055
transform 1 0 19488 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_194
timestamp 1621261055
transform 1 0 19776 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_202
timestamp 1621261055
transform 1 0 20544 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_44_210
timestamp 1621261055
transform 1 0 21312 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _121_
timestamp 1621261055
transform 1 0 21408 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_44_214
timestamp 1621261055
transform 1 0 21696 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_222
timestamp 1621261055
transform 1 0 22464 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_230
timestamp 1621261055
transform 1 0 23232 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_640
timestamp 1621261055
transform 1 0 24960 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_238
timestamp 1621261055
transform 1 0 24000 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_246
timestamp 1621261055
transform 1 0 24768 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_249
timestamp 1621261055
transform 1 0 25056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _055_
timestamp 1621261055
transform 1 0 26016 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _159_
timestamp 1621261055
transform 1 0 27168 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_257
timestamp 1621261055
transform 1 0 25824 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_262
timestamp 1621261055
transform 1 0 26304 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_44_270
timestamp 1621261055
transform 1 0 27072 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_274
timestamp 1621261055
transform 1 0 27456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_282
timestamp 1621261055
transform 1 0 28224 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_290
timestamp 1621261055
transform 1 0 28992 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_641
timestamp 1621261055
transform 1 0 30240 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_298
timestamp 1621261055
transform 1 0 29760 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_44_302
timestamp 1621261055
transform 1 0 30144 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_304
timestamp 1621261055
transform 1 0 30336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_312
timestamp 1621261055
transform 1 0 31104 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_320
timestamp 1621261055
transform 1 0 31872 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_328
timestamp 1621261055
transform 1 0 32640 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_336
timestamp 1621261055
transform 1 0 33408 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_344
timestamp 1621261055
transform 1 0 34176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_352
timestamp 1621261055
transform 1 0 34944 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_356
timestamp 1621261055
transform 1 0 35328 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_642
timestamp 1621261055
transform 1 0 35520 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_359
timestamp 1621261055
transform 1 0 35616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_367
timestamp 1621261055
transform 1 0 36384 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_375
timestamp 1621261055
transform 1 0 37152 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_383
timestamp 1621261055
transform 1 0 37920 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_391
timestamp 1621261055
transform 1 0 38688 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_399
timestamp 1621261055
transform 1 0 39456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_643
timestamp 1621261055
transform 1 0 40800 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_407
timestamp 1621261055
transform 1 0 40224 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_411
timestamp 1621261055
transform 1 0 40608 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_414
timestamp 1621261055
transform 1 0 40896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_422
timestamp 1621261055
transform 1 0 41664 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_430
timestamp 1621261055
transform 1 0 42432 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_438
timestamp 1621261055
transform 1 0 43200 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_446
timestamp 1621261055
transform 1 0 43968 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_454
timestamp 1621261055
transform 1 0 44736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_462
timestamp 1621261055
transform 1 0 45504 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_644
timestamp 1621261055
transform 1 0 46080 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_466
timestamp 1621261055
transform 1 0 45888 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_469
timestamp 1621261055
transform 1 0 46176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_477
timestamp 1621261055
transform 1 0 46944 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_485
timestamp 1621261055
transform 1 0 47712 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_493
timestamp 1621261055
transform 1 0 48480 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_501
timestamp 1621261055
transform 1 0 49248 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_645
timestamp 1621261055
transform 1 0 51360 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_509
timestamp 1621261055
transform 1 0 50016 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_517
timestamp 1621261055
transform 1 0 50784 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_521
timestamp 1621261055
transform 1 0 51168 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_524
timestamp 1621261055
transform 1 0 51456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_532
timestamp 1621261055
transform 1 0 52224 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_540
timestamp 1621261055
transform 1 0 52992 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_548
timestamp 1621261055
transform 1 0 53760 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_556
timestamp 1621261055
transform 1 0 54528 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_564
timestamp 1621261055
transform 1 0 55296 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_646
timestamp 1621261055
transform 1 0 56640 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_572
timestamp 1621261055
transform 1 0 56064 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_576
timestamp 1621261055
transform 1 0 56448 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_579
timestamp 1621261055
transform 1 0 56736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_587
timestamp 1621261055
transform 1 0 57504 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_89
timestamp 1621261055
transform -1 0 58848 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_595
timestamp 1621261055
transform 1 0 58272 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_90
timestamp 1621261055
transform 1 0 1152 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_4
timestamp 1621261055
transform 1 0 1536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_12
timestamp 1621261055
transform 1 0 2304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_20
timestamp 1621261055
transform 1 0 3072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_28
timestamp 1621261055
transform 1 0 3840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_36
timestamp 1621261055
transform 1 0 4608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_647
timestamp 1621261055
transform 1 0 6432 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_44
timestamp 1621261055
transform 1 0 5376 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_52
timestamp 1621261055
transform 1 0 6144 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_54
timestamp 1621261055
transform 1 0 6336 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_56
timestamp 1621261055
transform 1 0 6528 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_64
timestamp 1621261055
transform 1 0 7296 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_72
timestamp 1621261055
transform 1 0 8064 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_80
timestamp 1621261055
transform 1 0 8832 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_88
timestamp 1621261055
transform 1 0 9600 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_96
timestamp 1621261055
transform 1 0 10368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_104
timestamp 1621261055
transform 1 0 11136 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_648
timestamp 1621261055
transform 1 0 11712 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_108
timestamp 1621261055
transform 1 0 11520 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_111
timestamp 1621261055
transform 1 0 11808 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_119
timestamp 1621261055
transform 1 0 12576 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_127
timestamp 1621261055
transform 1 0 13344 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_135
timestamp 1621261055
transform 1 0 14112 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_143
timestamp 1621261055
transform 1 0 14880 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_649
timestamp 1621261055
transform 1 0 16992 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_151
timestamp 1621261055
transform 1 0 15648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_159
timestamp 1621261055
transform 1 0 16416 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_163
timestamp 1621261055
transform 1 0 16800 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_166
timestamp 1621261055
transform 1 0 17088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_174
timestamp 1621261055
transform 1 0 17856 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_182
timestamp 1621261055
transform 1 0 18624 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_190
timestamp 1621261055
transform 1 0 19392 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_198
timestamp 1621261055
transform 1 0 20160 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_206
timestamp 1621261055
transform 1 0 20928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_650
timestamp 1621261055
transform 1 0 22272 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_214
timestamp 1621261055
transform 1 0 21696 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_218
timestamp 1621261055
transform 1 0 22080 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_221
timestamp 1621261055
transform 1 0 22368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_229
timestamp 1621261055
transform 1 0 23136 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_237
timestamp 1621261055
transform 1 0 23904 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_245
timestamp 1621261055
transform 1 0 24672 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_253
timestamp 1621261055
transform 1 0 25440 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_261
timestamp 1621261055
transform 1 0 26208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_269
timestamp 1621261055
transform 1 0 26976 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_273
timestamp 1621261055
transform 1 0 27360 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_651
timestamp 1621261055
transform 1 0 27552 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_276
timestamp 1621261055
transform 1 0 27648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_284
timestamp 1621261055
transform 1 0 28416 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_292
timestamp 1621261055
transform 1 0 29184 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_300
timestamp 1621261055
transform 1 0 29952 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_308
timestamp 1621261055
transform 1 0 30720 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_652
timestamp 1621261055
transform 1 0 32832 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_316
timestamp 1621261055
transform 1 0 31488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_324
timestamp 1621261055
transform 1 0 32256 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_328
timestamp 1621261055
transform 1 0 32640 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_331
timestamp 1621261055
transform 1 0 32928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_339
timestamp 1621261055
transform 1 0 33696 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_347
timestamp 1621261055
transform 1 0 34464 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_355
timestamp 1621261055
transform 1 0 35232 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_363
timestamp 1621261055
transform 1 0 36000 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_371
timestamp 1621261055
transform 1 0 36768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_653
timestamp 1621261055
transform 1 0 38112 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_379
timestamp 1621261055
transform 1 0 37536 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_383
timestamp 1621261055
transform 1 0 37920 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_386
timestamp 1621261055
transform 1 0 38208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_394
timestamp 1621261055
transform 1 0 38976 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_398
timestamp 1621261055
transform 1 0 39360 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _021_
timestamp 1621261055
transform 1 0 39552 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_45_403
timestamp 1621261055
transform 1 0 39840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_411
timestamp 1621261055
transform 1 0 40608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_419
timestamp 1621261055
transform 1 0 41376 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_654
timestamp 1621261055
transform 1 0 43392 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_427
timestamp 1621261055
transform 1 0 42144 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_435
timestamp 1621261055
transform 1 0 42912 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_45_439
timestamp 1621261055
transform 1 0 43296 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_441
timestamp 1621261055
transform 1 0 43488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_449
timestamp 1621261055
transform 1 0 44256 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_457
timestamp 1621261055
transform 1 0 45024 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_465
timestamp 1621261055
transform 1 0 45792 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_473
timestamp 1621261055
transform 1 0 46560 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_481
timestamp 1621261055
transform 1 0 47328 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_655
timestamp 1621261055
transform 1 0 48672 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_489
timestamp 1621261055
transform 1 0 48096 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_493
timestamp 1621261055
transform 1 0 48480 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_496
timestamp 1621261055
transform 1 0 48768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_504
timestamp 1621261055
transform 1 0 49536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_512
timestamp 1621261055
transform 1 0 50304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_520
timestamp 1621261055
transform 1 0 51072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_528
timestamp 1621261055
transform 1 0 51840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_536
timestamp 1621261055
transform 1 0 52608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_544
timestamp 1621261055
transform 1 0 53376 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_656
timestamp 1621261055
transform 1 0 53952 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_548
timestamp 1621261055
transform 1 0 53760 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_551
timestamp 1621261055
transform 1 0 54048 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_559
timestamp 1621261055
transform 1 0 54816 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_567
timestamp 1621261055
transform 1 0 55584 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_575
timestamp 1621261055
transform 1 0 56352 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_583
timestamp 1621261055
transform 1 0 57120 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_91
timestamp 1621261055
transform -1 0 58848 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_45_591
timestamp 1621261055
transform 1 0 57888 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_595
timestamp 1621261055
transform 1 0 58272 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_92
timestamp 1621261055
transform 1 0 1152 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_94
timestamp 1621261055
transform 1 0 1152 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_4
timestamp 1621261055
transform 1 0 1536 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_12
timestamp 1621261055
transform 1 0 2304 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_20
timestamp 1621261055
transform 1 0 3072 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_4
timestamp 1621261055
transform 1 0 1536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_12
timestamp 1621261055
transform 1 0 2304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_20
timestamp 1621261055
transform 1 0 3072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_657
timestamp 1621261055
transform 1 0 3840 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_29
timestamp 1621261055
transform 1 0 3936 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_37
timestamp 1621261055
transform 1 0 4704 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_28
timestamp 1621261055
transform 1 0 3840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_36
timestamp 1621261055
transform 1 0 4608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_668
timestamp 1621261055
transform 1 0 6432 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_45
timestamp 1621261055
transform 1 0 5472 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_53
timestamp 1621261055
transform 1 0 6240 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_61
timestamp 1621261055
transform 1 0 7008 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_44
timestamp 1621261055
transform 1 0 5376 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_52
timestamp 1621261055
transform 1 0 6144 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_47_54
timestamp 1621261055
transform 1 0 6336 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_56
timestamp 1621261055
transform 1 0 6528 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_658
timestamp 1621261055
transform 1 0 9120 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_69
timestamp 1621261055
transform 1 0 7776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_77
timestamp 1621261055
transform 1 0 8544 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_81
timestamp 1621261055
transform 1 0 8928 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_84
timestamp 1621261055
transform 1 0 9216 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_64
timestamp 1621261055
transform 1 0 7296 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_72
timestamp 1621261055
transform 1 0 8064 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_80
timestamp 1621261055
transform 1 0 8832 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_92
timestamp 1621261055
transform 1 0 9984 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_100
timestamp 1621261055
transform 1 0 10752 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_88
timestamp 1621261055
transform 1 0 9600 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_96
timestamp 1621261055
transform 1 0 10368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_104
timestamp 1621261055
transform 1 0 11136 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_669
timestamp 1621261055
transform 1 0 11712 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_108
timestamp 1621261055
transform 1 0 11520 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_116
timestamp 1621261055
transform 1 0 12288 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_124
timestamp 1621261055
transform 1 0 13056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_108
timestamp 1621261055
transform 1 0 11520 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_111
timestamp 1621261055
transform 1 0 11808 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_119
timestamp 1621261055
transform 1 0 12576 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_659
timestamp 1621261055
transform 1 0 14400 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_132
timestamp 1621261055
transform 1 0 13824 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_136
timestamp 1621261055
transform 1 0 14208 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_139
timestamp 1621261055
transform 1 0 14496 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_147
timestamp 1621261055
transform 1 0 15264 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_127
timestamp 1621261055
transform 1 0 13344 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_135
timestamp 1621261055
transform 1 0 14112 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_143
timestamp 1621261055
transform 1 0 14880 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _211_
timestamp 1621261055
transform 1 0 16608 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_670
timestamp 1621261055
transform 1 0 16992 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_155
timestamp 1621261055
transform 1 0 16032 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_159
timestamp 1621261055
transform 1 0 16416 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_164
timestamp 1621261055
transform 1 0 16896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_151
timestamp 1621261055
transform 1 0 15648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_159
timestamp 1621261055
transform 1 0 16416 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_163
timestamp 1621261055
transform 1 0 16800 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_166
timestamp 1621261055
transform 1 0 17088 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_172
timestamp 1621261055
transform 1 0 17664 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_180
timestamp 1621261055
transform 1 0 18432 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_188
timestamp 1621261055
transform 1 0 19200 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_174
timestamp 1621261055
transform 1 0 17856 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_182
timestamp 1621261055
transform 1 0 18624 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_660
timestamp 1621261055
transform 1 0 19680 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_46_192
timestamp 1621261055
transform 1 0 19584 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_194
timestamp 1621261055
transform 1 0 19776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_202
timestamp 1621261055
transform 1 0 20544 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_210
timestamp 1621261055
transform 1 0 21312 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_190
timestamp 1621261055
transform 1 0 19392 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_198
timestamp 1621261055
transform 1 0 20160 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_206
timestamp 1621261055
transform 1 0 20928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_671
timestamp 1621261055
transform 1 0 22272 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_218
timestamp 1621261055
transform 1 0 22080 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_226
timestamp 1621261055
transform 1 0 22848 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_214
timestamp 1621261055
transform 1 0 21696 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_218
timestamp 1621261055
transform 1 0 22080 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_221
timestamp 1621261055
transform 1 0 22368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_229
timestamp 1621261055
transform 1 0 23136 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_661
timestamp 1621261055
transform 1 0 24960 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_234
timestamp 1621261055
transform 1 0 23616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_242
timestamp 1621261055
transform 1 0 24384 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_246
timestamp 1621261055
transform 1 0 24768 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_249
timestamp 1621261055
transform 1 0 25056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_237
timestamp 1621261055
transform 1 0 23904 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_245
timestamp 1621261055
transform 1 0 24672 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _057_
timestamp 1621261055
transform 1 0 26496 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_46_257
timestamp 1621261055
transform 1 0 25824 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_261
timestamp 1621261055
transform 1 0 26208 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_46_263
timestamp 1621261055
transform 1 0 26400 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_267
timestamp 1621261055
transform 1 0 26784 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_253
timestamp 1621261055
transform 1 0 25440 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_261
timestamp 1621261055
transform 1 0 26208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_269
timestamp 1621261055
transform 1 0 26976 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_273
timestamp 1621261055
transform 1 0 27360 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _166_
timestamp 1621261055
transform 1 0 28032 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_672
timestamp 1621261055
transform 1 0 27552 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_275
timestamp 1621261055
transform 1 0 27552 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_283
timestamp 1621261055
transform 1 0 28320 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_291
timestamp 1621261055
transform 1 0 29088 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_276
timestamp 1621261055
transform 1 0 27648 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_283
timestamp 1621261055
transform 1 0 28320 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_291
timestamp 1621261055
transform 1 0 29088 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_662
timestamp 1621261055
transform 1 0 30240 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_299
timestamp 1621261055
transform 1 0 29856 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_304
timestamp 1621261055
transform 1 0 30336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_312
timestamp 1621261055
transform 1 0 31104 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_299
timestamp 1621261055
transform 1 0 29856 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_307
timestamp 1621261055
transform 1 0 30624 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_315
timestamp 1621261055
transform 1 0 31392 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_673
timestamp 1621261055
transform 1 0 32832 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_320
timestamp 1621261055
transform 1 0 31872 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_328
timestamp 1621261055
transform 1 0 32640 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_336
timestamp 1621261055
transform 1 0 33408 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_323
timestamp 1621261055
transform 1 0 32160 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_327
timestamp 1621261055
transform 1 0 32544 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_47_329
timestamp 1621261055
transform 1 0 32736 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_331
timestamp 1621261055
transform 1 0 32928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_344
timestamp 1621261055
transform 1 0 34176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_352
timestamp 1621261055
transform 1 0 34944 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_356
timestamp 1621261055
transform 1 0 35328 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_339
timestamp 1621261055
transform 1 0 33696 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_347
timestamp 1621261055
transform 1 0 34464 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_355
timestamp 1621261055
transform 1 0 35232 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _124_
timestamp 1621261055
transform 1 0 36000 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_663
timestamp 1621261055
transform 1 0 35520 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_190
timestamp 1621261055
transform 1 0 35808 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_359
timestamp 1621261055
transform 1 0 35616 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_366
timestamp 1621261055
transform 1 0 36288 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_374
timestamp 1621261055
transform 1 0 37056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_363
timestamp 1621261055
transform 1 0 36000 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_371
timestamp 1621261055
transform 1 0 36768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_674
timestamp 1621261055
transform 1 0 38112 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_382
timestamp 1621261055
transform 1 0 37824 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_390
timestamp 1621261055
transform 1 0 38592 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_398
timestamp 1621261055
transform 1 0 39360 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_379
timestamp 1621261055
transform 1 0 37536 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_383
timestamp 1621261055
transform 1 0 37920 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_386
timestamp 1621261055
transform 1 0 38208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_394
timestamp 1621261055
transform 1 0 38976 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_664
timestamp 1621261055
transform 1 0 40800 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_406
timestamp 1621261055
transform 1 0 40128 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_410
timestamp 1621261055
transform 1 0 40512 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_46_412
timestamp 1621261055
transform 1 0 40704 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_414
timestamp 1621261055
transform 1 0 40896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_402
timestamp 1621261055
transform 1 0 39744 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_410
timestamp 1621261055
transform 1 0 40512 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_418
timestamp 1621261055
transform 1 0 41280 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_675
timestamp 1621261055
transform 1 0 43392 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_422
timestamp 1621261055
transform 1 0 41664 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_430
timestamp 1621261055
transform 1 0 42432 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_438
timestamp 1621261055
transform 1 0 43200 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_426
timestamp 1621261055
transform 1 0 42048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_434
timestamp 1621261055
transform 1 0 42816 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_438
timestamp 1621261055
transform 1 0 43200 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_441
timestamp 1621261055
transform 1 0 43488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_446
timestamp 1621261055
transform 1 0 43968 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_454
timestamp 1621261055
transform 1 0 44736 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_462
timestamp 1621261055
transform 1 0 45504 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_449
timestamp 1621261055
transform 1 0 44256 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_457
timestamp 1621261055
transform 1 0 45024 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_665
timestamp 1621261055
transform 1 0 46080 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_466
timestamp 1621261055
transform 1 0 45888 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_469
timestamp 1621261055
transform 1 0 46176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_477
timestamp 1621261055
transform 1 0 46944 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_465
timestamp 1621261055
transform 1 0 45792 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_473
timestamp 1621261055
transform 1 0 46560 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_481
timestamp 1621261055
transform 1 0 47328 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_676
timestamp 1621261055
transform 1 0 48672 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_485
timestamp 1621261055
transform 1 0 47712 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_493
timestamp 1621261055
transform 1 0 48480 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_501
timestamp 1621261055
transform 1 0 49248 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_489
timestamp 1621261055
transform 1 0 48096 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_493
timestamp 1621261055
transform 1 0 48480 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_496
timestamp 1621261055
transform 1 0 48768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_504
timestamp 1621261055
transform 1 0 49536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_666
timestamp 1621261055
transform 1 0 51360 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_509
timestamp 1621261055
transform 1 0 50016 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_517
timestamp 1621261055
transform 1 0 50784 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_521
timestamp 1621261055
transform 1 0 51168 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_524
timestamp 1621261055
transform 1 0 51456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_512
timestamp 1621261055
transform 1 0 50304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_520
timestamp 1621261055
transform 1 0 51072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_532
timestamp 1621261055
transform 1 0 52224 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_540
timestamp 1621261055
transform 1 0 52992 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_528
timestamp 1621261055
transform 1 0 51840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_536
timestamp 1621261055
transform 1 0 52608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_544
timestamp 1621261055
transform 1 0 53376 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_677
timestamp 1621261055
transform 1 0 53952 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_548
timestamp 1621261055
transform 1 0 53760 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_556
timestamp 1621261055
transform 1 0 54528 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_564
timestamp 1621261055
transform 1 0 55296 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_548
timestamp 1621261055
transform 1 0 53760 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_551
timestamp 1621261055
transform 1 0 54048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_559
timestamp 1621261055
transform 1 0 54816 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_567
timestamp 1621261055
transform 1 0 55584 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_667
timestamp 1621261055
transform 1 0 56640 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_572
timestamp 1621261055
transform 1 0 56064 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_576
timestamp 1621261055
transform 1 0 56448 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_579
timestamp 1621261055
transform 1 0 56736 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_587
timestamp 1621261055
transform 1 0 57504 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_575
timestamp 1621261055
transform 1 0 56352 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_583
timestamp 1621261055
transform 1 0 57120 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_587
timestamp 1621261055
transform 1 0 57504 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _026_
timestamp 1621261055
transform 1 0 57792 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_93
timestamp 1621261055
transform -1 0 58848 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_95
timestamp 1621261055
transform -1 0 58848 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_595
timestamp 1621261055
transform 1 0 58272 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_47_589
timestamp 1621261055
transform 1 0 57696 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_47_593
timestamp 1621261055
transform 1 0 58080 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_96
timestamp 1621261055
transform 1 0 1152 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_4
timestamp 1621261055
transform 1 0 1536 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_12
timestamp 1621261055
transform 1 0 2304 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_20
timestamp 1621261055
transform 1 0 3072 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_678
timestamp 1621261055
transform 1 0 3840 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_29
timestamp 1621261055
transform 1 0 3936 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_37
timestamp 1621261055
transform 1 0 4704 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_45
timestamp 1621261055
transform 1 0 5472 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_53
timestamp 1621261055
transform 1 0 6240 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_61
timestamp 1621261055
transform 1 0 7008 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_679
timestamp 1621261055
transform 1 0 9120 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_69
timestamp 1621261055
transform 1 0 7776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_77
timestamp 1621261055
transform 1 0 8544 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_81
timestamp 1621261055
transform 1 0 8928 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_84
timestamp 1621261055
transform 1 0 9216 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_92
timestamp 1621261055
transform 1 0 9984 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_100
timestamp 1621261055
transform 1 0 10752 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_108
timestamp 1621261055
transform 1 0 11520 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_116
timestamp 1621261055
transform 1 0 12288 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_124
timestamp 1621261055
transform 1 0 13056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_680
timestamp 1621261055
transform 1 0 14400 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_132
timestamp 1621261055
transform 1 0 13824 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_136
timestamp 1621261055
transform 1 0 14208 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_139
timestamp 1621261055
transform 1 0 14496 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_147
timestamp 1621261055
transform 1 0 15264 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _093_
timestamp 1621261055
transform 1 0 15648 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_164
timestamp 1621261055
transform 1 0 15456 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_154
timestamp 1621261055
transform 1 0 15936 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_162
timestamp 1621261055
transform 1 0 16704 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_170
timestamp 1621261055
transform 1 0 17472 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_178
timestamp 1621261055
transform 1 0 18240 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_186
timestamp 1621261055
transform 1 0 19008 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_681
timestamp 1621261055
transform 1 0 19680 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_190
timestamp 1621261055
transform 1 0 19392 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_192
timestamp 1621261055
transform 1 0 19584 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_194
timestamp 1621261055
transform 1 0 19776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_202
timestamp 1621261055
transform 1 0 20544 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_210
timestamp 1621261055
transform 1 0 21312 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_218
timestamp 1621261055
transform 1 0 22080 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_226
timestamp 1621261055
transform 1 0 22848 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_682
timestamp 1621261055
transform 1 0 24960 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_234
timestamp 1621261055
transform 1 0 23616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_242
timestamp 1621261055
transform 1 0 24384 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_246
timestamp 1621261055
transform 1 0 24768 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_249
timestamp 1621261055
transform 1 0 25056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_257
timestamp 1621261055
transform 1 0 25824 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_265
timestamp 1621261055
transform 1 0 26592 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_273
timestamp 1621261055
transform 1 0 27360 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_281
timestamp 1621261055
transform 1 0 28128 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_289
timestamp 1621261055
transform 1 0 28896 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _050_
timestamp 1621261055
transform 1 0 30720 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_683
timestamp 1621261055
transform 1 0 30240 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_217
timestamp 1621261055
transform -1 0 31488 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_297
timestamp 1621261055
transform 1 0 29664 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_301
timestamp 1621261055
transform 1 0 30048 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_304
timestamp 1621261055
transform 1 0 30336 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_311
timestamp 1621261055
transform 1 0 31008 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_313
timestamp 1621261055
transform 1 0 31200 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _200_
timestamp 1621261055
transform -1 0 31776 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_48_319
timestamp 1621261055
transform 1 0 31776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_327
timestamp 1621261055
transform 1 0 32544 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_335
timestamp 1621261055
transform 1 0 33312 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_343
timestamp 1621261055
transform 1 0 34080 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_351
timestamp 1621261055
transform 1 0 34848 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_355
timestamp 1621261055
transform 1 0 35232 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_357
timestamp 1621261055
transform 1 0 35424 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_684
timestamp 1621261055
transform 1 0 35520 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_359
timestamp 1621261055
transform 1 0 35616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_367
timestamp 1621261055
transform 1 0 36384 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_375
timestamp 1621261055
transform 1 0 37152 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_383
timestamp 1621261055
transform 1 0 37920 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_391
timestamp 1621261055
transform 1 0 38688 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_399
timestamp 1621261055
transform 1 0 39456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_685
timestamp 1621261055
transform 1 0 40800 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_407
timestamp 1621261055
transform 1 0 40224 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_411
timestamp 1621261055
transform 1 0 40608 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_414
timestamp 1621261055
transform 1 0 40896 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_422
timestamp 1621261055
transform 1 0 41664 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_430
timestamp 1621261055
transform 1 0 42432 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_438
timestamp 1621261055
transform 1 0 43200 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_446
timestamp 1621261055
transform 1 0 43968 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_454
timestamp 1621261055
transform 1 0 44736 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_462
timestamp 1621261055
transform 1 0 45504 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_686
timestamp 1621261055
transform 1 0 46080 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_466
timestamp 1621261055
transform 1 0 45888 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_469
timestamp 1621261055
transform 1 0 46176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_477
timestamp 1621261055
transform 1 0 46944 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_485
timestamp 1621261055
transform 1 0 47712 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_493
timestamp 1621261055
transform 1 0 48480 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_501
timestamp 1621261055
transform 1 0 49248 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_687
timestamp 1621261055
transform 1 0 51360 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_509
timestamp 1621261055
transform 1 0 50016 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_517
timestamp 1621261055
transform 1 0 50784 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_521
timestamp 1621261055
transform 1 0 51168 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_524
timestamp 1621261055
transform 1 0 51456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _186_
timestamp 1621261055
transform -1 0 53472 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_211
timestamp 1621261055
transform -1 0 53184 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_532
timestamp 1621261055
transform 1 0 52224 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_545
timestamp 1621261055
transform 1 0 53472 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_553
timestamp 1621261055
transform 1 0 54240 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_561
timestamp 1621261055
transform 1 0 55008 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _091_
timestamp 1621261055
transform -1 0 57504 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_688
timestamp 1621261055
transform 1 0 56640 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_160
timestamp 1621261055
transform -1 0 57216 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_569
timestamp 1621261055
transform 1 0 55776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_48_577
timestamp 1621261055
transform 1 0 56544 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_579
timestamp 1621261055
transform 1 0 56736 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_581
timestamp 1621261055
transform 1 0 56928 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_587
timestamp 1621261055
transform 1 0 57504 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_97
timestamp 1621261055
transform -1 0 58848 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_595
timestamp 1621261055
transform 1 0 58272 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_98
timestamp 1621261055
transform 1 0 1152 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_49_4
timestamp 1621261055
transform 1 0 1536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_12
timestamp 1621261055
transform 1 0 2304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_20
timestamp 1621261055
transform 1 0 3072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_28
timestamp 1621261055
transform 1 0 3840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_36
timestamp 1621261055
transform 1 0 4608 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_689
timestamp 1621261055
transform 1 0 6432 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_44
timestamp 1621261055
transform 1 0 5376 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_52
timestamp 1621261055
transform 1 0 6144 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_54
timestamp 1621261055
transform 1 0 6336 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_56
timestamp 1621261055
transform 1 0 6528 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_64
timestamp 1621261055
transform 1 0 7296 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_72
timestamp 1621261055
transform 1 0 8064 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_80
timestamp 1621261055
transform 1 0 8832 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _191_
timestamp 1621261055
transform -1 0 11136 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_235
timestamp 1621261055
transform -1 0 10848 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_88
timestamp 1621261055
transform 1 0 9600 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_96
timestamp 1621261055
transform 1 0 10368 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_98
timestamp 1621261055
transform 1 0 10560 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_104
timestamp 1621261055
transform 1 0 11136 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_690
timestamp 1621261055
transform 1 0 11712 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_108
timestamp 1621261055
transform 1 0 11520 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_111
timestamp 1621261055
transform 1 0 11808 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_119
timestamp 1621261055
transform 1 0 12576 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_127
timestamp 1621261055
transform 1 0 13344 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_135
timestamp 1621261055
transform 1 0 14112 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_143
timestamp 1621261055
transform 1 0 14880 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_691
timestamp 1621261055
transform 1 0 16992 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_151
timestamp 1621261055
transform 1 0 15648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_159
timestamp 1621261055
transform 1 0 16416 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_163
timestamp 1621261055
transform 1 0 16800 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_166
timestamp 1621261055
transform 1 0 17088 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_174
timestamp 1621261055
transform 1 0 17856 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_182
timestamp 1621261055
transform 1 0 18624 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _085_
timestamp 1621261055
transform 1 0 20448 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _163_
timestamp 1621261055
transform 1 0 21120 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_108
timestamp 1621261055
transform 1 0 20928 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_148
timestamp 1621261055
transform 1 0 20256 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_190
timestamp 1621261055
transform 1 0 19392 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_49_198
timestamp 1621261055
transform 1 0 20160 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_204
timestamp 1621261055
transform 1 0 20736 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_692
timestamp 1621261055
transform 1 0 22272 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_211
timestamp 1621261055
transform 1 0 21408 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_49_219
timestamp 1621261055
transform 1 0 22176 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_221
timestamp 1621261055
transform 1 0 22368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_229
timestamp 1621261055
transform 1 0 23136 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_237
timestamp 1621261055
transform 1 0 23904 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_245
timestamp 1621261055
transform 1 0 24672 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_253
timestamp 1621261055
transform 1 0 25440 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_261
timestamp 1621261055
transform 1 0 26208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_269
timestamp 1621261055
transform 1 0 26976 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_273
timestamp 1621261055
transform 1 0 27360 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_693
timestamp 1621261055
transform 1 0 27552 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_276
timestamp 1621261055
transform 1 0 27648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_284
timestamp 1621261055
transform 1 0 28416 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_292
timestamp 1621261055
transform 1 0 29184 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_300
timestamp 1621261055
transform 1 0 29952 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_308
timestamp 1621261055
transform 1 0 30720 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_694
timestamp 1621261055
transform 1 0 32832 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_316
timestamp 1621261055
transform 1 0 31488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_324
timestamp 1621261055
transform 1 0 32256 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_328
timestamp 1621261055
transform 1 0 32640 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_331
timestamp 1621261055
transform 1 0 32928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_339
timestamp 1621261055
transform 1 0 33696 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_347
timestamp 1621261055
transform 1 0 34464 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_355
timestamp 1621261055
transform 1 0 35232 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_363
timestamp 1621261055
transform 1 0 36000 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_371
timestamp 1621261055
transform 1 0 36768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_695
timestamp 1621261055
transform 1 0 38112 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_379
timestamp 1621261055
transform 1 0 37536 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_383
timestamp 1621261055
transform 1 0 37920 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_386
timestamp 1621261055
transform 1 0 38208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_394
timestamp 1621261055
transform 1 0 38976 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_402
timestamp 1621261055
transform 1 0 39744 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_410
timestamp 1621261055
transform 1 0 40512 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_418
timestamp 1621261055
transform 1 0 41280 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_696
timestamp 1621261055
transform 1 0 43392 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_426
timestamp 1621261055
transform 1 0 42048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_434
timestamp 1621261055
transform 1 0 42816 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_438
timestamp 1621261055
transform 1 0 43200 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_441
timestamp 1621261055
transform 1 0 43488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_449
timestamp 1621261055
transform 1 0 44256 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_457
timestamp 1621261055
transform 1 0 45024 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_465
timestamp 1621261055
transform 1 0 45792 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_473
timestamp 1621261055
transform 1 0 46560 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_481
timestamp 1621261055
transform 1 0 47328 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_697
timestamp 1621261055
transform 1 0 48672 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_489
timestamp 1621261055
transform 1 0 48096 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_493
timestamp 1621261055
transform 1 0 48480 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_496
timestamp 1621261055
transform 1 0 48768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_504
timestamp 1621261055
transform 1 0 49536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_512
timestamp 1621261055
transform 1 0 50304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_520
timestamp 1621261055
transform 1 0 51072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _068_
timestamp 1621261055
transform -1 0 53088 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_110
timestamp 1621261055
transform -1 0 52800 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_528
timestamp 1621261055
transform 1 0 51840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_541
timestamp 1621261055
transform 1 0 53088 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_698
timestamp 1621261055
transform 1 0 53952 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_49_549
timestamp 1621261055
transform 1 0 53856 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_551
timestamp 1621261055
transform 1 0 54048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_559
timestamp 1621261055
transform 1 0 54816 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_567
timestamp 1621261055
transform 1 0 55584 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _201_
timestamp 1621261055
transform -1 0 56928 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_219
timestamp 1621261055
transform -1 0 56640 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_575
timestamp 1621261055
transform 1 0 56352 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_581
timestamp 1621261055
transform 1 0 56928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_99
timestamp 1621261055
transform -1 0 58848 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_49_589
timestamp 1621261055
transform 1 0 57696 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_100
timestamp 1621261055
transform 1 0 1152 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_4
timestamp 1621261055
transform 1 0 1536 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_12
timestamp 1621261055
transform 1 0 2304 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_20
timestamp 1621261055
transform 1 0 3072 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_699
timestamp 1621261055
transform 1 0 3840 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_29
timestamp 1621261055
transform 1 0 3936 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_37
timestamp 1621261055
transform 1 0 4704 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_45
timestamp 1621261055
transform 1 0 5472 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_53
timestamp 1621261055
transform 1 0 6240 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_61
timestamp 1621261055
transform 1 0 7008 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_700
timestamp 1621261055
transform 1 0 9120 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_69
timestamp 1621261055
transform 1 0 7776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_77
timestamp 1621261055
transform 1 0 8544 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_81
timestamp 1621261055
transform 1 0 8928 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_50_84
timestamp 1621261055
transform 1 0 9216 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _079_
timestamp 1621261055
transform 1 0 9600 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_50_91
timestamp 1621261055
transform 1 0 9888 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_99
timestamp 1621261055
transform 1 0 10656 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_107
timestamp 1621261055
transform 1 0 11424 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_115
timestamp 1621261055
transform 1 0 12192 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_123
timestamp 1621261055
transform 1 0 12960 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_701
timestamp 1621261055
transform 1 0 14400 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_131
timestamp 1621261055
transform 1 0 13728 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_135
timestamp 1621261055
transform 1 0 14112 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_50_137
timestamp 1621261055
transform 1 0 14304 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_139
timestamp 1621261055
transform 1 0 14496 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_147
timestamp 1621261055
transform 1 0 15264 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _189_
timestamp 1621261055
transform -1 0 17376 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_231
timestamp 1621261055
transform -1 0 17088 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_155
timestamp 1621261055
transform 1 0 16032 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_50_163
timestamp 1621261055
transform 1 0 16800 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_169
timestamp 1621261055
transform 1 0 17376 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_177
timestamp 1621261055
transform 1 0 18144 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_185
timestamp 1621261055
transform 1 0 18912 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _071_
timestamp 1621261055
transform -1 0 21120 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_702
timestamp 1621261055
transform 1 0 19680 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_132
timestamp 1621261055
transform -1 0 20832 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_194
timestamp 1621261055
transform 1 0 19776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_50_202
timestamp 1621261055
transform 1 0 20544 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_208
timestamp 1621261055
transform 1 0 21120 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_216
timestamp 1621261055
transform 1 0 21888 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_224
timestamp 1621261055
transform 1 0 22656 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_703
timestamp 1621261055
transform 1 0 24960 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_232
timestamp 1621261055
transform 1 0 23424 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_240
timestamp 1621261055
transform 1 0 24192 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_249
timestamp 1621261055
transform 1 0 25056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_257
timestamp 1621261055
transform 1 0 25824 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_265
timestamp 1621261055
transform 1 0 26592 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_273
timestamp 1621261055
transform 1 0 27360 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_281
timestamp 1621261055
transform 1 0 28128 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_289
timestamp 1621261055
transform 1 0 28896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_704
timestamp 1621261055
transform 1 0 30240 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_297
timestamp 1621261055
transform 1 0 29664 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_301
timestamp 1621261055
transform 1 0 30048 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_304
timestamp 1621261055
transform 1 0 30336 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_312
timestamp 1621261055
transform 1 0 31104 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_320
timestamp 1621261055
transform 1 0 31872 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_328
timestamp 1621261055
transform 1 0 32640 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_336
timestamp 1621261055
transform 1 0 33408 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_344
timestamp 1621261055
transform 1 0 34176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_352
timestamp 1621261055
transform 1 0 34944 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_356
timestamp 1621261055
transform 1 0 35328 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_705
timestamp 1621261055
transform 1 0 35520 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_359
timestamp 1621261055
transform 1 0 35616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_367
timestamp 1621261055
transform 1 0 36384 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_375
timestamp 1621261055
transform 1 0 37152 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_383
timestamp 1621261055
transform 1 0 37920 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_391
timestamp 1621261055
transform 1 0 38688 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_399
timestamp 1621261055
transform 1 0 39456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_706
timestamp 1621261055
transform 1 0 40800 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_407
timestamp 1621261055
transform 1 0 40224 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_411
timestamp 1621261055
transform 1 0 40608 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_414
timestamp 1621261055
transform 1 0 40896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_422
timestamp 1621261055
transform 1 0 41664 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_430
timestamp 1621261055
transform 1 0 42432 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_438
timestamp 1621261055
transform 1 0 43200 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _209_
timestamp 1621261055
transform -1 0 44832 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_223
timestamp 1621261055
transform -1 0 44544 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_50_446
timestamp 1621261055
transform 1 0 43968 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_455
timestamp 1621261055
transform 1 0 44832 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_707
timestamp 1621261055
transform 1 0 46080 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_463
timestamp 1621261055
transform 1 0 45600 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_50_467
timestamp 1621261055
transform 1 0 45984 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_469
timestamp 1621261055
transform 1 0 46176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_477
timestamp 1621261055
transform 1 0 46944 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_485
timestamp 1621261055
transform 1 0 47712 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_493
timestamp 1621261055
transform 1 0 48480 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_501
timestamp 1621261055
transform 1 0 49248 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_708
timestamp 1621261055
transform 1 0 51360 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_509
timestamp 1621261055
transform 1 0 50016 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_517
timestamp 1621261055
transform 1 0 50784 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_521
timestamp 1621261055
transform 1 0 51168 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_524
timestamp 1621261055
transform 1 0 51456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_532
timestamp 1621261055
transform 1 0 52224 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_540
timestamp 1621261055
transform 1 0 52992 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_548
timestamp 1621261055
transform 1 0 53760 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_556
timestamp 1621261055
transform 1 0 54528 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_564
timestamp 1621261055
transform 1 0 55296 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_709
timestamp 1621261055
transform 1 0 56640 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_572
timestamp 1621261055
transform 1 0 56064 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_576
timestamp 1621261055
transform 1 0 56448 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_579
timestamp 1621261055
transform 1 0 56736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_587
timestamp 1621261055
transform 1 0 57504 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_101
timestamp 1621261055
transform -1 0 58848 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_595
timestamp 1621261055
transform 1 0 58272 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_102
timestamp 1621261055
transform 1 0 1152 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_4
timestamp 1621261055
transform 1 0 1536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_12
timestamp 1621261055
transform 1 0 2304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_20
timestamp 1621261055
transform 1 0 3072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_28
timestamp 1621261055
transform 1 0 3840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_36
timestamp 1621261055
transform 1 0 4608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_710
timestamp 1621261055
transform 1 0 6432 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_44
timestamp 1621261055
transform 1 0 5376 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_52
timestamp 1621261055
transform 1 0 6144 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_54
timestamp 1621261055
transform 1 0 6336 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_56
timestamp 1621261055
transform 1 0 6528 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_64
timestamp 1621261055
transform 1 0 7296 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_72
timestamp 1621261055
transform 1 0 8064 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_80
timestamp 1621261055
transform 1 0 8832 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_88
timestamp 1621261055
transform 1 0 9600 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_96
timestamp 1621261055
transform 1 0 10368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_104
timestamp 1621261055
transform 1 0 11136 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_711
timestamp 1621261055
transform 1 0 11712 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_108
timestamp 1621261055
transform 1 0 11520 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_111
timestamp 1621261055
transform 1 0 11808 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_119
timestamp 1621261055
transform 1 0 12576 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _109_
timestamp 1621261055
transform 1 0 14688 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_182
timestamp 1621261055
transform 1 0 14496 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_127
timestamp 1621261055
transform 1 0 13344 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_135
timestamp 1621261055
transform 1 0 14112 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_144
timestamp 1621261055
transform 1 0 14976 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_712
timestamp 1621261055
transform 1 0 16992 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_152
timestamp 1621261055
transform 1 0 15744 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_160
timestamp 1621261055
transform 1 0 16512 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_51_164
timestamp 1621261055
transform 1 0 16896 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_166
timestamp 1621261055
transform 1 0 17088 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_174
timestamp 1621261055
transform 1 0 17856 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_182
timestamp 1621261055
transform 1 0 18624 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_190
timestamp 1621261055
transform 1 0 19392 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_198
timestamp 1621261055
transform 1 0 20160 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_206
timestamp 1621261055
transform 1 0 20928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_713
timestamp 1621261055
transform 1 0 22272 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_214
timestamp 1621261055
transform 1 0 21696 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_218
timestamp 1621261055
transform 1 0 22080 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_221
timestamp 1621261055
transform 1 0 22368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_229
timestamp 1621261055
transform 1 0 23136 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _070_
timestamp 1621261055
transform -1 0 24288 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_130
timestamp 1621261055
transform -1 0 24000 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_233
timestamp 1621261055
transform 1 0 23520 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_235
timestamp 1621261055
transform 1 0 23712 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_241
timestamp 1621261055
transform 1 0 24288 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_249
timestamp 1621261055
transform 1 0 25056 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_257
timestamp 1621261055
transform 1 0 25824 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_265
timestamp 1621261055
transform 1 0 26592 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_273
timestamp 1621261055
transform 1 0 27360 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_714
timestamp 1621261055
transform 1 0 27552 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_276
timestamp 1621261055
transform 1 0 27648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_284
timestamp 1621261055
transform 1 0 28416 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_292
timestamp 1621261055
transform 1 0 29184 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_300
timestamp 1621261055
transform 1 0 29952 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_308
timestamp 1621261055
transform 1 0 30720 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_715
timestamp 1621261055
transform 1 0 32832 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_316
timestamp 1621261055
transform 1 0 31488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_324
timestamp 1621261055
transform 1 0 32256 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_328
timestamp 1621261055
transform 1 0 32640 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_331
timestamp 1621261055
transform 1 0 32928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_339
timestamp 1621261055
transform 1 0 33696 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_347
timestamp 1621261055
transform 1 0 34464 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_355
timestamp 1621261055
transform 1 0 35232 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_363
timestamp 1621261055
transform 1 0 36000 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_371
timestamp 1621261055
transform 1 0 36768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_716
timestamp 1621261055
transform 1 0 38112 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_379
timestamp 1621261055
transform 1 0 37536 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_383
timestamp 1621261055
transform 1 0 37920 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_386
timestamp 1621261055
transform 1 0 38208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_394
timestamp 1621261055
transform 1 0 38976 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_402
timestamp 1621261055
transform 1 0 39744 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_410
timestamp 1621261055
transform 1 0 40512 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_418
timestamp 1621261055
transform 1 0 41280 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_717
timestamp 1621261055
transform 1 0 43392 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_426
timestamp 1621261055
transform 1 0 42048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_434
timestamp 1621261055
transform 1 0 42816 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_438
timestamp 1621261055
transform 1 0 43200 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_441
timestamp 1621261055
transform 1 0 43488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_449
timestamp 1621261055
transform 1 0 44256 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_457
timestamp 1621261055
transform 1 0 45024 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_465
timestamp 1621261055
transform 1 0 45792 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_473
timestamp 1621261055
transform 1 0 46560 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_481
timestamp 1621261055
transform 1 0 47328 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_718
timestamp 1621261055
transform 1 0 48672 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_489
timestamp 1621261055
transform 1 0 48096 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_493
timestamp 1621261055
transform 1 0 48480 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_496
timestamp 1621261055
transform 1 0 48768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_504
timestamp 1621261055
transform 1 0 49536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_512
timestamp 1621261055
transform 1 0 50304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_520
timestamp 1621261055
transform 1 0 51072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_528
timestamp 1621261055
transform 1 0 51840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_536
timestamp 1621261055
transform 1 0 52608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_544
timestamp 1621261055
transform 1 0 53376 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_719
timestamp 1621261055
transform 1 0 53952 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_548
timestamp 1621261055
transform 1 0 53760 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_551
timestamp 1621261055
transform 1 0 54048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_559
timestamp 1621261055
transform 1 0 54816 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_567
timestamp 1621261055
transform 1 0 55584 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_575
timestamp 1621261055
transform 1 0 56352 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_583
timestamp 1621261055
transform 1 0 57120 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_103
timestamp 1621261055
transform -1 0 58848 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_51_591
timestamp 1621261055
transform 1 0 57888 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_595
timestamp 1621261055
transform 1 0 58272 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_104
timestamp 1621261055
transform 1 0 1152 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_52_4
timestamp 1621261055
transform 1 0 1536 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_12
timestamp 1621261055
transform 1 0 2304 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_20
timestamp 1621261055
transform 1 0 3072 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _032_
timestamp 1621261055
transform 1 0 4800 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_720
timestamp 1621261055
transform 1 0 3840 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_29
timestamp 1621261055
transform 1 0 3936 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_52_37
timestamp 1621261055
transform 1 0 4704 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_41
timestamp 1621261055
transform 1 0 5088 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _063_
timestamp 1621261055
transform 1 0 5856 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_185
timestamp 1621261055
transform 1 0 5664 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_45
timestamp 1621261055
transform 1 0 5472 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_52
timestamp 1621261055
transform 1 0 6144 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_60
timestamp 1621261055
transform 1 0 6912 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_721
timestamp 1621261055
transform 1 0 9120 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_68
timestamp 1621261055
transform 1 0 7680 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_76
timestamp 1621261055
transform 1 0 8448 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_80
timestamp 1621261055
transform 1 0 8832 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_82
timestamp 1621261055
transform 1 0 9024 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_84
timestamp 1621261055
transform 1 0 9216 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_92
timestamp 1621261055
transform 1 0 9984 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_100
timestamp 1621261055
transform 1 0 10752 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_108
timestamp 1621261055
transform 1 0 11520 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_116
timestamp 1621261055
transform 1 0 12288 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_124
timestamp 1621261055
transform 1 0 13056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_722
timestamp 1621261055
transform 1 0 14400 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_132
timestamp 1621261055
transform 1 0 13824 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_136
timestamp 1621261055
transform 1 0 14208 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_139
timestamp 1621261055
transform 1 0 14496 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_147
timestamp 1621261055
transform 1 0 15264 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_155
timestamp 1621261055
transform 1 0 16032 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_163
timestamp 1621261055
transform 1 0 16800 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_171
timestamp 1621261055
transform 1 0 17568 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_179
timestamp 1621261055
transform 1 0 18336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_187
timestamp 1621261055
transform 1 0 19104 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_723
timestamp 1621261055
transform 1 0 19680 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_191
timestamp 1621261055
transform 1 0 19488 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_194
timestamp 1621261055
transform 1 0 19776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_202
timestamp 1621261055
transform 1 0 20544 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_210
timestamp 1621261055
transform 1 0 21312 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_218
timestamp 1621261055
transform 1 0 22080 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_226
timestamp 1621261055
transform 1 0 22848 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_724
timestamp 1621261055
transform 1 0 24960 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_234
timestamp 1621261055
transform 1 0 23616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_242
timestamp 1621261055
transform 1 0 24384 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_246
timestamp 1621261055
transform 1 0 24768 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_249
timestamp 1621261055
transform 1 0 25056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_257
timestamp 1621261055
transform 1 0 25824 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_265
timestamp 1621261055
transform 1 0 26592 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_273
timestamp 1621261055
transform 1 0 27360 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_281
timestamp 1621261055
transform 1 0 28128 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_289
timestamp 1621261055
transform 1 0 28896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_725
timestamp 1621261055
transform 1 0 30240 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_297
timestamp 1621261055
transform 1 0 29664 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_301
timestamp 1621261055
transform 1 0 30048 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_304
timestamp 1621261055
transform 1 0 30336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_312
timestamp 1621261055
transform 1 0 31104 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_320
timestamp 1621261055
transform 1 0 31872 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_328
timestamp 1621261055
transform 1 0 32640 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_336
timestamp 1621261055
transform 1 0 33408 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_344
timestamp 1621261055
transform 1 0 34176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_352
timestamp 1621261055
transform 1 0 34944 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_356
timestamp 1621261055
transform 1 0 35328 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_726
timestamp 1621261055
transform 1 0 35520 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_359
timestamp 1621261055
transform 1 0 35616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_367
timestamp 1621261055
transform 1 0 36384 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_375
timestamp 1621261055
transform 1 0 37152 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_383
timestamp 1621261055
transform 1 0 37920 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_391
timestamp 1621261055
transform 1 0 38688 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_399
timestamp 1621261055
transform 1 0 39456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_727
timestamp 1621261055
transform 1 0 40800 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_407
timestamp 1621261055
transform 1 0 40224 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_411
timestamp 1621261055
transform 1 0 40608 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_414
timestamp 1621261055
transform 1 0 40896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _028_
timestamp 1621261055
transform 1 0 43104 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_52_422
timestamp 1621261055
transform 1 0 41664 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_430
timestamp 1621261055
transform 1 0 42432 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_434
timestamp 1621261055
transform 1 0 42816 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_436
timestamp 1621261055
transform 1 0 43008 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_440
timestamp 1621261055
transform 1 0 43392 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_448
timestamp 1621261055
transform 1 0 44160 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_456
timestamp 1621261055
transform 1 0 44928 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_728
timestamp 1621261055
transform 1 0 46080 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_464
timestamp 1621261055
transform 1 0 45696 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_52_469
timestamp 1621261055
transform 1 0 46176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_477
timestamp 1621261055
transform 1 0 46944 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_485
timestamp 1621261055
transform 1 0 47712 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_493
timestamp 1621261055
transform 1 0 48480 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_501
timestamp 1621261055
transform 1 0 49248 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_729
timestamp 1621261055
transform 1 0 51360 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_509
timestamp 1621261055
transform 1 0 50016 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_517
timestamp 1621261055
transform 1 0 50784 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_521
timestamp 1621261055
transform 1 0 51168 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_524
timestamp 1621261055
transform 1 0 51456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_532
timestamp 1621261055
transform 1 0 52224 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_540
timestamp 1621261055
transform 1 0 52992 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_548
timestamp 1621261055
transform 1 0 53760 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_556
timestamp 1621261055
transform 1 0 54528 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_564
timestamp 1621261055
transform 1 0 55296 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_730
timestamp 1621261055
transform 1 0 56640 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_572
timestamp 1621261055
transform 1 0 56064 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_576
timestamp 1621261055
transform 1 0 56448 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_579
timestamp 1621261055
transform 1 0 56736 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_587
timestamp 1621261055
transform 1 0 57504 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_105
timestamp 1621261055
transform -1 0 58848 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_595
timestamp 1621261055
transform 1 0 58272 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_106
timestamp 1621261055
transform 1 0 1152 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_4
timestamp 1621261055
transform 1 0 1536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_12
timestamp 1621261055
transform 1 0 2304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_20
timestamp 1621261055
transform 1 0 3072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_28
timestamp 1621261055
transform 1 0 3840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_36
timestamp 1621261055
transform 1 0 4608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_731
timestamp 1621261055
transform 1 0 6432 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_44
timestamp 1621261055
transform 1 0 5376 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_52
timestamp 1621261055
transform 1 0 6144 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_54
timestamp 1621261055
transform 1 0 6336 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_56
timestamp 1621261055
transform 1 0 6528 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_64
timestamp 1621261055
transform 1 0 7296 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_72
timestamp 1621261055
transform 1 0 8064 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_80
timestamp 1621261055
transform 1 0 8832 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_88
timestamp 1621261055
transform 1 0 9600 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_96
timestamp 1621261055
transform 1 0 10368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_104
timestamp 1621261055
transform 1 0 11136 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_732
timestamp 1621261055
transform 1 0 11712 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_108
timestamp 1621261055
transform 1 0 11520 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_111
timestamp 1621261055
transform 1 0 11808 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_119
timestamp 1621261055
transform 1 0 12576 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_127
timestamp 1621261055
transform 1 0 13344 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_135
timestamp 1621261055
transform 1 0 14112 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_143
timestamp 1621261055
transform 1 0 14880 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_733
timestamp 1621261055
transform 1 0 16992 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_151
timestamp 1621261055
transform 1 0 15648 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_159
timestamp 1621261055
transform 1 0 16416 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_163
timestamp 1621261055
transform 1 0 16800 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_166
timestamp 1621261055
transform 1 0 17088 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_174
timestamp 1621261055
transform 1 0 17856 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_182
timestamp 1621261055
transform 1 0 18624 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_190
timestamp 1621261055
transform 1 0 19392 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_198
timestamp 1621261055
transform 1 0 20160 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_206
timestamp 1621261055
transform 1 0 20928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_734
timestamp 1621261055
transform 1 0 22272 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_214
timestamp 1621261055
transform 1 0 21696 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_218
timestamp 1621261055
transform 1 0 22080 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_221
timestamp 1621261055
transform 1 0 22368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_229
timestamp 1621261055
transform 1 0 23136 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_237
timestamp 1621261055
transform 1 0 23904 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_245
timestamp 1621261055
transform 1 0 24672 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_253
timestamp 1621261055
transform 1 0 25440 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_261
timestamp 1621261055
transform 1 0 26208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_269
timestamp 1621261055
transform 1 0 26976 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_273
timestamp 1621261055
transform 1 0 27360 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_735
timestamp 1621261055
transform 1 0 27552 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_276
timestamp 1621261055
transform 1 0 27648 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_284
timestamp 1621261055
transform 1 0 28416 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_292
timestamp 1621261055
transform 1 0 29184 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_300
timestamp 1621261055
transform 1 0 29952 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_308
timestamp 1621261055
transform 1 0 30720 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_736
timestamp 1621261055
transform 1 0 32832 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_316
timestamp 1621261055
transform 1 0 31488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_324
timestamp 1621261055
transform 1 0 32256 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_328
timestamp 1621261055
transform 1 0 32640 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_331
timestamp 1621261055
transform 1 0 32928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _097_
timestamp 1621261055
transform -1 0 34656 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_170
timestamp 1621261055
transform -1 0 34368 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_53_339
timestamp 1621261055
transform 1 0 33696 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_53_343
timestamp 1621261055
transform 1 0 34080 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_349
timestamp 1621261055
transform 1 0 34656 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_357
timestamp 1621261055
transform 1 0 35424 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_365
timestamp 1621261055
transform 1 0 36192 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_373
timestamp 1621261055
transform 1 0 36960 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_737
timestamp 1621261055
transform 1 0 38112 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_381
timestamp 1621261055
transform 1 0 37728 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_386
timestamp 1621261055
transform 1 0 38208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_394
timestamp 1621261055
transform 1 0 38976 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_402
timestamp 1621261055
transform 1 0 39744 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_410
timestamp 1621261055
transform 1 0 40512 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_418
timestamp 1621261055
transform 1 0 41280 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_738
timestamp 1621261055
transform 1 0 43392 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_426
timestamp 1621261055
transform 1 0 42048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_434
timestamp 1621261055
transform 1 0 42816 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_438
timestamp 1621261055
transform 1 0 43200 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_441
timestamp 1621261055
transform 1 0 43488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_449
timestamp 1621261055
transform 1 0 44256 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_457
timestamp 1621261055
transform 1 0 45024 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_465
timestamp 1621261055
transform 1 0 45792 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_473
timestamp 1621261055
transform 1 0 46560 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_481
timestamp 1621261055
transform 1 0 47328 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_739
timestamp 1621261055
transform 1 0 48672 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_489
timestamp 1621261055
transform 1 0 48096 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_493
timestamp 1621261055
transform 1 0 48480 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_496
timestamp 1621261055
transform 1 0 48768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_504
timestamp 1621261055
transform 1 0 49536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_512
timestamp 1621261055
transform 1 0 50304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_520
timestamp 1621261055
transform 1 0 51072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_528
timestamp 1621261055
transform 1 0 51840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_536
timestamp 1621261055
transform 1 0 52608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_544
timestamp 1621261055
transform 1 0 53376 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _039_
timestamp 1621261055
transform 1 0 54432 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _198_
timestamp 1621261055
transform -1 0 55680 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_740
timestamp 1621261055
transform 1 0 53952 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_215
timestamp 1621261055
transform -1 0 55392 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_548
timestamp 1621261055
transform 1 0 53760 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_53_551
timestamp 1621261055
transform 1 0 54048 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_53_558
timestamp 1621261055
transform 1 0 54720 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_53_562
timestamp 1621261055
transform 1 0 55104 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_568
timestamp 1621261055
transform 1 0 55680 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_576
timestamp 1621261055
transform 1 0 56448 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_584
timestamp 1621261055
transform 1 0 57216 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_107
timestamp 1621261055
transform -1 0 58848 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_53_592
timestamp 1621261055
transform 1 0 57984 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_53_596
timestamp 1621261055
transform 1 0 58368 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_108
timestamp 1621261055
transform 1 0 1152 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_110
timestamp 1621261055
transform 1 0 1152 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_4
timestamp 1621261055
transform 1 0 1536 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_12
timestamp 1621261055
transform 1 0 2304 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_20
timestamp 1621261055
transform 1 0 3072 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_4
timestamp 1621261055
transform 1 0 1536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_12
timestamp 1621261055
transform 1 0 2304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_20
timestamp 1621261055
transform 1 0 3072 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_741
timestamp 1621261055
transform 1 0 3840 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_29
timestamp 1621261055
transform 1 0 3936 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_37
timestamp 1621261055
transform 1 0 4704 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_28
timestamp 1621261055
transform 1 0 3840 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_36
timestamp 1621261055
transform 1 0 4608 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_752
timestamp 1621261055
transform 1 0 6432 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_45
timestamp 1621261055
transform 1 0 5472 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_53
timestamp 1621261055
transform 1 0 6240 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_61
timestamp 1621261055
transform 1 0 7008 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_44
timestamp 1621261055
transform 1 0 5376 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_52
timestamp 1621261055
transform 1 0 6144 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_55_54
timestamp 1621261055
transform 1 0 6336 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_56
timestamp 1621261055
transform 1 0 6528 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_742
timestamp 1621261055
transform 1 0 9120 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_69
timestamp 1621261055
transform 1 0 7776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_77
timestamp 1621261055
transform 1 0 8544 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_81
timestamp 1621261055
transform 1 0 8928 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_84
timestamp 1621261055
transform 1 0 9216 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_64
timestamp 1621261055
transform 1 0 7296 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_72
timestamp 1621261055
transform 1 0 8064 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_80
timestamp 1621261055
transform 1 0 8832 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _088_
timestamp 1621261055
transform 1 0 10464 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_154
timestamp 1621261055
transform 1 0 10272 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_92
timestamp 1621261055
transform 1 0 9984 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_54_94
timestamp 1621261055
transform 1 0 10176 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_100
timestamp 1621261055
transform 1 0 10752 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_88
timestamp 1621261055
transform 1 0 9600 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_96
timestamp 1621261055
transform 1 0 10368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_104
timestamp 1621261055
transform 1 0 11136 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_753
timestamp 1621261055
transform 1 0 11712 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_108
timestamp 1621261055
transform 1 0 11520 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_116
timestamp 1621261055
transform 1 0 12288 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_124
timestamp 1621261055
transform 1 0 13056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_108
timestamp 1621261055
transform 1 0 11520 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_111
timestamp 1621261055
transform 1 0 11808 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_119
timestamp 1621261055
transform 1 0 12576 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_743
timestamp 1621261055
transform 1 0 14400 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_132
timestamp 1621261055
transform 1 0 13824 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_136
timestamp 1621261055
transform 1 0 14208 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_139
timestamp 1621261055
transform 1 0 14496 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_147
timestamp 1621261055
transform 1 0 15264 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_127
timestamp 1621261055
transform 1 0 13344 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_135
timestamp 1621261055
transform 1 0 14112 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_143
timestamp 1621261055
transform 1 0 14880 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_754
timestamp 1621261055
transform 1 0 16992 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_155
timestamp 1621261055
transform 1 0 16032 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_163
timestamp 1621261055
transform 1 0 16800 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_151
timestamp 1621261055
transform 1 0 15648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_159
timestamp 1621261055
transform 1 0 16416 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_163
timestamp 1621261055
transform 1 0 16800 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_166
timestamp 1621261055
transform 1 0 17088 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_171
timestamp 1621261055
transform 1 0 17568 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_179
timestamp 1621261055
transform 1 0 18336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_187
timestamp 1621261055
transform 1 0 19104 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_174
timestamp 1621261055
transform 1 0 17856 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_182
timestamp 1621261055
transform 1 0 18624 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_744
timestamp 1621261055
transform 1 0 19680 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_191
timestamp 1621261055
transform 1 0 19488 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_194
timestamp 1621261055
transform 1 0 19776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_202
timestamp 1621261055
transform 1 0 20544 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_210
timestamp 1621261055
transform 1 0 21312 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_190
timestamp 1621261055
transform 1 0 19392 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_198
timestamp 1621261055
transform 1 0 20160 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_206
timestamp 1621261055
transform 1 0 20928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_755
timestamp 1621261055
transform 1 0 22272 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_218
timestamp 1621261055
transform 1 0 22080 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_226
timestamp 1621261055
transform 1 0 22848 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_214
timestamp 1621261055
transform 1 0 21696 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_218
timestamp 1621261055
transform 1 0 22080 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_221
timestamp 1621261055
transform 1 0 22368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_229
timestamp 1621261055
transform 1 0 23136 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _104_
timestamp 1621261055
transform 1 0 24192 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_745
timestamp 1621261055
transform 1 0 24960 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_176
timestamp 1621261055
transform 1 0 24000 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_234
timestamp 1621261055
transform 1 0 23616 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_54_243
timestamp 1621261055
transform 1 0 24480 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_54_247
timestamp 1621261055
transform 1 0 24864 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_249
timestamp 1621261055
transform 1 0 25056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_237
timestamp 1621261055
transform 1 0 23904 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_245
timestamp 1621261055
transform 1 0 24672 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _017_
timestamp 1621261055
transform 1 0 26592 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_54_257
timestamp 1621261055
transform 1 0 25824 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_268
timestamp 1621261055
transform 1 0 26880 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_253
timestamp 1621261055
transform 1 0 25440 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_261
timestamp 1621261055
transform 1 0 26208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_269
timestamp 1621261055
transform 1 0 26976 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_273
timestamp 1621261055
transform 1 0 27360 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_756
timestamp 1621261055
transform 1 0 27552 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_276
timestamp 1621261055
transform 1 0 27648 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_284
timestamp 1621261055
transform 1 0 28416 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_292
timestamp 1621261055
transform 1 0 29184 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_276
timestamp 1621261055
transform 1 0 27648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_284
timestamp 1621261055
transform 1 0 28416 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_292
timestamp 1621261055
transform 1 0 29184 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_300
timestamp 1621261055
transform 1 0 29952 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_302
timestamp 1621261055
transform 1 0 30144 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_300
timestamp 1621261055
transform 1 0 29952 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_308
timestamp 1621261055
transform 1 0 30720 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_311
timestamp 1621261055
transform 1 0 31008 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_304
timestamp 1621261055
transform 1 0 30336 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_746
timestamp 1621261055
transform 1 0 30240 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _003_
timestamp 1621261055
transform 1 0 30720 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_188
timestamp 1621261055
transform 1 0 31200 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _122_
timestamp 1621261055
transform 1 0 31392 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_757
timestamp 1621261055
transform 1 0 32832 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_318
timestamp 1621261055
transform 1 0 31680 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_326
timestamp 1621261055
transform 1 0 32448 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_334
timestamp 1621261055
transform 1 0 33216 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_316
timestamp 1621261055
transform 1 0 31488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_324
timestamp 1621261055
transform 1 0 32256 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_328
timestamp 1621261055
transform 1 0 32640 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_331
timestamp 1621261055
transform 1 0 32928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_342
timestamp 1621261055
transform 1 0 33984 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_350
timestamp 1621261055
transform 1 0 34752 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_339
timestamp 1621261055
transform 1 0 33696 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_347
timestamp 1621261055
transform 1 0 34464 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_355
timestamp 1621261055
transform 1 0 35232 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_747
timestamp 1621261055
transform 1 0 35520 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_359
timestamp 1621261055
transform 1 0 35616 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_367
timestamp 1621261055
transform 1 0 36384 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_375
timestamp 1621261055
transform 1 0 37152 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_363
timestamp 1621261055
transform 1 0 36000 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_371
timestamp 1621261055
transform 1 0 36768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_758
timestamp 1621261055
transform 1 0 38112 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_383
timestamp 1621261055
transform 1 0 37920 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_391
timestamp 1621261055
transform 1 0 38688 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_399
timestamp 1621261055
transform 1 0 39456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_379
timestamp 1621261055
transform 1 0 37536 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_383
timestamp 1621261055
transform 1 0 37920 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_386
timestamp 1621261055
transform 1 0 38208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_394
timestamp 1621261055
transform 1 0 38976 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_748
timestamp 1621261055
transform 1 0 40800 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_407
timestamp 1621261055
transform 1 0 40224 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_411
timestamp 1621261055
transform 1 0 40608 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_414
timestamp 1621261055
transform 1 0 40896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_402
timestamp 1621261055
transform 1 0 39744 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_410
timestamp 1621261055
transform 1 0 40512 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_418
timestamp 1621261055
transform 1 0 41280 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_759
timestamp 1621261055
transform 1 0 43392 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_422
timestamp 1621261055
transform 1 0 41664 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_430
timestamp 1621261055
transform 1 0 42432 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_438
timestamp 1621261055
transform 1 0 43200 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_426
timestamp 1621261055
transform 1 0 42048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_434
timestamp 1621261055
transform 1 0 42816 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_438
timestamp 1621261055
transform 1 0 43200 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_441
timestamp 1621261055
transform 1 0 43488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_446
timestamp 1621261055
transform 1 0 43968 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_454
timestamp 1621261055
transform 1 0 44736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_462
timestamp 1621261055
transform 1 0 45504 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_449
timestamp 1621261055
transform 1 0 44256 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_457
timestamp 1621261055
transform 1 0 45024 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_749
timestamp 1621261055
transform 1 0 46080 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_466
timestamp 1621261055
transform 1 0 45888 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_469
timestamp 1621261055
transform 1 0 46176 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_477
timestamp 1621261055
transform 1 0 46944 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_465
timestamp 1621261055
transform 1 0 45792 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_473
timestamp 1621261055
transform 1 0 46560 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_481
timestamp 1621261055
transform 1 0 47328 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_760
timestamp 1621261055
transform 1 0 48672 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_485
timestamp 1621261055
transform 1 0 47712 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_493
timestamp 1621261055
transform 1 0 48480 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_501
timestamp 1621261055
transform 1 0 49248 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_489
timestamp 1621261055
transform 1 0 48096 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_493
timestamp 1621261055
transform 1 0 48480 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_496
timestamp 1621261055
transform 1 0 48768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_504
timestamp 1621261055
transform 1 0 49536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_750
timestamp 1621261055
transform 1 0 51360 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_509
timestamp 1621261055
transform 1 0 50016 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_517
timestamp 1621261055
transform 1 0 50784 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_521
timestamp 1621261055
transform 1 0 51168 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_524
timestamp 1621261055
transform 1 0 51456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_512
timestamp 1621261055
transform 1 0 50304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_520
timestamp 1621261055
transform 1 0 51072 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_532
timestamp 1621261055
transform 1 0 52224 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_540
timestamp 1621261055
transform 1 0 52992 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_528
timestamp 1621261055
transform 1 0 51840 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_536
timestamp 1621261055
transform 1 0 52608 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_544
timestamp 1621261055
transform 1 0 53376 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_761
timestamp 1621261055
transform 1 0 53952 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_548
timestamp 1621261055
transform 1 0 53760 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_556
timestamp 1621261055
transform 1 0 54528 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_564
timestamp 1621261055
transform 1 0 55296 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_548
timestamp 1621261055
transform 1 0 53760 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_551
timestamp 1621261055
transform 1 0 54048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_559
timestamp 1621261055
transform 1 0 54816 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_567
timestamp 1621261055
transform 1 0 55584 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_575
timestamp 1621261055
transform 1 0 56352 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_576
timestamp 1621261055
transform 1 0 56448 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_572
timestamp 1621261055
transform 1 0 56064 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_55_583
timestamp 1621261055
transform 1 0 57120 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_579
timestamp 1621261055
transform 1 0 56736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_751
timestamp 1621261055
transform 1 0 56640 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_55_587
timestamp 1621261055
transform 1 0 57504 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_54_587
timestamp 1621261055
transform 1 0 57504 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_208
timestamp 1621261055
transform -1 0 57792 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_118
timestamp 1621261055
transform -1 0 57792 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _149_
timestamp 1621261055
transform -1 0 58080 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _177_
timestamp 1621261055
transform -1 0 58080 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_109
timestamp 1621261055
transform -1 0 58848 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_111
timestamp 1621261055
transform -1 0 58848 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_54_593
timestamp 1621261055
transform 1 0 58080 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_55_593
timestamp 1621261055
transform 1 0 58080 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_112
timestamp 1621261055
transform 1 0 1152 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_56_4
timestamp 1621261055
transform 1 0 1536 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_12
timestamp 1621261055
transform 1 0 2304 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_20
timestamp 1621261055
transform 1 0 3072 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_762
timestamp 1621261055
transform 1 0 3840 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_29
timestamp 1621261055
transform 1 0 3936 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_37
timestamp 1621261055
transform 1 0 4704 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_45
timestamp 1621261055
transform 1 0 5472 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_53
timestamp 1621261055
transform 1 0 6240 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_61
timestamp 1621261055
transform 1 0 7008 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_763
timestamp 1621261055
transform 1 0 9120 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_69
timestamp 1621261055
transform 1 0 7776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_77
timestamp 1621261055
transform 1 0 8544 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_81
timestamp 1621261055
transform 1 0 8928 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_84
timestamp 1621261055
transform 1 0 9216 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_92
timestamp 1621261055
transform 1 0 9984 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_100
timestamp 1621261055
transform 1 0 10752 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_108
timestamp 1621261055
transform 1 0 11520 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_116
timestamp 1621261055
transform 1 0 12288 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_124
timestamp 1621261055
transform 1 0 13056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_764
timestamp 1621261055
transform 1 0 14400 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_132
timestamp 1621261055
transform 1 0 13824 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_136
timestamp 1621261055
transform 1 0 14208 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_139
timestamp 1621261055
transform 1 0 14496 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_147
timestamp 1621261055
transform 1 0 15264 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_155
timestamp 1621261055
transform 1 0 16032 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_163
timestamp 1621261055
transform 1 0 16800 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_171
timestamp 1621261055
transform 1 0 17568 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_179
timestamp 1621261055
transform 1 0 18336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_187
timestamp 1621261055
transform 1 0 19104 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_765
timestamp 1621261055
transform 1 0 19680 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_191
timestamp 1621261055
transform 1 0 19488 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_194
timestamp 1621261055
transform 1 0 19776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_202
timestamp 1621261055
transform 1 0 20544 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_210
timestamp 1621261055
transform 1 0 21312 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_218
timestamp 1621261055
transform 1 0 22080 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_226
timestamp 1621261055
transform 1 0 22848 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_766
timestamp 1621261055
transform 1 0 24960 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_234
timestamp 1621261055
transform 1 0 23616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_242
timestamp 1621261055
transform 1 0 24384 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_246
timestamp 1621261055
transform 1 0 24768 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_249
timestamp 1621261055
transform 1 0 25056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _090_
timestamp 1621261055
transform -1 0 27072 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_158
timestamp 1621261055
transform -1 0 26784 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_257
timestamp 1621261055
transform 1 0 25824 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_270
timestamp 1621261055
transform 1 0 27072 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_278
timestamp 1621261055
transform 1 0 27840 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_286
timestamp 1621261055
transform 1 0 28608 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_294
timestamp 1621261055
transform 1 0 29376 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_767
timestamp 1621261055
transform 1 0 30240 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_56_302
timestamp 1621261055
transform 1 0 30144 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_304
timestamp 1621261055
transform 1 0 30336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_312
timestamp 1621261055
transform 1 0 31104 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_320
timestamp 1621261055
transform 1 0 31872 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_328
timestamp 1621261055
transform 1 0 32640 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_336
timestamp 1621261055
transform 1 0 33408 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_344
timestamp 1621261055
transform 1 0 34176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_352
timestamp 1621261055
transform 1 0 34944 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_356
timestamp 1621261055
transform 1 0 35328 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_768
timestamp 1621261055
transform 1 0 35520 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_359
timestamp 1621261055
transform 1 0 35616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_367
timestamp 1621261055
transform 1 0 36384 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_375
timestamp 1621261055
transform 1 0 37152 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_383
timestamp 1621261055
transform 1 0 37920 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_391
timestamp 1621261055
transform 1 0 38688 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_399
timestamp 1621261055
transform 1 0 39456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_769
timestamp 1621261055
transform 1 0 40800 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_407
timestamp 1621261055
transform 1 0 40224 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_411
timestamp 1621261055
transform 1 0 40608 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_414
timestamp 1621261055
transform 1 0 40896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_422
timestamp 1621261055
transform 1 0 41664 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_430
timestamp 1621261055
transform 1 0 42432 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_438
timestamp 1621261055
transform 1 0 43200 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _012_
timestamp 1621261055
transform 1 0 44928 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_56_446
timestamp 1621261055
transform 1 0 43968 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_454
timestamp 1621261055
transform 1 0 44736 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_459
timestamp 1621261055
transform 1 0 45216 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_770
timestamp 1621261055
transform 1 0 46080 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_56_467
timestamp 1621261055
transform 1 0 45984 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_469
timestamp 1621261055
transform 1 0 46176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_477
timestamp 1621261055
transform 1 0 46944 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_485
timestamp 1621261055
transform 1 0 47712 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_493
timestamp 1621261055
transform 1 0 48480 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_501
timestamp 1621261055
transform 1 0 49248 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_771
timestamp 1621261055
transform 1 0 51360 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_509
timestamp 1621261055
transform 1 0 50016 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_517
timestamp 1621261055
transform 1 0 50784 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_521
timestamp 1621261055
transform 1 0 51168 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_524
timestamp 1621261055
transform 1 0 51456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_532
timestamp 1621261055
transform 1 0 52224 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_540
timestamp 1621261055
transform 1 0 52992 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_548
timestamp 1621261055
transform 1 0 53760 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_556
timestamp 1621261055
transform 1 0 54528 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_564
timestamp 1621261055
transform 1 0 55296 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _072_
timestamp 1621261055
transform -1 0 57792 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_772
timestamp 1621261055
transform 1 0 56640 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_134
timestamp 1621261055
transform -1 0 57504 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_56_572
timestamp 1621261055
transform 1 0 56064 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_576
timestamp 1621261055
transform 1 0 56448 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_56_579
timestamp 1621261055
transform 1 0 56736 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_583
timestamp 1621261055
transform 1 0 57120 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_113
timestamp 1621261055
transform -1 0 58848 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_56_590
timestamp 1621261055
transform 1 0 57792 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_594
timestamp 1621261055
transform 1 0 58176 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_56_596
timestamp 1621261055
transform 1 0 58368 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _102_
timestamp 1621261055
transform 1 0 1632 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_114
timestamp 1621261055
transform 1 0 1152 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_174
timestamp 1621261055
transform 1 0 1920 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_4
timestamp 1621261055
transform 1 0 1536 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_10
timestamp 1621261055
transform 1 0 2112 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_18
timestamp 1621261055
transform 1 0 2880 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_26
timestamp 1621261055
transform 1 0 3648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_34
timestamp 1621261055
transform 1 0 4416 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_42
timestamp 1621261055
transform 1 0 5184 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_773
timestamp 1621261055
transform 1 0 6432 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_50
timestamp 1621261055
transform 1 0 5952 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_57_54
timestamp 1621261055
transform 1 0 6336 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_56
timestamp 1621261055
transform 1 0 6528 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_64
timestamp 1621261055
transform 1 0 7296 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_72
timestamp 1621261055
transform 1 0 8064 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_80
timestamp 1621261055
transform 1 0 8832 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_88
timestamp 1621261055
transform 1 0 9600 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_96
timestamp 1621261055
transform 1 0 10368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_104
timestamp 1621261055
transform 1 0 11136 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_774
timestamp 1621261055
transform 1 0 11712 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_108
timestamp 1621261055
transform 1 0 11520 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_111
timestamp 1621261055
transform 1 0 11808 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_119
timestamp 1621261055
transform 1 0 12576 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_127
timestamp 1621261055
transform 1 0 13344 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_135
timestamp 1621261055
transform 1 0 14112 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_143
timestamp 1621261055
transform 1 0 14880 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_775
timestamp 1621261055
transform 1 0 16992 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_151
timestamp 1621261055
transform 1 0 15648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_159
timestamp 1621261055
transform 1 0 16416 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_163
timestamp 1621261055
transform 1 0 16800 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_166
timestamp 1621261055
transform 1 0 17088 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_174
timestamp 1621261055
transform 1 0 17856 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_182
timestamp 1621261055
transform 1 0 18624 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_190
timestamp 1621261055
transform 1 0 19392 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_198
timestamp 1621261055
transform 1 0 20160 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_206
timestamp 1621261055
transform 1 0 20928 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_776
timestamp 1621261055
transform 1 0 22272 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_214
timestamp 1621261055
transform 1 0 21696 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_218
timestamp 1621261055
transform 1 0 22080 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_221
timestamp 1621261055
transform 1 0 22368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_229
timestamp 1621261055
transform 1 0 23136 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_237
timestamp 1621261055
transform 1 0 23904 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_245
timestamp 1621261055
transform 1 0 24672 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_253
timestamp 1621261055
transform 1 0 25440 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_261
timestamp 1621261055
transform 1 0 26208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_269
timestamp 1621261055
transform 1 0 26976 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_273
timestamp 1621261055
transform 1 0 27360 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_777
timestamp 1621261055
transform 1 0 27552 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_276
timestamp 1621261055
transform 1 0 27648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_284
timestamp 1621261055
transform 1 0 28416 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_292
timestamp 1621261055
transform 1 0 29184 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_300
timestamp 1621261055
transform 1 0 29952 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_308
timestamp 1621261055
transform 1 0 30720 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _150_
timestamp 1621261055
transform 1 0 33312 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_778
timestamp 1621261055
transform 1 0 32832 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_316
timestamp 1621261055
transform 1 0 31488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_324
timestamp 1621261055
transform 1 0 32256 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_328
timestamp 1621261055
transform 1 0 32640 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_57_331
timestamp 1621261055
transform 1 0 32928 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _195_
timestamp 1621261055
transform -1 0 34368 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_237
timestamp 1621261055
transform -1 0 34080 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_338
timestamp 1621261055
transform 1 0 33600 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_340
timestamp 1621261055
transform 1 0 33792 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_346
timestamp 1621261055
transform 1 0 34368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_354
timestamp 1621261055
transform 1 0 35136 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_362
timestamp 1621261055
transform 1 0 35904 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_370
timestamp 1621261055
transform 1 0 36672 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_378
timestamp 1621261055
transform 1 0 37440 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_779
timestamp 1621261055
transform 1 0 38112 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_382
timestamp 1621261055
transform 1 0 37824 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_384
timestamp 1621261055
transform 1 0 38016 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_386
timestamp 1621261055
transform 1 0 38208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_394
timestamp 1621261055
transform 1 0 38976 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_402
timestamp 1621261055
transform 1 0 39744 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_410
timestamp 1621261055
transform 1 0 40512 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_418
timestamp 1621261055
transform 1 0 41280 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_780
timestamp 1621261055
transform 1 0 43392 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_426
timestamp 1621261055
transform 1 0 42048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_434
timestamp 1621261055
transform 1 0 42816 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_438
timestamp 1621261055
transform 1 0 43200 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_441
timestamp 1621261055
transform 1 0 43488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_449
timestamp 1621261055
transform 1 0 44256 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_457
timestamp 1621261055
transform 1 0 45024 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_465
timestamp 1621261055
transform 1 0 45792 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_473
timestamp 1621261055
transform 1 0 46560 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_481
timestamp 1621261055
transform 1 0 47328 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_781
timestamp 1621261055
transform 1 0 48672 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_489
timestamp 1621261055
transform 1 0 48096 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_493
timestamp 1621261055
transform 1 0 48480 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_496
timestamp 1621261055
transform 1 0 48768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_504
timestamp 1621261055
transform 1 0 49536 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_512
timestamp 1621261055
transform 1 0 50304 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_520
timestamp 1621261055
transform 1 0 51072 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_528
timestamp 1621261055
transform 1 0 51840 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_536
timestamp 1621261055
transform 1 0 52608 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_544
timestamp 1621261055
transform 1 0 53376 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_782
timestamp 1621261055
transform 1 0 53952 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_548
timestamp 1621261055
transform 1 0 53760 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_551
timestamp 1621261055
transform 1 0 54048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_559
timestamp 1621261055
transform 1 0 54816 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_567
timestamp 1621261055
transform 1 0 55584 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_575
timestamp 1621261055
transform 1 0 56352 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_583
timestamp 1621261055
transform 1 0 57120 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_115
timestamp 1621261055
transform -1 0 58848 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_57_591
timestamp 1621261055
transform 1 0 57888 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_595
timestamp 1621261055
transform 1 0 58272 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_116
timestamp 1621261055
transform 1 0 1152 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_58_4
timestamp 1621261055
transform 1 0 1536 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_12
timestamp 1621261055
transform 1 0 2304 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_20
timestamp 1621261055
transform 1 0 3072 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_783
timestamp 1621261055
transform 1 0 3840 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_29
timestamp 1621261055
transform 1 0 3936 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_37
timestamp 1621261055
transform 1 0 4704 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_45
timestamp 1621261055
transform 1 0 5472 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_53
timestamp 1621261055
transform 1 0 6240 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_61
timestamp 1621261055
transform 1 0 7008 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_784
timestamp 1621261055
transform 1 0 9120 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_69
timestamp 1621261055
transform 1 0 7776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_77
timestamp 1621261055
transform 1 0 8544 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_81
timestamp 1621261055
transform 1 0 8928 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_84
timestamp 1621261055
transform 1 0 9216 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_92
timestamp 1621261055
transform 1 0 9984 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_100
timestamp 1621261055
transform 1 0 10752 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_108
timestamp 1621261055
transform 1 0 11520 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_116
timestamp 1621261055
transform 1 0 12288 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_124
timestamp 1621261055
transform 1 0 13056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_785
timestamp 1621261055
transform 1 0 14400 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_132
timestamp 1621261055
transform 1 0 13824 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_136
timestamp 1621261055
transform 1 0 14208 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_139
timestamp 1621261055
transform 1 0 14496 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_147
timestamp 1621261055
transform 1 0 15264 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_155
timestamp 1621261055
transform 1 0 16032 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_163
timestamp 1621261055
transform 1 0 16800 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_171
timestamp 1621261055
transform 1 0 17568 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_179
timestamp 1621261055
transform 1 0 18336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_187
timestamp 1621261055
transform 1 0 19104 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_786
timestamp 1621261055
transform 1 0 19680 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_191
timestamp 1621261055
transform 1 0 19488 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_194
timestamp 1621261055
transform 1 0 19776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_202
timestamp 1621261055
transform 1 0 20544 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_210
timestamp 1621261055
transform 1 0 21312 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_218
timestamp 1621261055
transform 1 0 22080 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_226
timestamp 1621261055
transform 1 0 22848 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_787
timestamp 1621261055
transform 1 0 24960 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_234
timestamp 1621261055
transform 1 0 23616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_242
timestamp 1621261055
transform 1 0 24384 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_246
timestamp 1621261055
transform 1 0 24768 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_249
timestamp 1621261055
transform 1 0 25056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_257
timestamp 1621261055
transform 1 0 25824 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_265
timestamp 1621261055
transform 1 0 26592 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_273
timestamp 1621261055
transform 1 0 27360 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_281
timestamp 1621261055
transform 1 0 28128 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_289
timestamp 1621261055
transform 1 0 28896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_788
timestamp 1621261055
transform 1 0 30240 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_297
timestamp 1621261055
transform 1 0 29664 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_301
timestamp 1621261055
transform 1 0 30048 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_304
timestamp 1621261055
transform 1 0 30336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_312
timestamp 1621261055
transform 1 0 31104 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _080_
timestamp 1621261055
transform -1 0 33696 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_140
timestamp 1621261055
transform -1 0 33408 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_320
timestamp 1621261055
transform 1 0 31872 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_328
timestamp 1621261055
transform 1 0 32640 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_332
timestamp 1621261055
transform 1 0 33024 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_339
timestamp 1621261055
transform 1 0 33696 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_347
timestamp 1621261055
transform 1 0 34464 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_355
timestamp 1621261055
transform 1 0 35232 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_357
timestamp 1621261055
transform 1 0 35424 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_789
timestamp 1621261055
transform 1 0 35520 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_359
timestamp 1621261055
transform 1 0 35616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_367
timestamp 1621261055
transform 1 0 36384 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_375
timestamp 1621261055
transform 1 0 37152 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _001_
timestamp 1621261055
transform 1 0 38976 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_58_383
timestamp 1621261055
transform 1 0 37920 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_391
timestamp 1621261055
transform 1 0 38688 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_393
timestamp 1621261055
transform 1 0 38880 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_397
timestamp 1621261055
transform 1 0 39264 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_790
timestamp 1621261055
transform 1 0 40800 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_405
timestamp 1621261055
transform 1 0 40032 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_414
timestamp 1621261055
transform 1 0 40896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_422
timestamp 1621261055
transform 1 0 41664 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_430
timestamp 1621261055
transform 1 0 42432 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_438
timestamp 1621261055
transform 1 0 43200 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_446
timestamp 1621261055
transform 1 0 43968 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_454
timestamp 1621261055
transform 1 0 44736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_462
timestamp 1621261055
transform 1 0 45504 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_791
timestamp 1621261055
transform 1 0 46080 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_466
timestamp 1621261055
transform 1 0 45888 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_469
timestamp 1621261055
transform 1 0 46176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_477
timestamp 1621261055
transform 1 0 46944 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_485
timestamp 1621261055
transform 1 0 47712 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_493
timestamp 1621261055
transform 1 0 48480 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_501
timestamp 1621261055
transform 1 0 49248 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_792
timestamp 1621261055
transform 1 0 51360 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_509
timestamp 1621261055
transform 1 0 50016 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_517
timestamp 1621261055
transform 1 0 50784 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_521
timestamp 1621261055
transform 1 0 51168 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_524
timestamp 1621261055
transform 1 0 51456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_532
timestamp 1621261055
transform 1 0 52224 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_540
timestamp 1621261055
transform 1 0 52992 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_548
timestamp 1621261055
transform 1 0 53760 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_556
timestamp 1621261055
transform 1 0 54528 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_564
timestamp 1621261055
transform 1 0 55296 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_793
timestamp 1621261055
transform 1 0 56640 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_572
timestamp 1621261055
transform 1 0 56064 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_576
timestamp 1621261055
transform 1 0 56448 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_579
timestamp 1621261055
transform 1 0 56736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_587
timestamp 1621261055
transform 1 0 57504 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_117
timestamp 1621261055
transform -1 0 58848 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_595
timestamp 1621261055
transform 1 0 58272 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_118
timestamp 1621261055
transform 1 0 1152 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_4
timestamp 1621261055
transform 1 0 1536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_12
timestamp 1621261055
transform 1 0 2304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_20
timestamp 1621261055
transform 1 0 3072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_28
timestamp 1621261055
transform 1 0 3840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_36
timestamp 1621261055
transform 1 0 4608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_794
timestamp 1621261055
transform 1 0 6432 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_44
timestamp 1621261055
transform 1 0 5376 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_52
timestamp 1621261055
transform 1 0 6144 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_54
timestamp 1621261055
transform 1 0 6336 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_56
timestamp 1621261055
transform 1 0 6528 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_64
timestamp 1621261055
transform 1 0 7296 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_72
timestamp 1621261055
transform 1 0 8064 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_80
timestamp 1621261055
transform 1 0 8832 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_88
timestamp 1621261055
transform 1 0 9600 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_96
timestamp 1621261055
transform 1 0 10368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_104
timestamp 1621261055
transform 1 0 11136 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_795
timestamp 1621261055
transform 1 0 11712 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_108
timestamp 1621261055
transform 1 0 11520 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_111
timestamp 1621261055
transform 1 0 11808 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_119
timestamp 1621261055
transform 1 0 12576 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_127
timestamp 1621261055
transform 1 0 13344 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_135
timestamp 1621261055
transform 1 0 14112 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_143
timestamp 1621261055
transform 1 0 14880 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _130_
timestamp 1621261055
transform 1 0 16320 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_796
timestamp 1621261055
transform 1 0 16992 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_197
timestamp 1621261055
transform 1 0 16128 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_59_151
timestamp 1621261055
transform 1 0 15648 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_59_155
timestamp 1621261055
transform 1 0 16032 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_161
timestamp 1621261055
transform 1 0 16608 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_166
timestamp 1621261055
transform 1 0 17088 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_174
timestamp 1621261055
transform 1 0 17856 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_182
timestamp 1621261055
transform 1 0 18624 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_190
timestamp 1621261055
transform 1 0 19392 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_198
timestamp 1621261055
transform 1 0 20160 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_206
timestamp 1621261055
transform 1 0 20928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_797
timestamp 1621261055
transform 1 0 22272 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_214
timestamp 1621261055
transform 1 0 21696 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_218
timestamp 1621261055
transform 1 0 22080 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_221
timestamp 1621261055
transform 1 0 22368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_229
timestamp 1621261055
transform 1 0 23136 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_237
timestamp 1621261055
transform 1 0 23904 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_245
timestamp 1621261055
transform 1 0 24672 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_253
timestamp 1621261055
transform 1 0 25440 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_261
timestamp 1621261055
transform 1 0 26208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_269
timestamp 1621261055
transform 1 0 26976 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_273
timestamp 1621261055
transform 1 0 27360 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_798
timestamp 1621261055
transform 1 0 27552 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_276
timestamp 1621261055
transform 1 0 27648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_284
timestamp 1621261055
transform 1 0 28416 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_292
timestamp 1621261055
transform 1 0 29184 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_300
timestamp 1621261055
transform 1 0 29952 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_308
timestamp 1621261055
transform 1 0 30720 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_799
timestamp 1621261055
transform 1 0 32832 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_316
timestamp 1621261055
transform 1 0 31488 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_324
timestamp 1621261055
transform 1 0 32256 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_328
timestamp 1621261055
transform 1 0 32640 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_331
timestamp 1621261055
transform 1 0 32928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_339
timestamp 1621261055
transform 1 0 33696 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_347
timestamp 1621261055
transform 1 0 34464 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_355
timestamp 1621261055
transform 1 0 35232 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_363
timestamp 1621261055
transform 1 0 36000 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_371
timestamp 1621261055
transform 1 0 36768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_800
timestamp 1621261055
transform 1 0 38112 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_379
timestamp 1621261055
transform 1 0 37536 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_383
timestamp 1621261055
transform 1 0 37920 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_386
timestamp 1621261055
transform 1 0 38208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_394
timestamp 1621261055
transform 1 0 38976 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_402
timestamp 1621261055
transform 1 0 39744 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_410
timestamp 1621261055
transform 1 0 40512 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_418
timestamp 1621261055
transform 1 0 41280 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_801
timestamp 1621261055
transform 1 0 43392 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_426
timestamp 1621261055
transform 1 0 42048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_434
timestamp 1621261055
transform 1 0 42816 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_438
timestamp 1621261055
transform 1 0 43200 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_441
timestamp 1621261055
transform 1 0 43488 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_449
timestamp 1621261055
transform 1 0 44256 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_457
timestamp 1621261055
transform 1 0 45024 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_465
timestamp 1621261055
transform 1 0 45792 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_473
timestamp 1621261055
transform 1 0 46560 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_481
timestamp 1621261055
transform 1 0 47328 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _040_
timestamp 1621261055
transform 1 0 48000 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_802
timestamp 1621261055
transform 1 0 48672 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_485
timestamp 1621261055
transform 1 0 47712 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_487
timestamp 1621261055
transform 1 0 47904 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_491
timestamp 1621261055
transform 1 0 48288 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_496
timestamp 1621261055
transform 1 0 48768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_504
timestamp 1621261055
transform 1 0 49536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_512
timestamp 1621261055
transform 1 0 50304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_520
timestamp 1621261055
transform 1 0 51072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_528
timestamp 1621261055
transform 1 0 51840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_536
timestamp 1621261055
transform 1 0 52608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_544
timestamp 1621261055
transform 1 0 53376 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_803
timestamp 1621261055
transform 1 0 53952 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_548
timestamp 1621261055
transform 1 0 53760 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_551
timestamp 1621261055
transform 1 0 54048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_559
timestamp 1621261055
transform 1 0 54816 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_567
timestamp 1621261055
transform 1 0 55584 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_575
timestamp 1621261055
transform 1 0 56352 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_583
timestamp 1621261055
transform 1 0 57120 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_119
timestamp 1621261055
transform -1 0 58848 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_59_591
timestamp 1621261055
transform 1 0 57888 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_595
timestamp 1621261055
transform 1 0 58272 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_120
timestamp 1621261055
transform 1 0 1152 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_60_4
timestamp 1621261055
transform 1 0 1536 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_12
timestamp 1621261055
transform 1 0 2304 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_20
timestamp 1621261055
transform 1 0 3072 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_804
timestamp 1621261055
transform 1 0 3840 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_29
timestamp 1621261055
transform 1 0 3936 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_37
timestamp 1621261055
transform 1 0 4704 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_45
timestamp 1621261055
transform 1 0 5472 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_53
timestamp 1621261055
transform 1 0 6240 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_61
timestamp 1621261055
transform 1 0 7008 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_805
timestamp 1621261055
transform 1 0 9120 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_69
timestamp 1621261055
transform 1 0 7776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_77
timestamp 1621261055
transform 1 0 8544 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_81
timestamp 1621261055
transform 1 0 8928 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_84
timestamp 1621261055
transform 1 0 9216 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _092_
timestamp 1621261055
transform 1 0 11040 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_162
timestamp 1621261055
transform 1 0 10848 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_92
timestamp 1621261055
transform 1 0 9984 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_60_100
timestamp 1621261055
transform 1 0 10752 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_106
timestamp 1621261055
transform 1 0 11328 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_114
timestamp 1621261055
transform 1 0 12096 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_122
timestamp 1621261055
transform 1 0 12864 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_806
timestamp 1621261055
transform 1 0 14400 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_130
timestamp 1621261055
transform 1 0 13632 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_139
timestamp 1621261055
transform 1 0 14496 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_147
timestamp 1621261055
transform 1 0 15264 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_155
timestamp 1621261055
transform 1 0 16032 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_163
timestamp 1621261055
transform 1 0 16800 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_171
timestamp 1621261055
transform 1 0 17568 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_179
timestamp 1621261055
transform 1 0 18336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_187
timestamp 1621261055
transform 1 0 19104 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_807
timestamp 1621261055
transform 1 0 19680 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_191
timestamp 1621261055
transform 1 0 19488 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_194
timestamp 1621261055
transform 1 0 19776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_202
timestamp 1621261055
transform 1 0 20544 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_210
timestamp 1621261055
transform 1 0 21312 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_218
timestamp 1621261055
transform 1 0 22080 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_226
timestamp 1621261055
transform 1 0 22848 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_808
timestamp 1621261055
transform 1 0 24960 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_234
timestamp 1621261055
transform 1 0 23616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_242
timestamp 1621261055
transform 1 0 24384 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_246
timestamp 1621261055
transform 1 0 24768 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_249
timestamp 1621261055
transform 1 0 25056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _094_
timestamp 1621261055
transform 1 0 26016 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_166
timestamp 1621261055
transform 1 0 25824 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_262
timestamp 1621261055
transform 1 0 26304 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_270
timestamp 1621261055
transform 1 0 27072 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_278
timestamp 1621261055
transform 1 0 27840 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_286
timestamp 1621261055
transform 1 0 28608 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_294
timestamp 1621261055
transform 1 0 29376 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_809
timestamp 1621261055
transform 1 0 30240 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_60_302
timestamp 1621261055
transform 1 0 30144 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_304
timestamp 1621261055
transform 1 0 30336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_312
timestamp 1621261055
transform 1 0 31104 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_320
timestamp 1621261055
transform 1 0 31872 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_328
timestamp 1621261055
transform 1 0 32640 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_336
timestamp 1621261055
transform 1 0 33408 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_344
timestamp 1621261055
transform 1 0 34176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_352
timestamp 1621261055
transform 1 0 34944 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_356
timestamp 1621261055
transform 1 0 35328 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_810
timestamp 1621261055
transform 1 0 35520 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_359
timestamp 1621261055
transform 1 0 35616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_367
timestamp 1621261055
transform 1 0 36384 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_375
timestamp 1621261055
transform 1 0 37152 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_383
timestamp 1621261055
transform 1 0 37920 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_391
timestamp 1621261055
transform 1 0 38688 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_399
timestamp 1621261055
transform 1 0 39456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_811
timestamp 1621261055
transform 1 0 40800 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_407
timestamp 1621261055
transform 1 0 40224 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_411
timestamp 1621261055
transform 1 0 40608 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_414
timestamp 1621261055
transform 1 0 40896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_422
timestamp 1621261055
transform 1 0 41664 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_430
timestamp 1621261055
transform 1 0 42432 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_438
timestamp 1621261055
transform 1 0 43200 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _212_
timestamp 1621261055
transform -1 0 45696 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_225
timestamp 1621261055
transform -1 0 45408 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_446
timestamp 1621261055
transform 1 0 43968 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_454
timestamp 1621261055
transform 1 0 44736 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_60_458
timestamp 1621261055
transform 1 0 45120 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_812
timestamp 1621261055
transform 1 0 46080 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_464
timestamp 1621261055
transform 1 0 45696 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_60_469
timestamp 1621261055
transform 1 0 46176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_477
timestamp 1621261055
transform 1 0 46944 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_485
timestamp 1621261055
transform 1 0 47712 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_493
timestamp 1621261055
transform 1 0 48480 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_501
timestamp 1621261055
transform 1 0 49248 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_813
timestamp 1621261055
transform 1 0 51360 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_509
timestamp 1621261055
transform 1 0 50016 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_517
timestamp 1621261055
transform 1 0 50784 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_521
timestamp 1621261055
transform 1 0 51168 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_524
timestamp 1621261055
transform 1 0 51456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_532
timestamp 1621261055
transform 1 0 52224 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_540
timestamp 1621261055
transform 1 0 52992 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_548
timestamp 1621261055
transform 1 0 53760 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_556
timestamp 1621261055
transform 1 0 54528 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_564
timestamp 1621261055
transform 1 0 55296 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_814
timestamp 1621261055
transform 1 0 56640 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_572
timestamp 1621261055
transform 1 0 56064 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_576
timestamp 1621261055
transform 1 0 56448 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_579
timestamp 1621261055
transform 1 0 56736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_587
timestamp 1621261055
transform 1 0 57504 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_121
timestamp 1621261055
transform -1 0 58848 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_595
timestamp 1621261055
transform 1 0 58272 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_122
timestamp 1621261055
transform 1 0 1152 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_124
timestamp 1621261055
transform 1 0 1152 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_4
timestamp 1621261055
transform 1 0 1536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_12
timestamp 1621261055
transform 1 0 2304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_20
timestamp 1621261055
transform 1 0 3072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_4
timestamp 1621261055
transform 1 0 1536 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_12
timestamp 1621261055
transform 1 0 2304 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_20
timestamp 1621261055
transform 1 0 3072 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_825
timestamp 1621261055
transform 1 0 3840 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_28
timestamp 1621261055
transform 1 0 3840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_36
timestamp 1621261055
transform 1 0 4608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_29
timestamp 1621261055
transform 1 0 3936 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_37
timestamp 1621261055
transform 1 0 4704 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_815
timestamp 1621261055
transform 1 0 6432 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_44
timestamp 1621261055
transform 1 0 5376 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_52
timestamp 1621261055
transform 1 0 6144 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_61_54
timestamp 1621261055
transform 1 0 6336 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_56
timestamp 1621261055
transform 1 0 6528 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_45
timestamp 1621261055
transform 1 0 5472 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_53
timestamp 1621261055
transform 1 0 6240 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_61
timestamp 1621261055
transform 1 0 7008 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_826
timestamp 1621261055
transform 1 0 9120 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_64
timestamp 1621261055
transform 1 0 7296 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_72
timestamp 1621261055
transform 1 0 8064 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_80
timestamp 1621261055
transform 1 0 8832 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_69
timestamp 1621261055
transform 1 0 7776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_77
timestamp 1621261055
transform 1 0 8544 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_81
timestamp 1621261055
transform 1 0 8928 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_84
timestamp 1621261055
transform 1 0 9216 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_88
timestamp 1621261055
transform 1 0 9600 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_96
timestamp 1621261055
transform 1 0 10368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_104
timestamp 1621261055
transform 1 0 11136 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_92
timestamp 1621261055
transform 1 0 9984 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_100
timestamp 1621261055
transform 1 0 10752 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_816
timestamp 1621261055
transform 1 0 11712 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_108
timestamp 1621261055
transform 1 0 11520 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_111
timestamp 1621261055
transform 1 0 11808 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_119
timestamp 1621261055
transform 1 0 12576 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_108
timestamp 1621261055
transform 1 0 11520 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_116
timestamp 1621261055
transform 1 0 12288 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_124
timestamp 1621261055
transform 1 0 13056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _218_
timestamp 1621261055
transform 1 0 13536 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_827
timestamp 1621261055
transform 1 0 14400 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_127
timestamp 1621261055
transform 1 0 13344 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_132
timestamp 1621261055
transform 1 0 13824 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_140
timestamp 1621261055
transform 1 0 14592 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_132
timestamp 1621261055
transform 1 0 13824 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_136
timestamp 1621261055
transform 1 0 14208 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_139
timestamp 1621261055
transform 1 0 14496 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_147
timestamp 1621261055
transform 1 0 15264 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_817
timestamp 1621261055
transform 1 0 16992 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_148
timestamp 1621261055
transform 1 0 15360 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_156
timestamp 1621261055
transform 1 0 16128 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_164
timestamp 1621261055
transform 1 0 16896 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_166
timestamp 1621261055
transform 1 0 17088 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_155
timestamp 1621261055
transform 1 0 16032 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_163
timestamp 1621261055
transform 1 0 16800 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_174
timestamp 1621261055
transform 1 0 17856 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_182
timestamp 1621261055
transform 1 0 18624 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_171
timestamp 1621261055
transform 1 0 17568 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_179
timestamp 1621261055
transform 1 0 18336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_187
timestamp 1621261055
transform 1 0 19104 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_828
timestamp 1621261055
transform 1 0 19680 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_190
timestamp 1621261055
transform 1 0 19392 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_198
timestamp 1621261055
transform 1 0 20160 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_206
timestamp 1621261055
transform 1 0 20928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_191
timestamp 1621261055
transform 1 0 19488 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_194
timestamp 1621261055
transform 1 0 19776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_202
timestamp 1621261055
transform 1 0 20544 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_210
timestamp 1621261055
transform 1 0 21312 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_818
timestamp 1621261055
transform 1 0 22272 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_214
timestamp 1621261055
transform 1 0 21696 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_218
timestamp 1621261055
transform 1 0 22080 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_221
timestamp 1621261055
transform 1 0 22368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_229
timestamp 1621261055
transform 1 0 23136 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_218
timestamp 1621261055
transform 1 0 22080 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_226
timestamp 1621261055
transform 1 0 22848 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_829
timestamp 1621261055
transform 1 0 24960 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_237
timestamp 1621261055
transform 1 0 23904 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_245
timestamp 1621261055
transform 1 0 24672 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_234
timestamp 1621261055
transform 1 0 23616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_242
timestamp 1621261055
transform 1 0 24384 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_246
timestamp 1621261055
transform 1 0 24768 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_249
timestamp 1621261055
transform 1 0 25056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_253
timestamp 1621261055
transform 1 0 25440 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_261
timestamp 1621261055
transform 1 0 26208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_269
timestamp 1621261055
transform 1 0 26976 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_273
timestamp 1621261055
transform 1 0 27360 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_257
timestamp 1621261055
transform 1 0 25824 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_265
timestamp 1621261055
transform 1 0 26592 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_273
timestamp 1621261055
transform 1 0 27360 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_819
timestamp 1621261055
transform 1 0 27552 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_276
timestamp 1621261055
transform 1 0 27648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_284
timestamp 1621261055
transform 1 0 28416 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_292
timestamp 1621261055
transform 1 0 29184 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_281
timestamp 1621261055
transform 1 0 28128 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_289
timestamp 1621261055
transform 1 0 28896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_830
timestamp 1621261055
transform 1 0 30240 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_300
timestamp 1621261055
transform 1 0 29952 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_308
timestamp 1621261055
transform 1 0 30720 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_297
timestamp 1621261055
transform 1 0 29664 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_301
timestamp 1621261055
transform 1 0 30048 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_304
timestamp 1621261055
transform 1 0 30336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_312
timestamp 1621261055
transform 1 0 31104 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_820
timestamp 1621261055
transform 1 0 32832 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_316
timestamp 1621261055
transform 1 0 31488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_324
timestamp 1621261055
transform 1 0 32256 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_328
timestamp 1621261055
transform 1 0 32640 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_331
timestamp 1621261055
transform 1 0 32928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_320
timestamp 1621261055
transform 1 0 31872 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_328
timestamp 1621261055
transform 1 0 32640 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_336
timestamp 1621261055
transform 1 0 33408 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_339
timestamp 1621261055
transform 1 0 33696 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_347
timestamp 1621261055
transform 1 0 34464 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_355
timestamp 1621261055
transform 1 0 35232 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_344
timestamp 1621261055
transform 1 0 34176 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_352
timestamp 1621261055
transform 1 0 34944 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_356
timestamp 1621261055
transform 1 0 35328 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _172_
timestamp 1621261055
transform 1 0 37152 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_831
timestamp 1621261055
transform 1 0 35520 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_112
timestamp 1621261055
transform 1 0 36960 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_363
timestamp 1621261055
transform 1 0 36000 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_371
timestamp 1621261055
transform 1 0 36768 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_61_378
timestamp 1621261055
transform 1 0 37440 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_359
timestamp 1621261055
transform 1 0 35616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_367
timestamp 1621261055
transform 1 0 36384 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_375
timestamp 1621261055
transform 1 0 37152 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_383
timestamp 1621261055
transform 1 0 37920 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_386
timestamp 1621261055
transform 1 0 38208 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_61_384
timestamp 1621261055
transform 1 0 38016 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_382
timestamp 1621261055
transform 1 0 37824 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_821
timestamp 1621261055
transform 1 0 38112 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_391
timestamp 1621261055
transform 1 0 38688 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_393
timestamp 1621261055
transform 1 0 38880 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_142
timestamp 1621261055
transform -1 0 38592 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _082_
timestamp 1621261055
transform -1 0 38880 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_399
timestamp 1621261055
transform 1 0 39456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_832
timestamp 1621261055
transform 1 0 40800 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_401
timestamp 1621261055
transform 1 0 39648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_409
timestamp 1621261055
transform 1 0 40416 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_417
timestamp 1621261055
transform 1 0 41184 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_407
timestamp 1621261055
transform 1 0 40224 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_411
timestamp 1621261055
transform 1 0 40608 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_414
timestamp 1621261055
transform 1 0 40896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_822
timestamp 1621261055
transform 1 0 43392 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_425
timestamp 1621261055
transform 1 0 41952 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_433
timestamp 1621261055
transform 1 0 42720 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_437
timestamp 1621261055
transform 1 0 43104 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_61_439
timestamp 1621261055
transform 1 0 43296 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_441
timestamp 1621261055
transform 1 0 43488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_422
timestamp 1621261055
transform 1 0 41664 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_430
timestamp 1621261055
transform 1 0 42432 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_438
timestamp 1621261055
transform 1 0 43200 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_449
timestamp 1621261055
transform 1 0 44256 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_457
timestamp 1621261055
transform 1 0 45024 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_446
timestamp 1621261055
transform 1 0 43968 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_454
timestamp 1621261055
transform 1 0 44736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_462
timestamp 1621261055
transform 1 0 45504 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_62_469
timestamp 1621261055
transform 1 0 46176 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_466
timestamp 1621261055
transform 1 0 45888 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_465
timestamp 1621261055
transform 1 0 45792 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_833
timestamp 1621261055
transform 1 0 46080 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_473
timestamp 1621261055
transform 1 0 46560 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_473
timestamp 1621261055
transform 1 0 46560 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_221
timestamp 1621261055
transform -1 0 46944 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _207_
timestamp 1621261055
transform -1 0 47232 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_62_480
timestamp 1621261055
transform 1 0 47232 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_481
timestamp 1621261055
transform 1 0 47328 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _089_
timestamp 1621261055
transform -1 0 48096 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_823
timestamp 1621261055
transform 1 0 48672 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_156
timestamp 1621261055
transform -1 0 47808 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_61_489
timestamp 1621261055
transform 1 0 48096 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_493
timestamp 1621261055
transform 1 0 48480 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_496
timestamp 1621261055
transform 1 0 48768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_504
timestamp 1621261055
transform 1 0 49536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_489
timestamp 1621261055
transform 1 0 48096 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_497
timestamp 1621261055
transform 1 0 48864 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_834
timestamp 1621261055
transform 1 0 51360 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_512
timestamp 1621261055
transform 1 0 50304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_520
timestamp 1621261055
transform 1 0 51072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_505
timestamp 1621261055
transform 1 0 49632 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_513
timestamp 1621261055
transform 1 0 50400 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_521
timestamp 1621261055
transform 1 0 51168 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_524
timestamp 1621261055
transform 1 0 51456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _146_
timestamp 1621261055
transform 1 0 51840 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_61_531
timestamp 1621261055
transform 1 0 52128 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_539
timestamp 1621261055
transform 1 0 52896 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_532
timestamp 1621261055
transform 1 0 52224 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_540
timestamp 1621261055
transform 1 0 52992 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_824
timestamp 1621261055
transform 1 0 53952 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_547
timestamp 1621261055
transform 1 0 53664 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_61_549
timestamp 1621261055
transform 1 0 53856 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_551
timestamp 1621261055
transform 1 0 54048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_559
timestamp 1621261055
transform 1 0 54816 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_567
timestamp 1621261055
transform 1 0 55584 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_548
timestamp 1621261055
transform 1 0 53760 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_556
timestamp 1621261055
transform 1 0 54528 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_564
timestamp 1621261055
transform 1 0 55296 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_835
timestamp 1621261055
transform 1 0 56640 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_575
timestamp 1621261055
transform 1 0 56352 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_583
timestamp 1621261055
transform 1 0 57120 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_572
timestamp 1621261055
transform 1 0 56064 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_576
timestamp 1621261055
transform 1 0 56448 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_579
timestamp 1621261055
transform 1 0 56736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_587
timestamp 1621261055
transform 1 0 57504 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_123
timestamp 1621261055
transform -1 0 58848 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_125
timestamp 1621261055
transform -1 0 58848 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_61_591
timestamp 1621261055
transform 1 0 57888 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_595
timestamp 1621261055
transform 1 0 58272 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_595
timestamp 1621261055
transform 1 0 58272 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_126
timestamp 1621261055
transform 1 0 1152 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_4
timestamp 1621261055
transform 1 0 1536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_12
timestamp 1621261055
transform 1 0 2304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_20
timestamp 1621261055
transform 1 0 3072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_28
timestamp 1621261055
transform 1 0 3840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_36
timestamp 1621261055
transform 1 0 4608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_836
timestamp 1621261055
transform 1 0 6432 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_44
timestamp 1621261055
transform 1 0 5376 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_52
timestamp 1621261055
transform 1 0 6144 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_54
timestamp 1621261055
transform 1 0 6336 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_56
timestamp 1621261055
transform 1 0 6528 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_64
timestamp 1621261055
transform 1 0 7296 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_72
timestamp 1621261055
transform 1 0 8064 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_80
timestamp 1621261055
transform 1 0 8832 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_88
timestamp 1621261055
transform 1 0 9600 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_96
timestamp 1621261055
transform 1 0 10368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_104
timestamp 1621261055
transform 1 0 11136 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_837
timestamp 1621261055
transform 1 0 11712 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_108
timestamp 1621261055
transform 1 0 11520 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_111
timestamp 1621261055
transform 1 0 11808 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_119
timestamp 1621261055
transform 1 0 12576 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_127
timestamp 1621261055
transform 1 0 13344 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_135
timestamp 1621261055
transform 1 0 14112 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_143
timestamp 1621261055
transform 1 0 14880 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_838
timestamp 1621261055
transform 1 0 16992 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_151
timestamp 1621261055
transform 1 0 15648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_159
timestamp 1621261055
transform 1 0 16416 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_163
timestamp 1621261055
transform 1 0 16800 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_166
timestamp 1621261055
transform 1 0 17088 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_174
timestamp 1621261055
transform 1 0 17856 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_182
timestamp 1621261055
transform 1 0 18624 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_190
timestamp 1621261055
transform 1 0 19392 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_198
timestamp 1621261055
transform 1 0 20160 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_206
timestamp 1621261055
transform 1 0 20928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_839
timestamp 1621261055
transform 1 0 22272 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_214
timestamp 1621261055
transform 1 0 21696 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_218
timestamp 1621261055
transform 1 0 22080 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_221
timestamp 1621261055
transform 1 0 22368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_229
timestamp 1621261055
transform 1 0 23136 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_237
timestamp 1621261055
transform 1 0 23904 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_245
timestamp 1621261055
transform 1 0 24672 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_253
timestamp 1621261055
transform 1 0 25440 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_261
timestamp 1621261055
transform 1 0 26208 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_269
timestamp 1621261055
transform 1 0 26976 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_273
timestamp 1621261055
transform 1 0 27360 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_840
timestamp 1621261055
transform 1 0 27552 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_276
timestamp 1621261055
transform 1 0 27648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_284
timestamp 1621261055
transform 1 0 28416 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_292
timestamp 1621261055
transform 1 0 29184 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_300
timestamp 1621261055
transform 1 0 29952 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_308
timestamp 1621261055
transform 1 0 30720 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_841
timestamp 1621261055
transform 1 0 32832 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_316
timestamp 1621261055
transform 1 0 31488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_324
timestamp 1621261055
transform 1 0 32256 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_328
timestamp 1621261055
transform 1 0 32640 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_331
timestamp 1621261055
transform 1 0 32928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_339
timestamp 1621261055
transform 1 0 33696 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_347
timestamp 1621261055
transform 1 0 34464 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_355
timestamp 1621261055
transform 1 0 35232 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_363
timestamp 1621261055
transform 1 0 36000 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_371
timestamp 1621261055
transform 1 0 36768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _214_
timestamp 1621261055
transform -1 0 39360 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_842
timestamp 1621261055
transform 1 0 38112 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_227
timestamp 1621261055
transform -1 0 39072 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_63_379
timestamp 1621261055
transform 1 0 37536 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_383
timestamp 1621261055
transform 1 0 37920 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_63_386
timestamp 1621261055
transform 1 0 38208 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_390
timestamp 1621261055
transform 1 0 38592 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_392
timestamp 1621261055
transform 1 0 38784 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_398
timestamp 1621261055
transform 1 0 39360 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_406
timestamp 1621261055
transform 1 0 40128 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_414
timestamp 1621261055
transform 1 0 40896 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_843
timestamp 1621261055
transform 1 0 43392 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_422
timestamp 1621261055
transform 1 0 41664 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_430
timestamp 1621261055
transform 1 0 42432 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_438
timestamp 1621261055
transform 1 0 43200 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_441
timestamp 1621261055
transform 1 0 43488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_449
timestamp 1621261055
transform 1 0 44256 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_457
timestamp 1621261055
transform 1 0 45024 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_465
timestamp 1621261055
transform 1 0 45792 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_473
timestamp 1621261055
transform 1 0 46560 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_481
timestamp 1621261055
transform 1 0 47328 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_844
timestamp 1621261055
transform 1 0 48672 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_489
timestamp 1621261055
transform 1 0 48096 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_493
timestamp 1621261055
transform 1 0 48480 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_496
timestamp 1621261055
transform 1 0 48768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_504
timestamp 1621261055
transform 1 0 49536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_512
timestamp 1621261055
transform 1 0 50304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_520
timestamp 1621261055
transform 1 0 51072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_528
timestamp 1621261055
transform 1 0 51840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_536
timestamp 1621261055
transform 1 0 52608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_544
timestamp 1621261055
transform 1 0 53376 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_845
timestamp 1621261055
transform 1 0 53952 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_548
timestamp 1621261055
transform 1 0 53760 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_551
timestamp 1621261055
transform 1 0 54048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_559
timestamp 1621261055
transform 1 0 54816 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_567
timestamp 1621261055
transform 1 0 55584 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_575
timestamp 1621261055
transform 1 0 56352 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_583
timestamp 1621261055
transform 1 0 57120 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_127
timestamp 1621261055
transform -1 0 58848 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_63_591
timestamp 1621261055
transform 1 0 57888 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_595
timestamp 1621261055
transform 1 0 58272 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_128
timestamp 1621261055
transform 1 0 1152 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_64_4
timestamp 1621261055
transform 1 0 1536 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_12
timestamp 1621261055
transform 1 0 2304 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_20
timestamp 1621261055
transform 1 0 3072 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_846
timestamp 1621261055
transform 1 0 3840 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_29
timestamp 1621261055
transform 1 0 3936 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_37
timestamp 1621261055
transform 1 0 4704 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_45
timestamp 1621261055
transform 1 0 5472 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_53
timestamp 1621261055
transform 1 0 6240 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_61
timestamp 1621261055
transform 1 0 7008 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_847
timestamp 1621261055
transform 1 0 9120 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_69
timestamp 1621261055
transform 1 0 7776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_77
timestamp 1621261055
transform 1 0 8544 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_81
timestamp 1621261055
transform 1 0 8928 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_84
timestamp 1621261055
transform 1 0 9216 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_92
timestamp 1621261055
transform 1 0 9984 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_100
timestamp 1621261055
transform 1 0 10752 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_108
timestamp 1621261055
transform 1 0 11520 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_116
timestamp 1621261055
transform 1 0 12288 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_124
timestamp 1621261055
transform 1 0 13056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_848
timestamp 1621261055
transform 1 0 14400 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_132
timestamp 1621261055
transform 1 0 13824 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_136
timestamp 1621261055
transform 1 0 14208 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_139
timestamp 1621261055
transform 1 0 14496 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_147
timestamp 1621261055
transform 1 0 15264 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_155
timestamp 1621261055
transform 1 0 16032 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_163
timestamp 1621261055
transform 1 0 16800 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_171
timestamp 1621261055
transform 1 0 17568 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_179
timestamp 1621261055
transform 1 0 18336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_187
timestamp 1621261055
transform 1 0 19104 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_849
timestamp 1621261055
transform 1 0 19680 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_191
timestamp 1621261055
transform 1 0 19488 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_194
timestamp 1621261055
transform 1 0 19776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_202
timestamp 1621261055
transform 1 0 20544 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_210
timestamp 1621261055
transform 1 0 21312 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_218
timestamp 1621261055
transform 1 0 22080 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_226
timestamp 1621261055
transform 1 0 22848 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_850
timestamp 1621261055
transform 1 0 24960 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_234
timestamp 1621261055
transform 1 0 23616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_242
timestamp 1621261055
transform 1 0 24384 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_246
timestamp 1621261055
transform 1 0 24768 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_249
timestamp 1621261055
transform 1 0 25056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_257
timestamp 1621261055
transform 1 0 25824 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_265
timestamp 1621261055
transform 1 0 26592 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_273
timestamp 1621261055
transform 1 0 27360 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_281
timestamp 1621261055
transform 1 0 28128 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_289
timestamp 1621261055
transform 1 0 28896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_851
timestamp 1621261055
transform 1 0 30240 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_297
timestamp 1621261055
transform 1 0 29664 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_301
timestamp 1621261055
transform 1 0 30048 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_304
timestamp 1621261055
transform 1 0 30336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_312
timestamp 1621261055
transform 1 0 31104 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_320
timestamp 1621261055
transform 1 0 31872 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_328
timestamp 1621261055
transform 1 0 32640 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_336
timestamp 1621261055
transform 1 0 33408 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_344
timestamp 1621261055
transform 1 0 34176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_352
timestamp 1621261055
transform 1 0 34944 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_356
timestamp 1621261055
transform 1 0 35328 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_852
timestamp 1621261055
transform 1 0 35520 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_359
timestamp 1621261055
transform 1 0 35616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_367
timestamp 1621261055
transform 1 0 36384 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_375
timestamp 1621261055
transform 1 0 37152 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_383
timestamp 1621261055
transform 1 0 37920 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_391
timestamp 1621261055
transform 1 0 38688 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_399
timestamp 1621261055
transform 1 0 39456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_853
timestamp 1621261055
transform 1 0 40800 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_407
timestamp 1621261055
transform 1 0 40224 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_411
timestamp 1621261055
transform 1 0 40608 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_414
timestamp 1621261055
transform 1 0 40896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_422
timestamp 1621261055
transform 1 0 41664 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_430
timestamp 1621261055
transform 1 0 42432 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_438
timestamp 1621261055
transform 1 0 43200 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_446
timestamp 1621261055
transform 1 0 43968 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_454
timestamp 1621261055
transform 1 0 44736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_462
timestamp 1621261055
transform 1 0 45504 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_854
timestamp 1621261055
transform 1 0 46080 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_466
timestamp 1621261055
transform 1 0 45888 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_469
timestamp 1621261055
transform 1 0 46176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_477
timestamp 1621261055
transform 1 0 46944 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_485
timestamp 1621261055
transform 1 0 47712 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_493
timestamp 1621261055
transform 1 0 48480 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_501
timestamp 1621261055
transform 1 0 49248 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_855
timestamp 1621261055
transform 1 0 51360 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_509
timestamp 1621261055
transform 1 0 50016 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_517
timestamp 1621261055
transform 1 0 50784 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_521
timestamp 1621261055
transform 1 0 51168 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_524
timestamp 1621261055
transform 1 0 51456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_532
timestamp 1621261055
transform 1 0 52224 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_540
timestamp 1621261055
transform 1 0 52992 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_548
timestamp 1621261055
transform 1 0 53760 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_556
timestamp 1621261055
transform 1 0 54528 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_564
timestamp 1621261055
transform 1 0 55296 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_856
timestamp 1621261055
transform 1 0 56640 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_572
timestamp 1621261055
transform 1 0 56064 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_576
timestamp 1621261055
transform 1 0 56448 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_579
timestamp 1621261055
transform 1 0 56736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_587
timestamp 1621261055
transform 1 0 57504 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_129
timestamp 1621261055
transform -1 0 58848 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_595
timestamp 1621261055
transform 1 0 58272 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_130
timestamp 1621261055
transform 1 0 1152 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_4
timestamp 1621261055
transform 1 0 1536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_12
timestamp 1621261055
transform 1 0 2304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_20
timestamp 1621261055
transform 1 0 3072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_28
timestamp 1621261055
transform 1 0 3840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_36
timestamp 1621261055
transform 1 0 4608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_857
timestamp 1621261055
transform 1 0 6432 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_44
timestamp 1621261055
transform 1 0 5376 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_52
timestamp 1621261055
transform 1 0 6144 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_54
timestamp 1621261055
transform 1 0 6336 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_56
timestamp 1621261055
transform 1 0 6528 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_64
timestamp 1621261055
transform 1 0 7296 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_72
timestamp 1621261055
transform 1 0 8064 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_80
timestamp 1621261055
transform 1 0 8832 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_88
timestamp 1621261055
transform 1 0 9600 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_96
timestamp 1621261055
transform 1 0 10368 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_104
timestamp 1621261055
transform 1 0 11136 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_858
timestamp 1621261055
transform 1 0 11712 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_108
timestamp 1621261055
transform 1 0 11520 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_111
timestamp 1621261055
transform 1 0 11808 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_119
timestamp 1621261055
transform 1 0 12576 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_127
timestamp 1621261055
transform 1 0 13344 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_135
timestamp 1621261055
transform 1 0 14112 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_143
timestamp 1621261055
transform 1 0 14880 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_859
timestamp 1621261055
transform 1 0 16992 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_151
timestamp 1621261055
transform 1 0 15648 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_159
timestamp 1621261055
transform 1 0 16416 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_163
timestamp 1621261055
transform 1 0 16800 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_166
timestamp 1621261055
transform 1 0 17088 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_174
timestamp 1621261055
transform 1 0 17856 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_182
timestamp 1621261055
transform 1 0 18624 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_190
timestamp 1621261055
transform 1 0 19392 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_198
timestamp 1621261055
transform 1 0 20160 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_206
timestamp 1621261055
transform 1 0 20928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_860
timestamp 1621261055
transform 1 0 22272 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_214
timestamp 1621261055
transform 1 0 21696 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_218
timestamp 1621261055
transform 1 0 22080 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_221
timestamp 1621261055
transform 1 0 22368 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_229
timestamp 1621261055
transform 1 0 23136 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_237
timestamp 1621261055
transform 1 0 23904 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_245
timestamp 1621261055
transform 1 0 24672 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_253
timestamp 1621261055
transform 1 0 25440 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_261
timestamp 1621261055
transform 1 0 26208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_269
timestamp 1621261055
transform 1 0 26976 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_273
timestamp 1621261055
transform 1 0 27360 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _185_
timestamp 1621261055
transform 1 0 28032 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_861
timestamp 1621261055
transform 1 0 27552 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_127
timestamp 1621261055
transform 1 0 27840 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_276
timestamp 1621261055
transform 1 0 27648 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_283
timestamp 1621261055
transform 1 0 28320 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_291
timestamp 1621261055
transform 1 0 29088 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_299
timestamp 1621261055
transform 1 0 29856 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_307
timestamp 1621261055
transform 1 0 30624 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_315
timestamp 1621261055
transform 1 0 31392 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_862
timestamp 1621261055
transform 1 0 32832 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_323
timestamp 1621261055
transform 1 0 32160 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_327
timestamp 1621261055
transform 1 0 32544 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_329
timestamp 1621261055
transform 1 0 32736 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_331
timestamp 1621261055
transform 1 0 32928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_339
timestamp 1621261055
transform 1 0 33696 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_347
timestamp 1621261055
transform 1 0 34464 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_355
timestamp 1621261055
transform 1 0 35232 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_363
timestamp 1621261055
transform 1 0 36000 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_371
timestamp 1621261055
transform 1 0 36768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_863
timestamp 1621261055
transform 1 0 38112 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_379
timestamp 1621261055
transform 1 0 37536 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_383
timestamp 1621261055
transform 1 0 37920 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_386
timestamp 1621261055
transform 1 0 38208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_394
timestamp 1621261055
transform 1 0 38976 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _015_
timestamp 1621261055
transform 1 0 40224 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_65_402
timestamp 1621261055
transform 1 0 39744 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_65_406
timestamp 1621261055
transform 1 0 40128 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_410
timestamp 1621261055
transform 1 0 40512 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_418
timestamp 1621261055
transform 1 0 41280 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_864
timestamp 1621261055
transform 1 0 43392 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_426
timestamp 1621261055
transform 1 0 42048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_434
timestamp 1621261055
transform 1 0 42816 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_438
timestamp 1621261055
transform 1 0 43200 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_441
timestamp 1621261055
transform 1 0 43488 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_449
timestamp 1621261055
transform 1 0 44256 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_457
timestamp 1621261055
transform 1 0 45024 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_465
timestamp 1621261055
transform 1 0 45792 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_473
timestamp 1621261055
transform 1 0 46560 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_481
timestamp 1621261055
transform 1 0 47328 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_865
timestamp 1621261055
transform 1 0 48672 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_489
timestamp 1621261055
transform 1 0 48096 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_493
timestamp 1621261055
transform 1 0 48480 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_496
timestamp 1621261055
transform 1 0 48768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_504
timestamp 1621261055
transform 1 0 49536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_512
timestamp 1621261055
transform 1 0 50304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_520
timestamp 1621261055
transform 1 0 51072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_528
timestamp 1621261055
transform 1 0 51840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_536
timestamp 1621261055
transform 1 0 52608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_544
timestamp 1621261055
transform 1 0 53376 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_866
timestamp 1621261055
transform 1 0 53952 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_548
timestamp 1621261055
transform 1 0 53760 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_551
timestamp 1621261055
transform 1 0 54048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_559
timestamp 1621261055
transform 1 0 54816 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_567
timestamp 1621261055
transform 1 0 55584 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_575
timestamp 1621261055
transform 1 0 56352 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_583
timestamp 1621261055
transform 1 0 57120 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_131
timestamp 1621261055
transform -1 0 58848 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_65_591
timestamp 1621261055
transform 1 0 57888 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_595
timestamp 1621261055
transform 1 0 58272 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_132
timestamp 1621261055
transform 1 0 1152 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_66_4
timestamp 1621261055
transform 1 0 1536 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_12
timestamp 1621261055
transform 1 0 2304 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_20
timestamp 1621261055
transform 1 0 3072 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _179_
timestamp 1621261055
transform 1 0 4608 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_867
timestamp 1621261055
transform 1 0 3840 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_122
timestamp 1621261055
transform 1 0 4416 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_66_29
timestamp 1621261055
transform 1 0 3936 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_66_33
timestamp 1621261055
transform 1 0 4320 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_39
timestamp 1621261055
transform 1 0 4896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_47
timestamp 1621261055
transform 1 0 5664 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_55
timestamp 1621261055
transform 1 0 6432 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_63
timestamp 1621261055
transform 1 0 7200 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_868
timestamp 1621261055
transform 1 0 9120 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_71
timestamp 1621261055
transform 1 0 7968 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_79
timestamp 1621261055
transform 1 0 8736 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_66_84
timestamp 1621261055
transform 1 0 9216 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_92
timestamp 1621261055
transform 1 0 9984 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_100
timestamp 1621261055
transform 1 0 10752 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_108
timestamp 1621261055
transform 1 0 11520 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_116
timestamp 1621261055
transform 1 0 12288 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_124
timestamp 1621261055
transform 1 0 13056 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _083_
timestamp 1621261055
transform 1 0 13728 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_869
timestamp 1621261055
transform 1 0 14400 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_138
timestamp 1621261055
transform 1 0 15264 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_144
timestamp 1621261055
transform 1 0 13536 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_66_128
timestamp 1621261055
transform 1 0 13440 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_134
timestamp 1621261055
transform 1 0 14016 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_66_139
timestamp 1621261055
transform 1 0 14496 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _076_
timestamp 1621261055
transform 1 0 15456 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_66_152
timestamp 1621261055
transform 1 0 15744 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_160
timestamp 1621261055
transform 1 0 16512 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_168
timestamp 1621261055
transform 1 0 17280 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_176
timestamp 1621261055
transform 1 0 18048 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_184
timestamp 1621261055
transform 1 0 18816 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_870
timestamp 1621261055
transform 1 0 19680 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_66_192
timestamp 1621261055
transform 1 0 19584 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_194
timestamp 1621261055
transform 1 0 19776 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_202
timestamp 1621261055
transform 1 0 20544 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_210
timestamp 1621261055
transform 1 0 21312 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_218
timestamp 1621261055
transform 1 0 22080 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_226
timestamp 1621261055
transform 1 0 22848 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_871
timestamp 1621261055
transform 1 0 24960 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_234
timestamp 1621261055
transform 1 0 23616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_242
timestamp 1621261055
transform 1 0 24384 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_246
timestamp 1621261055
transform 1 0 24768 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_249
timestamp 1621261055
transform 1 0 25056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_257
timestamp 1621261055
transform 1 0 25824 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_265
timestamp 1621261055
transform 1 0 26592 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_273
timestamp 1621261055
transform 1 0 27360 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_281
timestamp 1621261055
transform 1 0 28128 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_289
timestamp 1621261055
transform 1 0 28896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_872
timestamp 1621261055
transform 1 0 30240 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_297
timestamp 1621261055
transform 1 0 29664 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_301
timestamp 1621261055
transform 1 0 30048 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_304
timestamp 1621261055
transform 1 0 30336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_312
timestamp 1621261055
transform 1 0 31104 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _010_
timestamp 1621261055
transform 1 0 31680 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_316
timestamp 1621261055
transform 1 0 31488 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_321
timestamp 1621261055
transform 1 0 31968 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_329
timestamp 1621261055
transform 1 0 32736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_337
timestamp 1621261055
transform 1 0 33504 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_345
timestamp 1621261055
transform 1 0 34272 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_353
timestamp 1621261055
transform 1 0 35040 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_66_357
timestamp 1621261055
transform 1 0 35424 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_873
timestamp 1621261055
transform 1 0 35520 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_359
timestamp 1621261055
transform 1 0 35616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_367
timestamp 1621261055
transform 1 0 36384 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_375
timestamp 1621261055
transform 1 0 37152 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_383
timestamp 1621261055
transform 1 0 37920 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_391
timestamp 1621261055
transform 1 0 38688 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_399
timestamp 1621261055
transform 1 0 39456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_874
timestamp 1621261055
transform 1 0 40800 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_407
timestamp 1621261055
transform 1 0 40224 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_411
timestamp 1621261055
transform 1 0 40608 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_414
timestamp 1621261055
transform 1 0 40896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_422
timestamp 1621261055
transform 1 0 41664 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_430
timestamp 1621261055
transform 1 0 42432 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_438
timestamp 1621261055
transform 1 0 43200 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _065_
timestamp 1621261055
transform -1 0 45696 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_201
timestamp 1621261055
transform -1 0 45408 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_446
timestamp 1621261055
transform 1 0 43968 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_454
timestamp 1621261055
transform 1 0 44736 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_66_458
timestamp 1621261055
transform 1 0 45120 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_875
timestamp 1621261055
transform 1 0 46080 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_464
timestamp 1621261055
transform 1 0 45696 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_66_469
timestamp 1621261055
transform 1 0 46176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_477
timestamp 1621261055
transform 1 0 46944 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_485
timestamp 1621261055
transform 1 0 47712 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_493
timestamp 1621261055
transform 1 0 48480 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_501
timestamp 1621261055
transform 1 0 49248 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_876
timestamp 1621261055
transform 1 0 51360 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_509
timestamp 1621261055
transform 1 0 50016 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_517
timestamp 1621261055
transform 1 0 50784 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_521
timestamp 1621261055
transform 1 0 51168 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_524
timestamp 1621261055
transform 1 0 51456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_532
timestamp 1621261055
transform 1 0 52224 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_540
timestamp 1621261055
transform 1 0 52992 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_548
timestamp 1621261055
transform 1 0 53760 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_556
timestamp 1621261055
transform 1 0 54528 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_564
timestamp 1621261055
transform 1 0 55296 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_877
timestamp 1621261055
transform 1 0 56640 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_572
timestamp 1621261055
transform 1 0 56064 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_576
timestamp 1621261055
transform 1 0 56448 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_579
timestamp 1621261055
transform 1 0 56736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_587
timestamp 1621261055
transform 1 0 57504 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_133
timestamp 1621261055
transform -1 0 58848 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_595
timestamp 1621261055
transform 1 0 58272 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_134
timestamp 1621261055
transform 1 0 1152 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_67_4
timestamp 1621261055
transform 1 0 1536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_12
timestamp 1621261055
transform 1 0 2304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_20
timestamp 1621261055
transform 1 0 3072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_28
timestamp 1621261055
transform 1 0 3840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_36
timestamp 1621261055
transform 1 0 4608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_878
timestamp 1621261055
transform 1 0 6432 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_44
timestamp 1621261055
transform 1 0 5376 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_52
timestamp 1621261055
transform 1 0 6144 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_54
timestamp 1621261055
transform 1 0 6336 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_56
timestamp 1621261055
transform 1 0 6528 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_64
timestamp 1621261055
transform 1 0 7296 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_72
timestamp 1621261055
transform 1 0 8064 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_80
timestamp 1621261055
transform 1 0 8832 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_88
timestamp 1621261055
transform 1 0 9600 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_96
timestamp 1621261055
transform 1 0 10368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_104
timestamp 1621261055
transform 1 0 11136 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_879
timestamp 1621261055
transform 1 0 11712 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_108
timestamp 1621261055
transform 1 0 11520 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_111
timestamp 1621261055
transform 1 0 11808 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_119
timestamp 1621261055
transform 1 0 12576 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_127
timestamp 1621261055
transform 1 0 13344 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_135
timestamp 1621261055
transform 1 0 14112 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_143
timestamp 1621261055
transform 1 0 14880 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_880
timestamp 1621261055
transform 1 0 16992 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_192
timestamp 1621261055
transform 1 0 17280 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_151
timestamp 1621261055
transform 1 0 15648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_159
timestamp 1621261055
transform 1 0 16416 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_163
timestamp 1621261055
transform 1 0 16800 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_166
timestamp 1621261055
transform 1 0 17088 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _127_
timestamp 1621261055
transform 1 0 17472 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_67_173
timestamp 1621261055
transform 1 0 17760 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_181
timestamp 1621261055
transform 1 0 18528 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_189
timestamp 1621261055
transform 1 0 19296 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_197
timestamp 1621261055
transform 1 0 20064 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_205
timestamp 1621261055
transform 1 0 20832 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _031_
timestamp 1621261055
transform 1 0 23328 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_881
timestamp 1621261055
transform 1 0 22272 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_213
timestamp 1621261055
transform 1 0 21600 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_217
timestamp 1621261055
transform 1 0 21984 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_219
timestamp 1621261055
transform 1 0 22176 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_221
timestamp 1621261055
transform 1 0 22368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_229
timestamp 1621261055
transform 1 0 23136 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_234
timestamp 1621261055
transform 1 0 23616 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_242
timestamp 1621261055
transform 1 0 24384 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_250
timestamp 1621261055
transform 1 0 25152 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_258
timestamp 1621261055
transform 1 0 25920 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_266
timestamp 1621261055
transform 1 0 26688 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_882
timestamp 1621261055
transform 1 0 27552 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_67_274
timestamp 1621261055
transform 1 0 27456 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_276
timestamp 1621261055
transform 1 0 27648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_284
timestamp 1621261055
transform 1 0 28416 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_292
timestamp 1621261055
transform 1 0 29184 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_300
timestamp 1621261055
transform 1 0 29952 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_308
timestamp 1621261055
transform 1 0 30720 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_883
timestamp 1621261055
transform 1 0 32832 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_316
timestamp 1621261055
transform 1 0 31488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_324
timestamp 1621261055
transform 1 0 32256 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_328
timestamp 1621261055
transform 1 0 32640 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_331
timestamp 1621261055
transform 1 0 32928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_339
timestamp 1621261055
transform 1 0 33696 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_347
timestamp 1621261055
transform 1 0 34464 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_355
timestamp 1621261055
transform 1 0 35232 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_363
timestamp 1621261055
transform 1 0 36000 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_371
timestamp 1621261055
transform 1 0 36768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_884
timestamp 1621261055
transform 1 0 38112 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_379
timestamp 1621261055
transform 1 0 37536 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_383
timestamp 1621261055
transform 1 0 37920 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_386
timestamp 1621261055
transform 1 0 38208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_394
timestamp 1621261055
transform 1 0 38976 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_402
timestamp 1621261055
transform 1 0 39744 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_410
timestamp 1621261055
transform 1 0 40512 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_418
timestamp 1621261055
transform 1 0 41280 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_885
timestamp 1621261055
transform 1 0 43392 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_426
timestamp 1621261055
transform 1 0 42048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_434
timestamp 1621261055
transform 1 0 42816 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_438
timestamp 1621261055
transform 1 0 43200 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_441
timestamp 1621261055
transform 1 0 43488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_449
timestamp 1621261055
transform 1 0 44256 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_457
timestamp 1621261055
transform 1 0 45024 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_465
timestamp 1621261055
transform 1 0 45792 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_473
timestamp 1621261055
transform 1 0 46560 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_481
timestamp 1621261055
transform 1 0 47328 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_886
timestamp 1621261055
transform 1 0 48672 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_489
timestamp 1621261055
transform 1 0 48096 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_493
timestamp 1621261055
transform 1 0 48480 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_496
timestamp 1621261055
transform 1 0 48768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_504
timestamp 1621261055
transform 1 0 49536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_512
timestamp 1621261055
transform 1 0 50304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_520
timestamp 1621261055
transform 1 0 51072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_528
timestamp 1621261055
transform 1 0 51840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_536
timestamp 1621261055
transform 1 0 52608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_544
timestamp 1621261055
transform 1 0 53376 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_887
timestamp 1621261055
transform 1 0 53952 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_548
timestamp 1621261055
transform 1 0 53760 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_551
timestamp 1621261055
transform 1 0 54048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_559
timestamp 1621261055
transform 1 0 54816 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_567
timestamp 1621261055
transform 1 0 55584 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_575
timestamp 1621261055
transform 1 0 56352 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_583
timestamp 1621261055
transform 1 0 57120 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_135
timestamp 1621261055
transform -1 0 58848 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_67_591
timestamp 1621261055
transform 1 0 57888 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_595
timestamp 1621261055
transform 1 0 58272 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_136
timestamp 1621261055
transform 1 0 1152 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_4
timestamp 1621261055
transform 1 0 1536 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_12
timestamp 1621261055
transform 1 0 2304 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_20
timestamp 1621261055
transform 1 0 3072 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _197_
timestamp 1621261055
transform 1 0 4320 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_888
timestamp 1621261055
transform 1 0 3840 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_213
timestamp 1621261055
transform 1 0 4128 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_29
timestamp 1621261055
transform 1 0 3936 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_36
timestamp 1621261055
transform 1 0 4608 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_44
timestamp 1621261055
transform 1 0 5376 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_52
timestamp 1621261055
transform 1 0 6144 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_60
timestamp 1621261055
transform 1 0 6912 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_889
timestamp 1621261055
transform 1 0 9120 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_68
timestamp 1621261055
transform 1 0 7680 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_76
timestamp 1621261055
transform 1 0 8448 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_80
timestamp 1621261055
transform 1 0 8832 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_68_82
timestamp 1621261055
transform 1 0 9024 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_84
timestamp 1621261055
transform 1 0 9216 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_92
timestamp 1621261055
transform 1 0 9984 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_100
timestamp 1621261055
transform 1 0 10752 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_108
timestamp 1621261055
transform 1 0 11520 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_116
timestamp 1621261055
transform 1 0 12288 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_124
timestamp 1621261055
transform 1 0 13056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_890
timestamp 1621261055
transform 1 0 14400 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_132
timestamp 1621261055
transform 1 0 13824 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_136
timestamp 1621261055
transform 1 0 14208 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_139
timestamp 1621261055
transform 1 0 14496 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_147
timestamp 1621261055
transform 1 0 15264 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_155
timestamp 1621261055
transform 1 0 16032 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_163
timestamp 1621261055
transform 1 0 16800 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_171
timestamp 1621261055
transform 1 0 17568 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_179
timestamp 1621261055
transform 1 0 18336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_187
timestamp 1621261055
transform 1 0 19104 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_891
timestamp 1621261055
transform 1 0 19680 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_191
timestamp 1621261055
transform 1 0 19488 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_194
timestamp 1621261055
transform 1 0 19776 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_202
timestamp 1621261055
transform 1 0 20544 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_210
timestamp 1621261055
transform 1 0 21312 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_218
timestamp 1621261055
transform 1 0 22080 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_226
timestamp 1621261055
transform 1 0 22848 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_892
timestamp 1621261055
transform 1 0 24960 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_234
timestamp 1621261055
transform 1 0 23616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_242
timestamp 1621261055
transform 1 0 24384 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_246
timestamp 1621261055
transform 1 0 24768 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_249
timestamp 1621261055
transform 1 0 25056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_257
timestamp 1621261055
transform 1 0 25824 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_265
timestamp 1621261055
transform 1 0 26592 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_273
timestamp 1621261055
transform 1 0 27360 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_281
timestamp 1621261055
transform 1 0 28128 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_289
timestamp 1621261055
transform 1 0 28896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_893
timestamp 1621261055
transform 1 0 30240 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_297
timestamp 1621261055
transform 1 0 29664 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_301
timestamp 1621261055
transform 1 0 30048 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_304
timestamp 1621261055
transform 1 0 30336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_312
timestamp 1621261055
transform 1 0 31104 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_320
timestamp 1621261055
transform 1 0 31872 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_328
timestamp 1621261055
transform 1 0 32640 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_336
timestamp 1621261055
transform 1 0 33408 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_344
timestamp 1621261055
transform 1 0 34176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_352
timestamp 1621261055
transform 1 0 34944 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_356
timestamp 1621261055
transform 1 0 35328 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_894
timestamp 1621261055
transform 1 0 35520 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_359
timestamp 1621261055
transform 1 0 35616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_367
timestamp 1621261055
transform 1 0 36384 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_375
timestamp 1621261055
transform 1 0 37152 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_383
timestamp 1621261055
transform 1 0 37920 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_391
timestamp 1621261055
transform 1 0 38688 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_399
timestamp 1621261055
transform 1 0 39456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_895
timestamp 1621261055
transform 1 0 40800 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_407
timestamp 1621261055
transform 1 0 40224 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_411
timestamp 1621261055
transform 1 0 40608 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_414
timestamp 1621261055
transform 1 0 40896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_422
timestamp 1621261055
transform 1 0 41664 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_430
timestamp 1621261055
transform 1 0 42432 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_438
timestamp 1621261055
transform 1 0 43200 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_446
timestamp 1621261055
transform 1 0 43968 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_454
timestamp 1621261055
transform 1 0 44736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_462
timestamp 1621261055
transform 1 0 45504 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_896
timestamp 1621261055
transform 1 0 46080 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_466
timestamp 1621261055
transform 1 0 45888 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_469
timestamp 1621261055
transform 1 0 46176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_477
timestamp 1621261055
transform 1 0 46944 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_485
timestamp 1621261055
transform 1 0 47712 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_493
timestamp 1621261055
transform 1 0 48480 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_501
timestamp 1621261055
transform 1 0 49248 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_897
timestamp 1621261055
transform 1 0 51360 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_509
timestamp 1621261055
transform 1 0 50016 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_517
timestamp 1621261055
transform 1 0 50784 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_521
timestamp 1621261055
transform 1 0 51168 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_524
timestamp 1621261055
transform 1 0 51456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_532
timestamp 1621261055
transform 1 0 52224 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_540
timestamp 1621261055
transform 1 0 52992 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_548
timestamp 1621261055
transform 1 0 53760 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_556
timestamp 1621261055
transform 1 0 54528 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_564
timestamp 1621261055
transform 1 0 55296 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_898
timestamp 1621261055
transform 1 0 56640 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_572
timestamp 1621261055
transform 1 0 56064 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_576
timestamp 1621261055
transform 1 0 56448 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_579
timestamp 1621261055
transform 1 0 56736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_587
timestamp 1621261055
transform 1 0 57504 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _153_
timestamp 1621261055
transform 1 0 57792 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_137
timestamp 1621261055
transform -1 0 58848 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_68_589
timestamp 1621261055
transform 1 0 57696 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_593
timestamp 1621261055
transform 1 0 58080 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _084_
timestamp 1621261055
transform 1 0 1536 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_138
timestamp 1621261055
transform 1 0 1152 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_140
timestamp 1621261055
transform 1 0 1152 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_146
timestamp 1621261055
transform 1 0 1824 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_9
timestamp 1621261055
transform 1 0 2016 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_17
timestamp 1621261055
transform 1 0 2784 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_4
timestamp 1621261055
transform 1 0 1536 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_12
timestamp 1621261055
transform 1 0 2304 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_20
timestamp 1621261055
transform 1 0 3072 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_909
timestamp 1621261055
transform 1 0 3840 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_25
timestamp 1621261055
transform 1 0 3552 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_33
timestamp 1621261055
transform 1 0 4320 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_41
timestamp 1621261055
transform 1 0 5088 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_29
timestamp 1621261055
transform 1 0 3936 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_37
timestamp 1621261055
transform 1 0 4704 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _004_
timestamp 1621261055
transform 1 0 6240 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _206_
timestamp 1621261055
transform 1 0 7008 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_899
timestamp 1621261055
transform 1 0 6432 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_49
timestamp 1621261055
transform 1 0 5856 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_53
timestamp 1621261055
transform 1 0 6240 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_56
timestamp 1621261055
transform 1 0 6528 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_69_60
timestamp 1621261055
transform 1 0 6912 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_45
timestamp 1621261055
transform 1 0 5472 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_56
timestamp 1621261055
transform 1 0 6528 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_910
timestamp 1621261055
transform 1 0 9120 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_64
timestamp 1621261055
transform 1 0 7296 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_72
timestamp 1621261055
transform 1 0 8064 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_80
timestamp 1621261055
transform 1 0 8832 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_64
timestamp 1621261055
transform 1 0 7296 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_72
timestamp 1621261055
transform 1 0 8064 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_80
timestamp 1621261055
transform 1 0 8832 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_70_82
timestamp 1621261055
transform 1 0 9024 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_84
timestamp 1621261055
transform 1 0 9216 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_88
timestamp 1621261055
transform 1 0 9600 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_96
timestamp 1621261055
transform 1 0 10368 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_104
timestamp 1621261055
transform 1 0 11136 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_92
timestamp 1621261055
transform 1 0 9984 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_100
timestamp 1621261055
transform 1 0 10752 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_900
timestamp 1621261055
transform 1 0 11712 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_108
timestamp 1621261055
transform 1 0 11520 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_111
timestamp 1621261055
transform 1 0 11808 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_119
timestamp 1621261055
transform 1 0 12576 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_108
timestamp 1621261055
transform 1 0 11520 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_116
timestamp 1621261055
transform 1 0 12288 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_124
timestamp 1621261055
transform 1 0 13056 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_911
timestamp 1621261055
transform 1 0 14400 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_127
timestamp 1621261055
transform 1 0 13344 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_135
timestamp 1621261055
transform 1 0 14112 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_143
timestamp 1621261055
transform 1 0 14880 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_132
timestamp 1621261055
transform 1 0 13824 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_136
timestamp 1621261055
transform 1 0 14208 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_139
timestamp 1621261055
transform 1 0 14496 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_147
timestamp 1621261055
transform 1 0 15264 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_901
timestamp 1621261055
transform 1 0 16992 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_151
timestamp 1621261055
transform 1 0 15648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_159
timestamp 1621261055
transform 1 0 16416 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_163
timestamp 1621261055
transform 1 0 16800 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_166
timestamp 1621261055
transform 1 0 17088 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_155
timestamp 1621261055
transform 1 0 16032 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_163
timestamp 1621261055
transform 1 0 16800 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_174
timestamp 1621261055
transform 1 0 17856 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_182
timestamp 1621261055
transform 1 0 18624 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_171
timestamp 1621261055
transform 1 0 17568 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_179
timestamp 1621261055
transform 1 0 18336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_187
timestamp 1621261055
transform 1 0 19104 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_912
timestamp 1621261055
transform 1 0 19680 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_190
timestamp 1621261055
transform 1 0 19392 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_198
timestamp 1621261055
transform 1 0 20160 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_206
timestamp 1621261055
transform 1 0 20928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_191
timestamp 1621261055
transform 1 0 19488 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_194
timestamp 1621261055
transform 1 0 19776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_202
timestamp 1621261055
transform 1 0 20544 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_210
timestamp 1621261055
transform 1 0 21312 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_902
timestamp 1621261055
transform 1 0 22272 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_214
timestamp 1621261055
transform 1 0 21696 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_218
timestamp 1621261055
transform 1 0 22080 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_221
timestamp 1621261055
transform 1 0 22368 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_229
timestamp 1621261055
transform 1 0 23136 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_218
timestamp 1621261055
transform 1 0 22080 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_226
timestamp 1621261055
transform 1 0 22848 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_913
timestamp 1621261055
transform 1 0 24960 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_237
timestamp 1621261055
transform 1 0 23904 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_245
timestamp 1621261055
transform 1 0 24672 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_234
timestamp 1621261055
transform 1 0 23616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_242
timestamp 1621261055
transform 1 0 24384 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_246
timestamp 1621261055
transform 1 0 24768 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_249
timestamp 1621261055
transform 1 0 25056 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_253
timestamp 1621261055
transform 1 0 25440 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_261
timestamp 1621261055
transform 1 0 26208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_269
timestamp 1621261055
transform 1 0 26976 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_273
timestamp 1621261055
transform 1 0 27360 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_257
timestamp 1621261055
transform 1 0 25824 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_265
timestamp 1621261055
transform 1 0 26592 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_273
timestamp 1621261055
transform 1 0 27360 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _009_
timestamp 1621261055
transform 1 0 28512 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_903
timestamp 1621261055
transform 1 0 27552 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_276
timestamp 1621261055
transform 1 0 27648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_284
timestamp 1621261055
transform 1 0 28416 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_288
timestamp 1621261055
transform 1 0 28800 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_281
timestamp 1621261055
transform 1 0 28128 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_289
timestamp 1621261055
transform 1 0 28896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_914
timestamp 1621261055
transform 1 0 30240 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_296
timestamp 1621261055
transform 1 0 29568 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_304
timestamp 1621261055
transform 1 0 30336 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_312
timestamp 1621261055
transform 1 0 31104 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_297
timestamp 1621261055
transform 1 0 29664 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_301
timestamp 1621261055
transform 1 0 30048 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_304
timestamp 1621261055
transform 1 0 30336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_312
timestamp 1621261055
transform 1 0 31104 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_904
timestamp 1621261055
transform 1 0 32832 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_320
timestamp 1621261055
transform 1 0 31872 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_328
timestamp 1621261055
transform 1 0 32640 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_331
timestamp 1621261055
transform 1 0 32928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_320
timestamp 1621261055
transform 1 0 31872 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_328
timestamp 1621261055
transform 1 0 32640 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_336
timestamp 1621261055
transform 1 0 33408 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_339
timestamp 1621261055
transform 1 0 33696 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_347
timestamp 1621261055
transform 1 0 34464 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_355
timestamp 1621261055
transform 1 0 35232 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_344
timestamp 1621261055
transform 1 0 34176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_352
timestamp 1621261055
transform 1 0 34944 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_356
timestamp 1621261055
transform 1 0 35328 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_915
timestamp 1621261055
transform 1 0 35520 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_363
timestamp 1621261055
transform 1 0 36000 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_371
timestamp 1621261055
transform 1 0 36768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_359
timestamp 1621261055
transform 1 0 35616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_367
timestamp 1621261055
transform 1 0 36384 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_375
timestamp 1621261055
transform 1 0 37152 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_905
timestamp 1621261055
transform 1 0 38112 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_379
timestamp 1621261055
transform 1 0 37536 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_383
timestamp 1621261055
transform 1 0 37920 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_386
timestamp 1621261055
transform 1 0 38208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_394
timestamp 1621261055
transform 1 0 38976 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_383
timestamp 1621261055
transform 1 0 37920 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_391
timestamp 1621261055
transform 1 0 38688 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_399
timestamp 1621261055
transform 1 0 39456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_916
timestamp 1621261055
transform 1 0 40800 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_152
timestamp 1621261055
transform -1 0 41568 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_402
timestamp 1621261055
transform 1 0 39744 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_410
timestamp 1621261055
transform 1 0 40512 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_418
timestamp 1621261055
transform 1 0 41280 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_70_407
timestamp 1621261055
transform 1 0 40224 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_411
timestamp 1621261055
transform 1 0 40608 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_414
timestamp 1621261055
transform 1 0 40896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _087_
timestamp 1621261055
transform -1 0 41856 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_906
timestamp 1621261055
transform 1 0 43392 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_424
timestamp 1621261055
transform 1 0 41856 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_432
timestamp 1621261055
transform 1 0 42624 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_441
timestamp 1621261055
transform 1 0 43488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_422
timestamp 1621261055
transform 1 0 41664 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_430
timestamp 1621261055
transform 1 0 42432 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_438
timestamp 1621261055
transform 1 0 43200 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _178_
timestamp 1621261055
transform 1 0 45024 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_120
timestamp 1621261055
transform 1 0 44832 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_449
timestamp 1621261055
transform 1 0 44256 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_457
timestamp 1621261055
transform 1 0 45024 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_446
timestamp 1621261055
transform 1 0 43968 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_70_454
timestamp 1621261055
transform 1 0 44736 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_460
timestamp 1621261055
transform 1 0 45312 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_917
timestamp 1621261055
transform 1 0 46080 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_465
timestamp 1621261055
transform 1 0 45792 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_473
timestamp 1621261055
transform 1 0 46560 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_481
timestamp 1621261055
transform 1 0 47328 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_469
timestamp 1621261055
transform 1 0 46176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_477
timestamp 1621261055
transform 1 0 46944 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_492
timestamp 1621261055
transform 1 0 48384 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_485
timestamp 1621261055
transform 1 0 47712 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_489
timestamp 1621261055
transform 1 0 48096 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_229
timestamp 1621261055
transform -1 0 48096 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _215_
timestamp 1621261055
transform -1 0 48384 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_500
timestamp 1621261055
transform 1 0 49152 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_496
timestamp 1621261055
transform 1 0 48768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_493
timestamp 1621261055
transform 1 0 48480 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_907
timestamp 1621261055
transform 1 0 48672 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_504
timestamp 1621261055
transform 1 0 49536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_918
timestamp 1621261055
transform 1 0 51360 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_512
timestamp 1621261055
transform 1 0 50304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_520
timestamp 1621261055
transform 1 0 51072 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_508
timestamp 1621261055
transform 1 0 49920 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_516
timestamp 1621261055
transform 1 0 50688 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_520
timestamp 1621261055
transform 1 0 51072 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_70_522
timestamp 1621261055
transform 1 0 51264 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_524
timestamp 1621261055
transform 1 0 51456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_528
timestamp 1621261055
transform 1 0 51840 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_536
timestamp 1621261055
transform 1 0 52608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_544
timestamp 1621261055
transform 1 0 53376 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_532
timestamp 1621261055
transform 1 0 52224 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_540
timestamp 1621261055
transform 1 0 52992 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_908
timestamp 1621261055
transform 1 0 53952 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_548
timestamp 1621261055
transform 1 0 53760 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_551
timestamp 1621261055
transform 1 0 54048 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_559
timestamp 1621261055
transform 1 0 54816 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_567
timestamp 1621261055
transform 1 0 55584 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_548
timestamp 1621261055
transform 1 0 53760 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_556
timestamp 1621261055
transform 1 0 54528 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_564
timestamp 1621261055
transform 1 0 55296 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_919
timestamp 1621261055
transform 1 0 56640 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_575
timestamp 1621261055
transform 1 0 56352 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_583
timestamp 1621261055
transform 1 0 57120 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_572
timestamp 1621261055
transform 1 0 56064 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_576
timestamp 1621261055
transform 1 0 56448 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_579
timestamp 1621261055
transform 1 0 56736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_587
timestamp 1621261055
transform 1 0 57504 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_139
timestamp 1621261055
transform -1 0 58848 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_141
timestamp 1621261055
transform -1 0 58848 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_69_591
timestamp 1621261055
transform 1 0 57888 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_595
timestamp 1621261055
transform 1 0 58272 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_595
timestamp 1621261055
transform 1 0 58272 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_142
timestamp 1621261055
transform 1 0 1152 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_71_4
timestamp 1621261055
transform 1 0 1536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_12
timestamp 1621261055
transform 1 0 2304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_20
timestamp 1621261055
transform 1 0 3072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _056_
timestamp 1621261055
transform 1 0 3936 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_71_28
timestamp 1621261055
transform 1 0 3840 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_32
timestamp 1621261055
transform 1 0 4224 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_40
timestamp 1621261055
transform 1 0 4992 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_920
timestamp 1621261055
transform 1 0 6432 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_48
timestamp 1621261055
transform 1 0 5760 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_52
timestamp 1621261055
transform 1 0 6144 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_54
timestamp 1621261055
transform 1 0 6336 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_56
timestamp 1621261055
transform 1 0 6528 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_64
timestamp 1621261055
transform 1 0 7296 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_72
timestamp 1621261055
transform 1 0 8064 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_80
timestamp 1621261055
transform 1 0 8832 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_88
timestamp 1621261055
transform 1 0 9600 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_96
timestamp 1621261055
transform 1 0 10368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_104
timestamp 1621261055
transform 1 0 11136 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_921
timestamp 1621261055
transform 1 0 11712 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_108
timestamp 1621261055
transform 1 0 11520 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_111
timestamp 1621261055
transform 1 0 11808 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_119
timestamp 1621261055
transform 1 0 12576 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_127
timestamp 1621261055
transform 1 0 13344 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_135
timestamp 1621261055
transform 1 0 14112 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_143
timestamp 1621261055
transform 1 0 14880 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_922
timestamp 1621261055
transform 1 0 16992 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_151
timestamp 1621261055
transform 1 0 15648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_159
timestamp 1621261055
transform 1 0 16416 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_163
timestamp 1621261055
transform 1 0 16800 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_166
timestamp 1621261055
transform 1 0 17088 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_174
timestamp 1621261055
transform 1 0 17856 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_182
timestamp 1621261055
transform 1 0 18624 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_190
timestamp 1621261055
transform 1 0 19392 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_198
timestamp 1621261055
transform 1 0 20160 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_206
timestamp 1621261055
transform 1 0 20928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_923
timestamp 1621261055
transform 1 0 22272 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_214
timestamp 1621261055
transform 1 0 21696 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_218
timestamp 1621261055
transform 1 0 22080 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_221
timestamp 1621261055
transform 1 0 22368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_229
timestamp 1621261055
transform 1 0 23136 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_237
timestamp 1621261055
transform 1 0 23904 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_245
timestamp 1621261055
transform 1 0 24672 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_253
timestamp 1621261055
transform 1 0 25440 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_261
timestamp 1621261055
transform 1 0 26208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_269
timestamp 1621261055
transform 1 0 26976 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_273
timestamp 1621261055
transform 1 0 27360 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_924
timestamp 1621261055
transform 1 0 27552 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_276
timestamp 1621261055
transform 1 0 27648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_284
timestamp 1621261055
transform 1 0 28416 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_292
timestamp 1621261055
transform 1 0 29184 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_300
timestamp 1621261055
transform 1 0 29952 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_308
timestamp 1621261055
transform 1 0 30720 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_925
timestamp 1621261055
transform 1 0 32832 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_316
timestamp 1621261055
transform 1 0 31488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_324
timestamp 1621261055
transform 1 0 32256 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_328
timestamp 1621261055
transform 1 0 32640 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_331
timestamp 1621261055
transform 1 0 32928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_339
timestamp 1621261055
transform 1 0 33696 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_347
timestamp 1621261055
transform 1 0 34464 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_355
timestamp 1621261055
transform 1 0 35232 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_363
timestamp 1621261055
transform 1 0 36000 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_371
timestamp 1621261055
transform 1 0 36768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_926
timestamp 1621261055
transform 1 0 38112 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_379
timestamp 1621261055
transform 1 0 37536 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_383
timestamp 1621261055
transform 1 0 37920 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_386
timestamp 1621261055
transform 1 0 38208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_394
timestamp 1621261055
transform 1 0 38976 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _096_
timestamp 1621261055
transform -1 0 41184 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_168
timestamp 1621261055
transform -1 0 40896 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_402
timestamp 1621261055
transform 1 0 39744 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_410
timestamp 1621261055
transform 1 0 40512 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_417
timestamp 1621261055
transform 1 0 41184 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_927
timestamp 1621261055
transform 1 0 43392 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_425
timestamp 1621261055
transform 1 0 41952 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_433
timestamp 1621261055
transform 1 0 42720 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_437
timestamp 1621261055
transform 1 0 43104 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_439
timestamp 1621261055
transform 1 0 43296 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_441
timestamp 1621261055
transform 1 0 43488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_449
timestamp 1621261055
transform 1 0 44256 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_457
timestamp 1621261055
transform 1 0 45024 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_465
timestamp 1621261055
transform 1 0 45792 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_473
timestamp 1621261055
transform 1 0 46560 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_481
timestamp 1621261055
transform 1 0 47328 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_928
timestamp 1621261055
transform 1 0 48672 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_489
timestamp 1621261055
transform 1 0 48096 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_493
timestamp 1621261055
transform 1 0 48480 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_496
timestamp 1621261055
transform 1 0 48768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_504
timestamp 1621261055
transform 1 0 49536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_512
timestamp 1621261055
transform 1 0 50304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_520
timestamp 1621261055
transform 1 0 51072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_528
timestamp 1621261055
transform 1 0 51840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_536
timestamp 1621261055
transform 1 0 52608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_544
timestamp 1621261055
transform 1 0 53376 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_929
timestamp 1621261055
transform 1 0 53952 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_548
timestamp 1621261055
transform 1 0 53760 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_551
timestamp 1621261055
transform 1 0 54048 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_559
timestamp 1621261055
transform 1 0 54816 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_567
timestamp 1621261055
transform 1 0 55584 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_575
timestamp 1621261055
transform 1 0 56352 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_583
timestamp 1621261055
transform 1 0 57120 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_143
timestamp 1621261055
transform -1 0 58848 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_71_591
timestamp 1621261055
transform 1 0 57888 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_595
timestamp 1621261055
transform 1 0 58272 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_144
timestamp 1621261055
transform 1 0 1152 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_72_4
timestamp 1621261055
transform 1 0 1536 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_12
timestamp 1621261055
transform 1 0 2304 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_20
timestamp 1621261055
transform 1 0 3072 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_930
timestamp 1621261055
transform 1 0 3840 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_29
timestamp 1621261055
transform 1 0 3936 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_37
timestamp 1621261055
transform 1 0 4704 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_45
timestamp 1621261055
transform 1 0 5472 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_53
timestamp 1621261055
transform 1 0 6240 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_61
timestamp 1621261055
transform 1 0 7008 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_931
timestamp 1621261055
transform 1 0 9120 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_69
timestamp 1621261055
transform 1 0 7776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_77
timestamp 1621261055
transform 1 0 8544 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_81
timestamp 1621261055
transform 1 0 8928 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_84
timestamp 1621261055
transform 1 0 9216 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_92
timestamp 1621261055
transform 1 0 9984 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_100
timestamp 1621261055
transform 1 0 10752 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _020_
timestamp 1621261055
transform 1 0 12480 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_72_108
timestamp 1621261055
transform 1 0 11520 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_116
timestamp 1621261055
transform 1 0 12288 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_121
timestamp 1621261055
transform 1 0 12768 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_932
timestamp 1621261055
transform 1 0 14400 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_129
timestamp 1621261055
transform 1 0 13536 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_72_137
timestamp 1621261055
transform 1 0 14304 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_139
timestamp 1621261055
transform 1 0 14496 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_147
timestamp 1621261055
transform 1 0 15264 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_155
timestamp 1621261055
transform 1 0 16032 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_163
timestamp 1621261055
transform 1 0 16800 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_171
timestamp 1621261055
transform 1 0 17568 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_179
timestamp 1621261055
transform 1 0 18336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_187
timestamp 1621261055
transform 1 0 19104 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_933
timestamp 1621261055
transform 1 0 19680 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_191
timestamp 1621261055
transform 1 0 19488 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_194
timestamp 1621261055
transform 1 0 19776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_202
timestamp 1621261055
transform 1 0 20544 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_210
timestamp 1621261055
transform 1 0 21312 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_218
timestamp 1621261055
transform 1 0 22080 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_226
timestamp 1621261055
transform 1 0 22848 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_934
timestamp 1621261055
transform 1 0 24960 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_234
timestamp 1621261055
transform 1 0 23616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_242
timestamp 1621261055
transform 1 0 24384 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_246
timestamp 1621261055
transform 1 0 24768 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_249
timestamp 1621261055
transform 1 0 25056 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_257
timestamp 1621261055
transform 1 0 25824 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_265
timestamp 1621261055
transform 1 0 26592 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_273
timestamp 1621261055
transform 1 0 27360 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_281
timestamp 1621261055
transform 1 0 28128 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_289
timestamp 1621261055
transform 1 0 28896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_935
timestamp 1621261055
transform 1 0 30240 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_297
timestamp 1621261055
transform 1 0 29664 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_301
timestamp 1621261055
transform 1 0 30048 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_304
timestamp 1621261055
transform 1 0 30336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_312
timestamp 1621261055
transform 1 0 31104 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _022_
timestamp 1621261055
transform 1 0 31968 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_72_320
timestamp 1621261055
transform 1 0 31872 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_324
timestamp 1621261055
transform 1 0 32256 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_332
timestamp 1621261055
transform 1 0 33024 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_340
timestamp 1621261055
transform 1 0 33792 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_348
timestamp 1621261055
transform 1 0 34560 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_356
timestamp 1621261055
transform 1 0 35328 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _182_
timestamp 1621261055
transform 1 0 37440 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_936
timestamp 1621261055
transform 1 0 35520 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_125
timestamp 1621261055
transform 1 0 37248 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_359
timestamp 1621261055
transform 1 0 35616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_367
timestamp 1621261055
transform 1 0 36384 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_72_375
timestamp 1621261055
transform 1 0 37152 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_381
timestamp 1621261055
transform 1 0 37728 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_389
timestamp 1621261055
transform 1 0 38496 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_397
timestamp 1621261055
transform 1 0 39264 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_937
timestamp 1621261055
transform 1 0 40800 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_405
timestamp 1621261055
transform 1 0 40032 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_414
timestamp 1621261055
transform 1 0 40896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_422
timestamp 1621261055
transform 1 0 41664 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_430
timestamp 1621261055
transform 1 0 42432 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_438
timestamp 1621261055
transform 1 0 43200 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_446
timestamp 1621261055
transform 1 0 43968 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_454
timestamp 1621261055
transform 1 0 44736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_462
timestamp 1621261055
transform 1 0 45504 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_938
timestamp 1621261055
transform 1 0 46080 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_466
timestamp 1621261055
transform 1 0 45888 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_469
timestamp 1621261055
transform 1 0 46176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_477
timestamp 1621261055
transform 1 0 46944 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_485
timestamp 1621261055
transform 1 0 47712 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_493
timestamp 1621261055
transform 1 0 48480 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_501
timestamp 1621261055
transform 1 0 49248 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_939
timestamp 1621261055
transform 1 0 51360 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_509
timestamp 1621261055
transform 1 0 50016 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_517
timestamp 1621261055
transform 1 0 50784 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_521
timestamp 1621261055
transform 1 0 51168 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_524
timestamp 1621261055
transform 1 0 51456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_532
timestamp 1621261055
transform 1 0 52224 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_540
timestamp 1621261055
transform 1 0 52992 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_548
timestamp 1621261055
transform 1 0 53760 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_556
timestamp 1621261055
transform 1 0 54528 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_564
timestamp 1621261055
transform 1 0 55296 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _147_
timestamp 1621261055
transform -1 0 57408 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_940
timestamp 1621261055
transform 1 0 56640 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_206
timestamp 1621261055
transform -1 0 57120 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_72_572
timestamp 1621261055
transform 1 0 56064 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_576
timestamp 1621261055
transform 1 0 56448 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_579
timestamp 1621261055
transform 1 0 56736 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_586
timestamp 1621261055
transform 1 0 57408 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_145
timestamp 1621261055
transform -1 0 58848 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_594
timestamp 1621261055
transform 1 0 58176 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_72_596
timestamp 1621261055
transform 1 0 58368 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _086_
timestamp 1621261055
transform 1 0 2592 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_146
timestamp 1621261055
transform 1 0 1152 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_150
timestamp 1621261055
transform 1 0 2400 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_4
timestamp 1621261055
transform 1 0 1536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_73_12
timestamp 1621261055
transform 1 0 2304 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_18
timestamp 1621261055
transform 1 0 2880 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_26
timestamp 1621261055
transform 1 0 3648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_34
timestamp 1621261055
transform 1 0 4416 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_42
timestamp 1621261055
transform 1 0 5184 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_941
timestamp 1621261055
transform 1 0 6432 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_50
timestamp 1621261055
transform 1 0 5952 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_73_54
timestamp 1621261055
transform 1 0 6336 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_56
timestamp 1621261055
transform 1 0 6528 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_64
timestamp 1621261055
transform 1 0 7296 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_72
timestamp 1621261055
transform 1 0 8064 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_80
timestamp 1621261055
transform 1 0 8832 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_88
timestamp 1621261055
transform 1 0 9600 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_96
timestamp 1621261055
transform 1 0 10368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_104
timestamp 1621261055
transform 1 0 11136 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_942
timestamp 1621261055
transform 1 0 11712 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_108
timestamp 1621261055
transform 1 0 11520 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_111
timestamp 1621261055
transform 1 0 11808 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_119
timestamp 1621261055
transform 1 0 12576 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_127
timestamp 1621261055
transform 1 0 13344 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_135
timestamp 1621261055
transform 1 0 14112 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_143
timestamp 1621261055
transform 1 0 14880 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_943
timestamp 1621261055
transform 1 0 16992 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_151
timestamp 1621261055
transform 1 0 15648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_159
timestamp 1621261055
transform 1 0 16416 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_163
timestamp 1621261055
transform 1 0 16800 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_166
timestamp 1621261055
transform 1 0 17088 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_174
timestamp 1621261055
transform 1 0 17856 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_182
timestamp 1621261055
transform 1 0 18624 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_190
timestamp 1621261055
transform 1 0 19392 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_198
timestamp 1621261055
transform 1 0 20160 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_206
timestamp 1621261055
transform 1 0 20928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_944
timestamp 1621261055
transform 1 0 22272 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_214
timestamp 1621261055
transform 1 0 21696 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_218
timestamp 1621261055
transform 1 0 22080 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_221
timestamp 1621261055
transform 1 0 22368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_229
timestamp 1621261055
transform 1 0 23136 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_237
timestamp 1621261055
transform 1 0 23904 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_245
timestamp 1621261055
transform 1 0 24672 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_253
timestamp 1621261055
transform 1 0 25440 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_261
timestamp 1621261055
transform 1 0 26208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_269
timestamp 1621261055
transform 1 0 26976 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_273
timestamp 1621261055
transform 1 0 27360 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_945
timestamp 1621261055
transform 1 0 27552 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_276
timestamp 1621261055
transform 1 0 27648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_284
timestamp 1621261055
transform 1 0 28416 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_292
timestamp 1621261055
transform 1 0 29184 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_300
timestamp 1621261055
transform 1 0 29952 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_308
timestamp 1621261055
transform 1 0 30720 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_946
timestamp 1621261055
transform 1 0 32832 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_316
timestamp 1621261055
transform 1 0 31488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_324
timestamp 1621261055
transform 1 0 32256 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_328
timestamp 1621261055
transform 1 0 32640 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_331
timestamp 1621261055
transform 1 0 32928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_339
timestamp 1621261055
transform 1 0 33696 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_347
timestamp 1621261055
transform 1 0 34464 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_355
timestamp 1621261055
transform 1 0 35232 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_363
timestamp 1621261055
transform 1 0 36000 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_371
timestamp 1621261055
transform 1 0 36768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_947
timestamp 1621261055
transform 1 0 38112 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_379
timestamp 1621261055
transform 1 0 37536 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_383
timestamp 1621261055
transform 1 0 37920 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_386
timestamp 1621261055
transform 1 0 38208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_394
timestamp 1621261055
transform 1 0 38976 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_402
timestamp 1621261055
transform 1 0 39744 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_410
timestamp 1621261055
transform 1 0 40512 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_418
timestamp 1621261055
transform 1 0 41280 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_948
timestamp 1621261055
transform 1 0 43392 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_426
timestamp 1621261055
transform 1 0 42048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_434
timestamp 1621261055
transform 1 0 42816 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_438
timestamp 1621261055
transform 1 0 43200 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_73_441
timestamp 1621261055
transform 1 0 43488 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _014_
timestamp 1621261055
transform 1 0 43872 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_73_448
timestamp 1621261055
transform 1 0 44160 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_456
timestamp 1621261055
transform 1 0 44928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_464
timestamp 1621261055
transform 1 0 45696 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_472
timestamp 1621261055
transform 1 0 46464 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_480
timestamp 1621261055
transform 1 0 47232 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_949
timestamp 1621261055
transform 1 0 48672 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_488
timestamp 1621261055
transform 1 0 48000 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_492
timestamp 1621261055
transform 1 0 48384 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_494
timestamp 1621261055
transform 1 0 48576 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_496
timestamp 1621261055
transform 1 0 48768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_504
timestamp 1621261055
transform 1 0 49536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_512
timestamp 1621261055
transform 1 0 50304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_520
timestamp 1621261055
transform 1 0 51072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_528
timestamp 1621261055
transform 1 0 51840 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_536
timestamp 1621261055
transform 1 0 52608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_544
timestamp 1621261055
transform 1 0 53376 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_950
timestamp 1621261055
transform 1 0 53952 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_548
timestamp 1621261055
transform 1 0 53760 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_551
timestamp 1621261055
transform 1 0 54048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_559
timestamp 1621261055
transform 1 0 54816 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_567
timestamp 1621261055
transform 1 0 55584 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_575
timestamp 1621261055
transform 1 0 56352 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_583
timestamp 1621261055
transform 1 0 57120 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_147
timestamp 1621261055
transform -1 0 58848 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_73_591
timestamp 1621261055
transform 1 0 57888 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_595
timestamp 1621261055
transform 1 0 58272 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_148
timestamp 1621261055
transform 1 0 1152 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_74_4
timestamp 1621261055
transform 1 0 1536 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_12
timestamp 1621261055
transform 1 0 2304 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_20
timestamp 1621261055
transform 1 0 3072 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_951
timestamp 1621261055
transform 1 0 3840 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_29
timestamp 1621261055
transform 1 0 3936 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_37
timestamp 1621261055
transform 1 0 4704 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_45
timestamp 1621261055
transform 1 0 5472 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_53
timestamp 1621261055
transform 1 0 6240 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_61
timestamp 1621261055
transform 1 0 7008 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_952
timestamp 1621261055
transform 1 0 9120 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_69
timestamp 1621261055
transform 1 0 7776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_77
timestamp 1621261055
transform 1 0 8544 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_81
timestamp 1621261055
transform 1 0 8928 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_84
timestamp 1621261055
transform 1 0 9216 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_92
timestamp 1621261055
transform 1 0 9984 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_100
timestamp 1621261055
transform 1 0 10752 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_108
timestamp 1621261055
transform 1 0 11520 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_116
timestamp 1621261055
transform 1 0 12288 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_124
timestamp 1621261055
transform 1 0 13056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_953
timestamp 1621261055
transform 1 0 14400 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_132
timestamp 1621261055
transform 1 0 13824 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_136
timestamp 1621261055
transform 1 0 14208 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_139
timestamp 1621261055
transform 1 0 14496 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_147
timestamp 1621261055
transform 1 0 15264 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_155
timestamp 1621261055
transform 1 0 16032 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_163
timestamp 1621261055
transform 1 0 16800 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_171
timestamp 1621261055
transform 1 0 17568 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_179
timestamp 1621261055
transform 1 0 18336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_187
timestamp 1621261055
transform 1 0 19104 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_954
timestamp 1621261055
transform 1 0 19680 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_191
timestamp 1621261055
transform 1 0 19488 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_194
timestamp 1621261055
transform 1 0 19776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_202
timestamp 1621261055
transform 1 0 20544 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_210
timestamp 1621261055
transform 1 0 21312 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_218
timestamp 1621261055
transform 1 0 22080 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_226
timestamp 1621261055
transform 1 0 22848 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_955
timestamp 1621261055
transform 1 0 24960 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_234
timestamp 1621261055
transform 1 0 23616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_242
timestamp 1621261055
transform 1 0 24384 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_246
timestamp 1621261055
transform 1 0 24768 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_249
timestamp 1621261055
transform 1 0 25056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_257
timestamp 1621261055
transform 1 0 25824 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_265
timestamp 1621261055
transform 1 0 26592 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_273
timestamp 1621261055
transform 1 0 27360 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_281
timestamp 1621261055
transform 1 0 28128 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_289
timestamp 1621261055
transform 1 0 28896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_956
timestamp 1621261055
transform 1 0 30240 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_297
timestamp 1621261055
transform 1 0 29664 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_301
timestamp 1621261055
transform 1 0 30048 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_304
timestamp 1621261055
transform 1 0 30336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_312
timestamp 1621261055
transform 1 0 31104 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_320
timestamp 1621261055
transform 1 0 31872 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_328
timestamp 1621261055
transform 1 0 32640 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_336
timestamp 1621261055
transform 1 0 33408 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_344
timestamp 1621261055
transform 1 0 34176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_352
timestamp 1621261055
transform 1 0 34944 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_356
timestamp 1621261055
transform 1 0 35328 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_957
timestamp 1621261055
transform 1 0 35520 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_359
timestamp 1621261055
transform 1 0 35616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_367
timestamp 1621261055
transform 1 0 36384 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_375
timestamp 1621261055
transform 1 0 37152 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_383
timestamp 1621261055
transform 1 0 37920 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_391
timestamp 1621261055
transform 1 0 38688 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_399
timestamp 1621261055
transform 1 0 39456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_958
timestamp 1621261055
transform 1 0 40800 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_407
timestamp 1621261055
transform 1 0 40224 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_411
timestamp 1621261055
transform 1 0 40608 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_414
timestamp 1621261055
transform 1 0 40896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_422
timestamp 1621261055
transform 1 0 41664 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_430
timestamp 1621261055
transform 1 0 42432 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_438
timestamp 1621261055
transform 1 0 43200 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_446
timestamp 1621261055
transform 1 0 43968 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_454
timestamp 1621261055
transform 1 0 44736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_462
timestamp 1621261055
transform 1 0 45504 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_959
timestamp 1621261055
transform 1 0 46080 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_466
timestamp 1621261055
transform 1 0 45888 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_469
timestamp 1621261055
transform 1 0 46176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_477
timestamp 1621261055
transform 1 0 46944 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_485
timestamp 1621261055
transform 1 0 47712 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_493
timestamp 1621261055
transform 1 0 48480 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_501
timestamp 1621261055
transform 1 0 49248 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_960
timestamp 1621261055
transform 1 0 51360 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_509
timestamp 1621261055
transform 1 0 50016 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_517
timestamp 1621261055
transform 1 0 50784 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_521
timestamp 1621261055
transform 1 0 51168 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_524
timestamp 1621261055
transform 1 0 51456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_532
timestamp 1621261055
transform 1 0 52224 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_540
timestamp 1621261055
transform 1 0 52992 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_548
timestamp 1621261055
transform 1 0 53760 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_556
timestamp 1621261055
transform 1 0 54528 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_564
timestamp 1621261055
transform 1 0 55296 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_961
timestamp 1621261055
transform 1 0 56640 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_572
timestamp 1621261055
transform 1 0 56064 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_576
timestamp 1621261055
transform 1 0 56448 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_579
timestamp 1621261055
transform 1 0 56736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_587
timestamp 1621261055
transform 1 0 57504 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_149
timestamp 1621261055
transform -1 0 58848 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_595
timestamp 1621261055
transform 1 0 58272 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _062_
timestamp 1621261055
transform 1 0 1824 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_150
timestamp 1621261055
transform 1 0 1152 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_180
timestamp 1621261055
transform 1 0 1632 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_4
timestamp 1621261055
transform 1 0 1536 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_10
timestamp 1621261055
transform 1 0 2112 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_18
timestamp 1621261055
transform 1 0 2880 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_26
timestamp 1621261055
transform 1 0 3648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_34
timestamp 1621261055
transform 1 0 4416 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_42
timestamp 1621261055
transform 1 0 5184 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_962
timestamp 1621261055
transform 1 0 6432 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_50
timestamp 1621261055
transform 1 0 5952 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_75_54
timestamp 1621261055
transform 1 0 6336 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_56
timestamp 1621261055
transform 1 0 6528 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_64
timestamp 1621261055
transform 1 0 7296 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_72
timestamp 1621261055
transform 1 0 8064 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_80
timestamp 1621261055
transform 1 0 8832 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_88
timestamp 1621261055
transform 1 0 9600 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_96
timestamp 1621261055
transform 1 0 10368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_104
timestamp 1621261055
transform 1 0 11136 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_963
timestamp 1621261055
transform 1 0 11712 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_108
timestamp 1621261055
transform 1 0 11520 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_111
timestamp 1621261055
transform 1 0 11808 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_119
timestamp 1621261055
transform 1 0 12576 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_127
timestamp 1621261055
transform 1 0 13344 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_135
timestamp 1621261055
transform 1 0 14112 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_143
timestamp 1621261055
transform 1 0 14880 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_964
timestamp 1621261055
transform 1 0 16992 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_151
timestamp 1621261055
transform 1 0 15648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_159
timestamp 1621261055
transform 1 0 16416 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_163
timestamp 1621261055
transform 1 0 16800 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_166
timestamp 1621261055
transform 1 0 17088 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_174
timestamp 1621261055
transform 1 0 17856 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_182
timestamp 1621261055
transform 1 0 18624 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_190
timestamp 1621261055
transform 1 0 19392 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_198
timestamp 1621261055
transform 1 0 20160 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_206
timestamp 1621261055
transform 1 0 20928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_965
timestamp 1621261055
transform 1 0 22272 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_214
timestamp 1621261055
transform 1 0 21696 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_218
timestamp 1621261055
transform 1 0 22080 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_221
timestamp 1621261055
transform 1 0 22368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_229
timestamp 1621261055
transform 1 0 23136 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_237
timestamp 1621261055
transform 1 0 23904 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_245
timestamp 1621261055
transform 1 0 24672 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_253
timestamp 1621261055
transform 1 0 25440 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_261
timestamp 1621261055
transform 1 0 26208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_269
timestamp 1621261055
transform 1 0 26976 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_273
timestamp 1621261055
transform 1 0 27360 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_966
timestamp 1621261055
transform 1 0 27552 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_276
timestamp 1621261055
transform 1 0 27648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_284
timestamp 1621261055
transform 1 0 28416 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_292
timestamp 1621261055
transform 1 0 29184 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _006_
timestamp 1621261055
transform 1 0 29952 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_75_303
timestamp 1621261055
transform 1 0 30240 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_311
timestamp 1621261055
transform 1 0 31008 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_967
timestamp 1621261055
transform 1 0 32832 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_319
timestamp 1621261055
transform 1 0 31776 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_327
timestamp 1621261055
transform 1 0 32544 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_329
timestamp 1621261055
transform 1 0 32736 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_331
timestamp 1621261055
transform 1 0 32928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_339
timestamp 1621261055
transform 1 0 33696 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_347
timestamp 1621261055
transform 1 0 34464 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_355
timestamp 1621261055
transform 1 0 35232 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_363
timestamp 1621261055
transform 1 0 36000 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_371
timestamp 1621261055
transform 1 0 36768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_968
timestamp 1621261055
transform 1 0 38112 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_379
timestamp 1621261055
transform 1 0 37536 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_383
timestamp 1621261055
transform 1 0 37920 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_386
timestamp 1621261055
transform 1 0 38208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_394
timestamp 1621261055
transform 1 0 38976 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_402
timestamp 1621261055
transform 1 0 39744 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_410
timestamp 1621261055
transform 1 0 40512 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_418
timestamp 1621261055
transform 1 0 41280 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_969
timestamp 1621261055
transform 1 0 43392 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_426
timestamp 1621261055
transform 1 0 42048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_434
timestamp 1621261055
transform 1 0 42816 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_438
timestamp 1621261055
transform 1 0 43200 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_441
timestamp 1621261055
transform 1 0 43488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_449
timestamp 1621261055
transform 1 0 44256 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_457
timestamp 1621261055
transform 1 0 45024 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_465
timestamp 1621261055
transform 1 0 45792 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_473
timestamp 1621261055
transform 1 0 46560 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_481
timestamp 1621261055
transform 1 0 47328 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_970
timestamp 1621261055
transform 1 0 48672 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_489
timestamp 1621261055
transform 1 0 48096 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_493
timestamp 1621261055
transform 1 0 48480 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_496
timestamp 1621261055
transform 1 0 48768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_504
timestamp 1621261055
transform 1 0 49536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _044_
timestamp 1621261055
transform 1 0 51264 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_75_512
timestamp 1621261055
transform 1 0 50304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_520
timestamp 1621261055
transform 1 0 51072 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_525
timestamp 1621261055
transform 1 0 51552 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_533
timestamp 1621261055
transform 1 0 52320 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_541
timestamp 1621261055
transform 1 0 53088 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_971
timestamp 1621261055
transform 1 0 53952 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_75_549
timestamp 1621261055
transform 1 0 53856 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_551
timestamp 1621261055
transform 1 0 54048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_559
timestamp 1621261055
transform 1 0 54816 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_567
timestamp 1621261055
transform 1 0 55584 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_575
timestamp 1621261055
transform 1 0 56352 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_583
timestamp 1621261055
transform 1 0 57120 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_151
timestamp 1621261055
transform -1 0 58848 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_75_591
timestamp 1621261055
transform 1 0 57888 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_595
timestamp 1621261055
transform 1 0 58272 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_152
timestamp 1621261055
transform 1 0 1152 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_76_4
timestamp 1621261055
transform 1 0 1536 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_12
timestamp 1621261055
transform 1 0 2304 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_20
timestamp 1621261055
transform 1 0 3072 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_972
timestamp 1621261055
transform 1 0 3840 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_29
timestamp 1621261055
transform 1 0 3936 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_37
timestamp 1621261055
transform 1 0 4704 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_45
timestamp 1621261055
transform 1 0 5472 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_53
timestamp 1621261055
transform 1 0 6240 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_61
timestamp 1621261055
transform 1 0 7008 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_973
timestamp 1621261055
transform 1 0 9120 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_69
timestamp 1621261055
transform 1 0 7776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_77
timestamp 1621261055
transform 1 0 8544 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_81
timestamp 1621261055
transform 1 0 8928 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_84
timestamp 1621261055
transform 1 0 9216 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_92
timestamp 1621261055
transform 1 0 9984 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_100
timestamp 1621261055
transform 1 0 10752 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_108
timestamp 1621261055
transform 1 0 11520 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_116
timestamp 1621261055
transform 1 0 12288 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_124
timestamp 1621261055
transform 1 0 13056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_974
timestamp 1621261055
transform 1 0 14400 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_132
timestamp 1621261055
transform 1 0 13824 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_136
timestamp 1621261055
transform 1 0 14208 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_139
timestamp 1621261055
transform 1 0 14496 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_147
timestamp 1621261055
transform 1 0 15264 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_155
timestamp 1621261055
transform 1 0 16032 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_163
timestamp 1621261055
transform 1 0 16800 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_171
timestamp 1621261055
transform 1 0 17568 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_179
timestamp 1621261055
transform 1 0 18336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_187
timestamp 1621261055
transform 1 0 19104 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_975
timestamp 1621261055
transform 1 0 19680 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_191
timestamp 1621261055
transform 1 0 19488 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_194
timestamp 1621261055
transform 1 0 19776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_202
timestamp 1621261055
transform 1 0 20544 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_210
timestamp 1621261055
transform 1 0 21312 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_218
timestamp 1621261055
transform 1 0 22080 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_226
timestamp 1621261055
transform 1 0 22848 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_976
timestamp 1621261055
transform 1 0 24960 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_234
timestamp 1621261055
transform 1 0 23616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_242
timestamp 1621261055
transform 1 0 24384 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_246
timestamp 1621261055
transform 1 0 24768 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_249
timestamp 1621261055
transform 1 0 25056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_257
timestamp 1621261055
transform 1 0 25824 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_265
timestamp 1621261055
transform 1 0 26592 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_273
timestamp 1621261055
transform 1 0 27360 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_281
timestamp 1621261055
transform 1 0 28128 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_289
timestamp 1621261055
transform 1 0 28896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_977
timestamp 1621261055
transform 1 0 30240 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_297
timestamp 1621261055
transform 1 0 29664 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_301
timestamp 1621261055
transform 1 0 30048 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_304
timestamp 1621261055
transform 1 0 30336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_312
timestamp 1621261055
transform 1 0 31104 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_320
timestamp 1621261055
transform 1 0 31872 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_328
timestamp 1621261055
transform 1 0 32640 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_336
timestamp 1621261055
transform 1 0 33408 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_344
timestamp 1621261055
transform 1 0 34176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_352
timestamp 1621261055
transform 1 0 34944 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_356
timestamp 1621261055
transform 1 0 35328 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_978
timestamp 1621261055
transform 1 0 35520 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_359
timestamp 1621261055
transform 1 0 35616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_367
timestamp 1621261055
transform 1 0 36384 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_375
timestamp 1621261055
transform 1 0 37152 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_383
timestamp 1621261055
transform 1 0 37920 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_391
timestamp 1621261055
transform 1 0 38688 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_399
timestamp 1621261055
transform 1 0 39456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_979
timestamp 1621261055
transform 1 0 40800 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_407
timestamp 1621261055
transform 1 0 40224 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_411
timestamp 1621261055
transform 1 0 40608 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_414
timestamp 1621261055
transform 1 0 40896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_422
timestamp 1621261055
transform 1 0 41664 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_430
timestamp 1621261055
transform 1 0 42432 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_438
timestamp 1621261055
transform 1 0 43200 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_446
timestamp 1621261055
transform 1 0 43968 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_454
timestamp 1621261055
transform 1 0 44736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_462
timestamp 1621261055
transform 1 0 45504 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_980
timestamp 1621261055
transform 1 0 46080 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_466
timestamp 1621261055
transform 1 0 45888 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_469
timestamp 1621261055
transform 1 0 46176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_477
timestamp 1621261055
transform 1 0 46944 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_485
timestamp 1621261055
transform 1 0 47712 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_493
timestamp 1621261055
transform 1 0 48480 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_501
timestamp 1621261055
transform 1 0 49248 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_981
timestamp 1621261055
transform 1 0 51360 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_509
timestamp 1621261055
transform 1 0 50016 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_517
timestamp 1621261055
transform 1 0 50784 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_521
timestamp 1621261055
transform 1 0 51168 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_524
timestamp 1621261055
transform 1 0 51456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_532
timestamp 1621261055
transform 1 0 52224 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_540
timestamp 1621261055
transform 1 0 52992 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_548
timestamp 1621261055
transform 1 0 53760 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_556
timestamp 1621261055
transform 1 0 54528 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_564
timestamp 1621261055
transform 1 0 55296 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_982
timestamp 1621261055
transform 1 0 56640 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_93
timestamp 1621261055
transform -1 0 57696 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_76_572
timestamp 1621261055
transform 1 0 56064 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_576
timestamp 1621261055
transform 1 0 56448 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_579
timestamp 1621261055
transform 1 0 56736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_153
timestamp 1621261055
transform -1 0 58848 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output436
timestamp 1621261055
transform -1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_94
timestamp 1621261055
transform -1 0 58272 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_595
timestamp 1621261055
transform 1 0 58272 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_154
timestamp 1621261055
transform 1 0 1152 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_156
timestamp 1621261055
transform 1 0 1152 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_4
timestamp 1621261055
transform 1 0 1536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_12
timestamp 1621261055
transform 1 0 2304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_20
timestamp 1621261055
transform 1 0 3072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_4
timestamp 1621261055
transform 1 0 1536 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_12
timestamp 1621261055
transform 1 0 2304 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_20
timestamp 1621261055
transform 1 0 3072 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_993
timestamp 1621261055
transform 1 0 3840 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_28
timestamp 1621261055
transform 1 0 3840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_36
timestamp 1621261055
transform 1 0 4608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_29
timestamp 1621261055
transform 1 0 3936 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_37
timestamp 1621261055
transform 1 0 4704 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_983
timestamp 1621261055
transform 1 0 6432 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_194
timestamp 1621261055
transform 1 0 7104 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_44
timestamp 1621261055
transform 1 0 5376 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_52
timestamp 1621261055
transform 1 0 6144 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_77_54
timestamp 1621261055
transform 1 0 6336 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_56
timestamp 1621261055
transform 1 0 6528 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_45
timestamp 1621261055
transform 1 0 5472 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_53
timestamp 1621261055
transform 1 0 6240 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_61
timestamp 1621261055
transform 1 0 7008 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _128_
timestamp 1621261055
transform 1 0 7296 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_994
timestamp 1621261055
transform 1 0 9120 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_64
timestamp 1621261055
transform 1 0 7296 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_72
timestamp 1621261055
transform 1 0 8064 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_80
timestamp 1621261055
transform 1 0 8832 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_67
timestamp 1621261055
transform 1 0 7584 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_75
timestamp 1621261055
transform 1 0 8352 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_84
timestamp 1621261055
transform 1 0 9216 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_88
timestamp 1621261055
transform 1 0 9600 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_96
timestamp 1621261055
transform 1 0 10368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_104
timestamp 1621261055
transform 1 0 11136 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_92
timestamp 1621261055
transform 1 0 9984 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_100
timestamp 1621261055
transform 1 0 10752 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_984
timestamp 1621261055
transform 1 0 11712 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_108
timestamp 1621261055
transform 1 0 11520 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_111
timestamp 1621261055
transform 1 0 11808 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_119
timestamp 1621261055
transform 1 0 12576 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_108
timestamp 1621261055
transform 1 0 11520 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_116
timestamp 1621261055
transform 1 0 12288 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_124
timestamp 1621261055
transform 1 0 13056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_995
timestamp 1621261055
transform 1 0 14400 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_127
timestamp 1621261055
transform 1 0 13344 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_135
timestamp 1621261055
transform 1 0 14112 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_143
timestamp 1621261055
transform 1 0 14880 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_132
timestamp 1621261055
transform 1 0 13824 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_136
timestamp 1621261055
transform 1 0 14208 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_139
timestamp 1621261055
transform 1 0 14496 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_147
timestamp 1621261055
transform 1 0 15264 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_985
timestamp 1621261055
transform 1 0 16992 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_151
timestamp 1621261055
transform 1 0 15648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_159
timestamp 1621261055
transform 1 0 16416 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_163
timestamp 1621261055
transform 1 0 16800 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_166
timestamp 1621261055
transform 1 0 17088 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_155
timestamp 1621261055
transform 1 0 16032 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_163
timestamp 1621261055
transform 1 0 16800 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_174
timestamp 1621261055
transform 1 0 17856 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_182
timestamp 1621261055
transform 1 0 18624 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_171
timestamp 1621261055
transform 1 0 17568 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_179
timestamp 1621261055
transform 1 0 18336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_187
timestamp 1621261055
transform 1 0 19104 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_78_196
timestamp 1621261055
transform 1 0 19968 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_194
timestamp 1621261055
transform 1 0 19776 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_191
timestamp 1621261055
transform 1 0 19488 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_190
timestamp 1621261055
transform 1 0 19392 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_178
timestamp 1621261055
transform 1 0 20064 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_996
timestamp 1621261055
transform 1 0 19680 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_202
timestamp 1621261055
transform 1 0 20544 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_206
timestamp 1621261055
transform 1 0 20928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_198
timestamp 1621261055
transform 1 0 20160 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _106_
timestamp 1621261055
transform 1 0 20256 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_210
timestamp 1621261055
transform 1 0 21312 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_218
timestamp 1621261055
transform 1 0 22080 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_218
timestamp 1621261055
transform 1 0 22080 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_214
timestamp 1621261055
transform 1 0 21696 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_226
timestamp 1621261055
transform 1 0 22848 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_220
timestamp 1621261055
transform 1 0 22272 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_221
timestamp 1621261055
transform 1 0 22368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_114
timestamp 1621261055
transform 1 0 22368 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_986
timestamp 1621261055
transform 1 0 22272 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _174_
timestamp 1621261055
transform 1 0 22560 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_77_229
timestamp 1621261055
transform 1 0 23136 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_997
timestamp 1621261055
transform 1 0 24960 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_237
timestamp 1621261055
transform 1 0 23904 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_245
timestamp 1621261055
transform 1 0 24672 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_234
timestamp 1621261055
transform 1 0 23616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_242
timestamp 1621261055
transform 1 0 24384 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_246
timestamp 1621261055
transform 1 0 24768 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_249
timestamp 1621261055
transform 1 0 25056 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _219_
timestamp 1621261055
transform 1 0 25440 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_77_253
timestamp 1621261055
transform 1 0 25440 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_261
timestamp 1621261055
transform 1 0 26208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_269
timestamp 1621261055
transform 1 0 26976 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_273
timestamp 1621261055
transform 1 0 27360 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_256
timestamp 1621261055
transform 1 0 25728 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_264
timestamp 1621261055
transform 1 0 26496 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_272
timestamp 1621261055
transform 1 0 27264 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_987
timestamp 1621261055
transform 1 0 27552 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_276
timestamp 1621261055
transform 1 0 27648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_284
timestamp 1621261055
transform 1 0 28416 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_292
timestamp 1621261055
transform 1 0 29184 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_280
timestamp 1621261055
transform 1 0 28032 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_288
timestamp 1621261055
transform 1 0 28800 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_998
timestamp 1621261055
transform 1 0 30240 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_300
timestamp 1621261055
transform 1 0 29952 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_308
timestamp 1621261055
transform 1 0 30720 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_296
timestamp 1621261055
transform 1 0 29568 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_300
timestamp 1621261055
transform 1 0 29952 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_78_302
timestamp 1621261055
transform 1 0 30144 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_304
timestamp 1621261055
transform 1 0 30336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_312
timestamp 1621261055
transform 1 0 31104 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_988
timestamp 1621261055
transform 1 0 32832 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_316
timestamp 1621261055
transform 1 0 31488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_324
timestamp 1621261055
transform 1 0 32256 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_328
timestamp 1621261055
transform 1 0 32640 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_331
timestamp 1621261055
transform 1 0 32928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_320
timestamp 1621261055
transform 1 0 31872 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_328
timestamp 1621261055
transform 1 0 32640 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_336
timestamp 1621261055
transform 1 0 33408 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_339
timestamp 1621261055
transform 1 0 33696 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_347
timestamp 1621261055
transform 1 0 34464 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_355
timestamp 1621261055
transform 1 0 35232 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_344
timestamp 1621261055
transform 1 0 34176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_352
timestamp 1621261055
transform 1 0 34944 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_356
timestamp 1621261055
transform 1 0 35328 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_999
timestamp 1621261055
transform 1 0 35520 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_363
timestamp 1621261055
transform 1 0 36000 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_371
timestamp 1621261055
transform 1 0 36768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_359
timestamp 1621261055
transform 1 0 35616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_367
timestamp 1621261055
transform 1 0 36384 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_375
timestamp 1621261055
transform 1 0 37152 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_989
timestamp 1621261055
transform 1 0 38112 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_77_379
timestamp 1621261055
transform 1 0 37536 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_383
timestamp 1621261055
transform 1 0 37920 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_386
timestamp 1621261055
transform 1 0 38208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_394
timestamp 1621261055
transform 1 0 38976 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_383
timestamp 1621261055
transform 1 0 37920 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_391
timestamp 1621261055
transform 1 0 38688 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_399
timestamp 1621261055
transform 1 0 39456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1000
timestamp 1621261055
transform 1 0 40800 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_402
timestamp 1621261055
transform 1 0 39744 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_410
timestamp 1621261055
transform 1 0 40512 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_418
timestamp 1621261055
transform 1 0 41280 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_407
timestamp 1621261055
transform 1 0 40224 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_411
timestamp 1621261055
transform 1 0 40608 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_414
timestamp 1621261055
transform 1 0 40896 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_426
timestamp 1621261055
transform 1 0 42048 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_422
timestamp 1621261055
transform 1 0 41664 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_426
timestamp 1621261055
transform 1 0 42048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _046_
timestamp 1621261055
transform 1 0 42144 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_430
timestamp 1621261055
transform 1 0 42432 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_434
timestamp 1621261055
transform 1 0 42816 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_438
timestamp 1621261055
transform 1 0 43200 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_441
timestamp 1621261055
transform 1 0 43488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_438
timestamp 1621261055
transform 1 0 43200 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_990
timestamp 1621261055
transform 1 0 43392 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_449
timestamp 1621261055
transform 1 0 44256 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_457
timestamp 1621261055
transform 1 0 45024 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_446
timestamp 1621261055
transform 1 0 43968 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_454
timestamp 1621261055
transform 1 0 44736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_462
timestamp 1621261055
transform 1 0 45504 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1001
timestamp 1621261055
transform 1 0 46080 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_465
timestamp 1621261055
transform 1 0 45792 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_473
timestamp 1621261055
transform 1 0 46560 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_481
timestamp 1621261055
transform 1 0 47328 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_466
timestamp 1621261055
transform 1 0 45888 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_469
timestamp 1621261055
transform 1 0 46176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_477
timestamp 1621261055
transform 1 0 46944 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_991
timestamp 1621261055
transform 1 0 48672 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_77_489
timestamp 1621261055
transform 1 0 48096 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_493
timestamp 1621261055
transform 1 0 48480 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_496
timestamp 1621261055
transform 1 0 48768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_504
timestamp 1621261055
transform 1 0 49536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_485
timestamp 1621261055
transform 1 0 47712 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_493
timestamp 1621261055
transform 1 0 48480 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_501
timestamp 1621261055
transform 1 0 49248 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1002
timestamp 1621261055
transform 1 0 51360 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_512
timestamp 1621261055
transform 1 0 50304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_520
timestamp 1621261055
transform 1 0 51072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_509
timestamp 1621261055
transform 1 0 50016 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_517
timestamp 1621261055
transform 1 0 50784 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_521
timestamp 1621261055
transform 1 0 51168 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_524
timestamp 1621261055
transform 1 0 51456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_528
timestamp 1621261055
transform 1 0 51840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_536
timestamp 1621261055
transform 1 0 52608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_544
timestamp 1621261055
transform 1 0 53376 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_532
timestamp 1621261055
transform 1 0 52224 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_540
timestamp 1621261055
transform 1 0 52992 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_992
timestamp 1621261055
transform 1 0 53952 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_548
timestamp 1621261055
transform 1 0 53760 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_551
timestamp 1621261055
transform 1 0 54048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_559
timestamp 1621261055
transform 1 0 54816 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_567
timestamp 1621261055
transform 1 0 55584 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_548
timestamp 1621261055
transform 1 0 53760 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_556
timestamp 1621261055
transform 1 0 54528 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_564
timestamp 1621261055
transform 1 0 55296 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1003
timestamp 1621261055
transform 1 0 56640 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_30
timestamp 1621261055
transform -1 0 57696 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_90
timestamp 1621261055
transform -1 0 57696 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_575
timestamp 1621261055
transform 1 0 56352 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_583
timestamp 1621261055
transform 1 0 57120 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_78_572
timestamp 1621261055
transform 1 0 56064 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_576
timestamp 1621261055
transform 1 0 56448 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_579
timestamp 1621261055
transform 1 0 56736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_155
timestamp 1621261055
transform -1 0 58848 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_157
timestamp 1621261055
transform -1 0 58848 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output398
timestamp 1621261055
transform -1 0 58080 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output435
timestamp 1621261055
transform -1 0 58080 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_91
timestamp 1621261055
transform -1 0 58272 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_595
timestamp 1621261055
transform 1 0 58272 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_593
timestamp 1621261055
transform 1 0 58080 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_158
timestamp 1621261055
transform 1 0 1152 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output406
timestamp 1621261055
transform 1 0 1536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_38
timestamp 1621261055
transform 1 0 1920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_10
timestamp 1621261055
transform 1 0 2112 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_18
timestamp 1621261055
transform 1 0 2880 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output428
timestamp 1621261055
transform 1 0 4320 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_79
timestamp 1621261055
transform 1 0 4128 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_26
timestamp 1621261055
transform 1 0 3648 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_30
timestamp 1621261055
transform 1 0 4032 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_37
timestamp 1621261055
transform 1 0 4704 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1004
timestamp 1621261055
transform 1 0 6432 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_45
timestamp 1621261055
transform 1 0 5472 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_53
timestamp 1621261055
transform 1 0 6240 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_56
timestamp 1621261055
transform 1 0 6528 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output438
timestamp 1621261055
transform 1 0 7488 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output439
timestamp 1621261055
transform -1 0 9504 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_98
timestamp 1621261055
transform 1 0 7296 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_100
timestamp 1621261055
transform -1 0 9120 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_70
timestamp 1621261055
transform 1 0 7872 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_78
timestamp 1621261055
transform 1 0 8640 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_80
timestamp 1621261055
transform 1 0 8832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_87
timestamp 1621261055
transform 1 0 9504 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_95
timestamp 1621261055
transform 1 0 10272 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_103
timestamp 1621261055
transform 1 0 11040 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1005
timestamp 1621261055
transform 1 0 11712 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_107
timestamp 1621261055
transform 1 0 11424 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_109
timestamp 1621261055
transform 1 0 11616 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_111
timestamp 1621261055
transform 1 0 11808 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_119
timestamp 1621261055
transform 1 0 12576 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output442
timestamp 1621261055
transform 1 0 13824 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_79_127
timestamp 1621261055
transform 1 0 13344 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_131
timestamp 1621261055
transform 1 0 13728 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_136
timestamp 1621261055
transform 1 0 14208 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_144
timestamp 1621261055
transform 1 0 14976 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1006
timestamp 1621261055
transform 1 0 16992 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_152
timestamp 1621261055
transform 1 0 15744 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_160
timestamp 1621261055
transform 1 0 16512 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_164
timestamp 1621261055
transform 1 0 16896 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_166
timestamp 1621261055
transform 1 0 17088 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_168
timestamp 1621261055
transform 1 0 17280 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _134_
timestamp 1621261055
transform 1 0 17568 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_199
timestamp 1621261055
transform 1 0 17376 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_174
timestamp 1621261055
transform 1 0 17856 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_182
timestamp 1621261055
transform 1 0 18624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _190_
timestamp 1621261055
transform -1 0 21216 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output409
timestamp 1621261055
transform -1 0 20544 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_44
timestamp 1621261055
transform -1 0 20160 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_233
timestamp 1621261055
transform -1 0 20928 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_190
timestamp 1621261055
transform 1 0 19392 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_194
timestamp 1621261055
transform 1 0 19776 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_202
timestamp 1621261055
transform 1 0 20544 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_209
timestamp 1621261055
transform 1 0 21216 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1007
timestamp 1621261055
transform 1 0 22272 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output411
timestamp 1621261055
transform 1 0 23328 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_48
timestamp 1621261055
transform 1 0 23136 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_217
timestamp 1621261055
transform 1 0 21984 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_219
timestamp 1621261055
transform 1 0 22176 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_221
timestamp 1621261055
transform 1 0 22368 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output412
timestamp 1621261055
transform -1 0 25248 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_50
timestamp 1621261055
transform -1 0 24864 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_235
timestamp 1621261055
transform 1 0 23712 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_243
timestamp 1621261055
transform 1 0 24480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_251
timestamp 1621261055
transform 1 0 25248 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_259
timestamp 1621261055
transform 1 0 26016 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_267
timestamp 1621261055
transform 1 0 26784 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1008
timestamp 1621261055
transform 1 0 27552 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_276
timestamp 1621261055
transform 1 0 27648 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_284
timestamp 1621261055
transform 1 0 28416 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_292
timestamp 1621261055
transform 1 0 29184 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_300
timestamp 1621261055
transform 1 0 29952 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_308
timestamp 1621261055
transform 1 0 30720 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1009
timestamp 1621261055
transform 1 0 32832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_316
timestamp 1621261055
transform 1 0 31488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_324
timestamp 1621261055
transform 1 0 32256 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_328
timestamp 1621261055
transform 1 0 32640 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_331
timestamp 1621261055
transform 1 0 32928 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_339
timestamp 1621261055
transform 1 0 33696 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_347
timestamp 1621261055
transform 1 0 34464 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_355
timestamp 1621261055
transform 1 0 35232 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_363
timestamp 1621261055
transform 1 0 36000 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_371
timestamp 1621261055
transform 1 0 36768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1010
timestamp 1621261055
transform 1 0 38112 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output422
timestamp 1621261055
transform -1 0 39456 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_67
timestamp 1621261055
transform -1 0 39072 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_379
timestamp 1621261055
transform 1 0 37536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_383
timestamp 1621261055
transform 1 0 37920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_386
timestamp 1621261055
transform 1 0 38208 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_390
timestamp 1621261055
transform 1 0 38592 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_392
timestamp 1621261055
transform 1 0 38784 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_399
timestamp 1621261055
transform 1 0 39456 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _075_
timestamp 1621261055
transform -1 0 40128 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output423
timestamp 1621261055
transform 1 0 40704 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_136
timestamp 1621261055
transform -1 0 39840 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_406
timestamp 1621261055
transform 1 0 40128 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_410
timestamp 1621261055
transform 1 0 40512 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_416
timestamp 1621261055
transform 1 0 41088 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1011
timestamp 1621261055
transform 1 0 43392 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_424
timestamp 1621261055
transform 1 0 41856 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_432
timestamp 1621261055
transform 1 0 42624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_441
timestamp 1621261055
transform 1 0 43488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output426
timestamp 1621261055
transform -1 0 45792 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_74
timestamp 1621261055
transform -1 0 45408 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_449
timestamp 1621261055
transform 1 0 44256 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_457
timestamp 1621261055
transform 1 0 45024 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _002_
timestamp 1621261055
transform 1 0 46272 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output427
timestamp 1621261055
transform -1 0 47328 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_75
timestamp 1621261055
transform -1 0 45984 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_77
timestamp 1621261055
transform -1 0 46944 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_467
timestamp 1621261055
transform 1 0 45984 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_469
timestamp 1621261055
transform 1 0 46176 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_473
timestamp 1621261055
transform 1 0 46560 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_481
timestamp 1621261055
transform 1 0 47328 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1012
timestamp 1621261055
transform 1 0 48672 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_79_489
timestamp 1621261055
transform 1 0 48096 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_493
timestamp 1621261055
transform 1 0 48480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_496
timestamp 1621261055
transform 1 0 48768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_504
timestamp 1621261055
transform 1 0 49536 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_512
timestamp 1621261055
transform 1 0 50304 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_520
timestamp 1621261055
transform 1 0 51072 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_524
timestamp 1621261055
transform 1 0 51456 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output431
timestamp 1621261055
transform 1 0 51744 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_526
timestamp 1621261055
transform 1 0 51648 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_531
timestamp 1621261055
transform 1 0 52128 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_539
timestamp 1621261055
transform 1 0 52896 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1013
timestamp 1621261055
transform 1 0 53952 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_172
timestamp 1621261055
transform -1 0 55776 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_547
timestamp 1621261055
transform 1 0 53664 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_549
timestamp 1621261055
transform 1 0 53856 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_551
timestamp 1621261055
transform 1 0 54048 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_559
timestamp 1621261055
transform 1 0 54816 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _061_
timestamp 1621261055
transform -1 0 56064 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output397
timestamp 1621261055
transform -1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output434
timestamp 1621261055
transform -1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_28
timestamp 1621261055
transform -1 0 57504 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_88
timestamp 1621261055
transform -1 0 56448 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_572
timestamp 1621261055
transform 1 0 56064 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_580
timestamp 1621261055
transform 1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_584
timestamp 1621261055
transform 1 0 57216 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_159
timestamp 1621261055
transform -1 0 58848 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_79_591
timestamp 1621261055
transform 1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_595
timestamp 1621261055
transform 1 0 58272 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_160
timestamp 1621261055
transform 1 0 1152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output368
timestamp 1621261055
transform 1 0 1536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output379
timestamp 1621261055
transform 1 0 2304 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output417
timestamp 1621261055
transform 1 0 3072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_11
timestamp 1621261055
transform 1 0 2112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_58
timestamp 1621261055
transform 1 0 2880 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_8
timestamp 1621261055
transform 1 0 1920 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_16
timestamp 1621261055
transform 1 0 2688 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1014
timestamp 1621261055
transform 1 0 3840 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output390
timestamp 1621261055
transform 1 0 4320 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_32
timestamp 1621261055
transform 1 0 5184 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_24
timestamp 1621261055
transform 1 0 3456 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_29
timestamp 1621261055
transform 1 0 3936 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_37
timestamp 1621261055
transform 1 0 4704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_41
timestamp 1621261055
transform 1 0 5088 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output399
timestamp 1621261055
transform 1 0 5376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output400
timestamp 1621261055
transform 1 0 7008 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output437
timestamp 1621261055
transform 1 0 6144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_96
timestamp 1621261055
transform 1 0 5952 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_48
timestamp 1621261055
transform 1 0 5760 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_56
timestamp 1621261055
transform 1 0 6528 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_60
timestamp 1621261055
transform 1 0 6912 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1015
timestamp 1621261055
transform 1 0 9120 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output401
timestamp 1621261055
transform 1 0 8352 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_34
timestamp 1621261055
transform 1 0 8160 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_65
timestamp 1621261055
transform 1 0 7392 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_79
timestamp 1621261055
transform 1 0 8736 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_84
timestamp 1621261055
transform 1 0 9216 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output402
timestamp 1621261055
transform 1 0 10176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output440
timestamp 1621261055
transform 1 0 10944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_102
timestamp 1621261055
transform 1 0 10752 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_92
timestamp 1621261055
transform 1 0 9984 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_98
timestamp 1621261055
transform 1 0 10560 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output403
timestamp 1621261055
transform 1 0 11712 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output441
timestamp 1621261055
transform 1 0 12480 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_36
timestamp 1621261055
transform 1 0 13152 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_106
timestamp 1621261055
transform 1 0 11328 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_114
timestamp 1621261055
transform 1 0 12096 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_122
timestamp 1621261055
transform 1 0 12864 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_124
timestamp 1621261055
transform 1 0 13056 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1016
timestamp 1621261055
transform 1 0 14400 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output404
timestamp 1621261055
transform 1 0 13344 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output405
timestamp 1621261055
transform 1 0 14880 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_131
timestamp 1621261055
transform 1 0 13728 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_135
timestamp 1621261055
transform 1 0 14112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_137
timestamp 1621261055
transform 1 0 14304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_139
timestamp 1621261055
transform 1 0 14496 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_147
timestamp 1621261055
transform 1 0 15264 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output407
timestamp 1621261055
transform 1 0 16992 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output443
timestamp 1621261055
transform -1 0 16032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_40
timestamp 1621261055
transform 1 0 16800 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_104
timestamp 1621261055
transform -1 0 15648 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_155
timestamp 1621261055
transform 1 0 16032 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output408
timestamp 1621261055
transform -1 0 18912 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_42
timestamp 1621261055
transform -1 0 18528 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_169
timestamp 1621261055
transform 1 0 17376 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_177
timestamp 1621261055
transform 1 0 18144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_185
timestamp 1621261055
transform 1 0 18912 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1017
timestamp 1621261055
transform 1 0 19680 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output371
timestamp 1621261055
transform 1 0 20160 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output372
timestamp 1621261055
transform 1 0 21216 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_5
timestamp 1621261055
transform 1 0 19968 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_7
timestamp 1621261055
transform 1 0 21024 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_194
timestamp 1621261055
transform 1 0 19776 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_202
timestamp 1621261055
transform 1 0 20544 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_206
timestamp 1621261055
transform 1 0 20928 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output373
timestamp 1621261055
transform 1 0 22752 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output410
timestamp 1621261055
transform -1 0 22368 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_46
timestamp 1621261055
transform -1 0 21984 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_213
timestamp 1621261055
transform 1 0 21600 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_221
timestamp 1621261055
transform 1 0 22368 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_229
timestamp 1621261055
transform 1 0 23136 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1018
timestamp 1621261055
transform 1 0 24960 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output374
timestamp 1621261055
transform 1 0 24192 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_237
timestamp 1621261055
transform 1 0 23904 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_239
timestamp 1621261055
transform 1 0 24096 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_244
timestamp 1621261055
transform 1 0 24576 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_249
timestamp 1621261055
transform 1 0 25056 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output375
timestamp 1621261055
transform 1 0 25920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output413
timestamp 1621261055
transform 1 0 26688 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_9
timestamp 1621261055
transform 1 0 27360 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_257
timestamp 1621261055
transform 1 0 25824 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_262
timestamp 1621261055
transform 1 0 26304 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_270
timestamp 1621261055
transform 1 0 27072 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_272
timestamp 1621261055
transform 1 0 27264 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output376
timestamp 1621261055
transform 1 0 27552 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output414
timestamp 1621261055
transform -1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_52
timestamp 1621261055
transform -1 0 28320 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_54
timestamp 1621261055
transform -1 0 29472 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_279
timestamp 1621261055
transform 1 0 27936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_287
timestamp 1621261055
transform 1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_291
timestamp 1621261055
transform 1 0 29088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1019
timestamp 1621261055
transform 1 0 30240 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output378
timestamp 1621261055
transform 1 0 30720 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output415
timestamp 1621261055
transform -1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_56
timestamp 1621261055
transform -1 0 31488 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_299
timestamp 1621261055
transform 1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_304
timestamp 1621261055
transform 1 0 30336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_312
timestamp 1621261055
transform 1 0 31104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output380
timestamp 1621261055
transform 1 0 32256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output416
timestamp 1621261055
transform -1 0 31872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output418
timestamp 1621261055
transform 1 0 33024 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_320
timestamp 1621261055
transform 1 0 31872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_328
timestamp 1621261055
transform 1 0 32640 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_336
timestamp 1621261055
transform 1 0 33408 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output381
timestamp 1621261055
transform 1 0 33792 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output419
timestamp 1621261055
transform 1 0 34560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_60
timestamp 1621261055
transform 1 0 34368 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_344
timestamp 1621261055
transform 1 0 34176 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_352
timestamp 1621261055
transform 1 0 34944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_356
timestamp 1621261055
transform 1 0 35328 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1020
timestamp 1621261055
transform 1 0 35520 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output382
timestamp 1621261055
transform 1 0 36000 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output420
timestamp 1621261055
transform -1 0 37152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_62
timestamp 1621261055
transform -1 0 36768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_64
timestamp 1621261055
transform -1 0 37536 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_359
timestamp 1621261055
transform 1 0 35616 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_367
timestamp 1621261055
transform 1 0 36384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_375
timestamp 1621261055
transform 1 0 37152 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output384
timestamp 1621261055
transform -1 0 38976 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output421
timestamp 1621261055
transform -1 0 37920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_16
timestamp 1621261055
transform -1 0 38592 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_65
timestamp 1621261055
transform -1 0 38112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_385
timestamp 1621261055
transform 1 0 38112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_387
timestamp 1621261055
transform 1 0 38304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_394
timestamp 1621261055
transform 1 0 38976 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1021
timestamp 1621261055
transform 1 0 40800 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output385
timestamp 1621261055
transform -1 0 40416 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_18
timestamp 1621261055
transform -1 0 40032 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_402
timestamp 1621261055
transform 1 0 39744 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_409
timestamp 1621261055
transform 1 0 40416 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_414
timestamp 1621261055
transform 1 0 40896 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_418
timestamp 1621261055
transform 1 0 41280 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_420
timestamp 1621261055
transform 1 0 41472 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output386
timestamp 1621261055
transform 1 0 41760 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output387
timestamp 1621261055
transform 1 0 43296 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output424
timestamp 1621261055
transform -1 0 42912 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_20
timestamp 1621261055
transform 1 0 41568 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_69
timestamp 1621261055
transform -1 0 42528 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_427
timestamp 1621261055
transform 1 0 42144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_435
timestamp 1621261055
transform 1 0 42912 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output388
timestamp 1621261055
transform 1 0 44928 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output425
timestamp 1621261055
transform -1 0 44448 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_71
timestamp 1621261055
transform -1 0 44064 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_72
timestamp 1621261055
transform -1 0 44640 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_443
timestamp 1621261055
transform 1 0 43680 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_453
timestamp 1621261055
transform 1 0 44640 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_455
timestamp 1621261055
transform 1 0 44832 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_460
timestamp 1621261055
transform 1 0 45312 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1022
timestamp 1621261055
transform 1 0 46080 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output389
timestamp 1621261055
transform -1 0 46944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_22
timestamp 1621261055
transform -1 0 46560 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_469
timestamp 1621261055
transform 1 0 46176 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_477
timestamp 1621261055
transform 1 0 46944 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output391
timestamp 1621261055
transform 1 0 48000 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output429
timestamp 1621261055
transform -1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_81
timestamp 1621261055
transform -1 0 48768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_485
timestamp 1621261055
transform 1 0 47712 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_487
timestamp 1621261055
transform 1 0 47904 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_492
timestamp 1621261055
transform 1 0 48384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_500
timestamp 1621261055
transform 1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_504
timestamp 1621261055
transform 1 0 49536 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1023
timestamp 1621261055
transform 1 0 51360 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output392
timestamp 1621261055
transform 1 0 49632 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output430
timestamp 1621261055
transform -1 0 50784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_83
timestamp 1621261055
transform -1 0 50400 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_509
timestamp 1621261055
transform 1 0 50016 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_517
timestamp 1621261055
transform 1 0 50784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_521
timestamp 1621261055
transform 1 0 51168 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_524
timestamp 1621261055
transform 1 0 51456 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output393
timestamp 1621261055
transform -1 0 52224 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output394
timestamp 1621261055
transform -1 0 53184 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output432
timestamp 1621261055
transform -1 0 53952 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_24
timestamp 1621261055
transform -1 0 51840 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_25
timestamp 1621261055
transform -1 0 52416 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_26
timestamp 1621261055
transform -1 0 52800 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_85
timestamp 1621261055
transform -1 0 53568 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_534
timestamp 1621261055
transform 1 0 52416 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_542
timestamp 1621261055
transform 1 0 53184 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output395
timestamp 1621261055
transform 1 0 54336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output433
timestamp 1621261055
transform -1 0 55488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_86
timestamp 1621261055
transform -1 0 54144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_87
timestamp 1621261055
transform -1 0 55104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_552
timestamp 1621261055
transform 1 0 54144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_558
timestamp 1621261055
transform 1 0 54720 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_566
timestamp 1621261055
transform 1 0 55488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1024
timestamp 1621261055
transform 1 0 56640 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input30
timestamp 1621261055
transform 1 0 57120 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output396
timestamp 1621261055
transform 1 0 55872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_574
timestamp 1621261055
transform 1 0 56256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_579
timestamp 1621261055
transform 1 0 56736 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_587
timestamp 1621261055
transform 1 0 57504 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_161
timestamp 1621261055
transform -1 0 58848 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_595
timestamp 1621261055
transform 1 0 58272 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_162
timestamp 1621261055
transform 1 0 1152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input12
timestamp 1621261055
transform 1 0 2400 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_9
timestamp 1621261055
transform 1 0 2016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_18
timestamp 1621261055
transform 1 0 2880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1025
timestamp 1621261055
transform 1 0 3840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input32
timestamp 1621261055
transform 1 0 4896 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_26
timestamp 1621261055
transform 1 0 3648 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_29
timestamp 1621261055
transform 1 0 3936 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_37
timestamp 1621261055
transform 1 0 4704 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1026
timestamp 1621261055
transform 1 0 6528 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input23
timestamp 1621261055
transform 1 0 5760 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input33
timestamp 1621261055
transform 1 0 7008 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_44
timestamp 1621261055
transform 1 0 5376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_52
timestamp 1621261055
transform 1 0 6144 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_57
timestamp 1621261055
transform 1 0 6624 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1027
timestamp 1621261055
transform 1 0 9216 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input34
timestamp 1621261055
transform 1 0 8064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_66
timestamp 1621261055
transform 1 0 7488 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_70
timestamp 1621261055
transform 1 0 7872 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_76
timestamp 1621261055
transform 1 0 8448 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  input35
timestamp 1621261055
transform 1 0 9696 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input36
timestamp 1621261055
transform 1 0 11040 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_85
timestamp 1621261055
transform 1 0 9312 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_93
timestamp 1621261055
transform 1 0 10080 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_101
timestamp 1621261055
transform 1 0 10848 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1028
timestamp 1621261055
transform 1 0 11904 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input37
timestamp 1621261055
transform 1 0 12768 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_108
timestamp 1621261055
transform 1 0 11520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_113
timestamp 1621261055
transform 1 0 12000 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_126
timestamp 1621261055
transform 1 0 13248 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1029
timestamp 1621261055
transform 1 0 14592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input38
timestamp 1621261055
transform 1 0 15072 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output369
timestamp 1621261055
transform 1 0 13824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_1
timestamp 1621261055
transform 1 0 13632 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_136
timestamp 1621261055
transform 1 0 14208 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_141
timestamp 1621261055
transform 1 0 14688 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1030
timestamp 1621261055
transform 1 0 17280 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input2
timestamp 1621261055
transform 1 0 15936 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_149
timestamp 1621261055
transform 1 0 15456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_153
timestamp 1621261055
transform 1 0 15840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_159
timestamp 1621261055
transform 1 0 16416 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_167
timestamp 1621261055
transform 1 0 17184 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input3
timestamp 1621261055
transform 1 0 17760 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input4
timestamp 1621261055
transform 1 0 19104 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_169
timestamp 1621261055
transform 1 0 17376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_177
timestamp 1621261055
transform 1 0 18144 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_185
timestamp 1621261055
transform 1 0 18912 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1031
timestamp 1621261055
transform 1 0 19968 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input5
timestamp 1621261055
transform 1 0 20640 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_3
timestamp 1621261055
transform 1 0 21216 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_192
timestamp 1621261055
transform 1 0 19584 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_197
timestamp 1621261055
transform 1 0 20064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_201
timestamp 1621261055
transform 1 0 20448 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_207
timestamp 1621261055
transform 1 0 21024 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1032
timestamp 1621261055
transform 1 0 22656 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input6
timestamp 1621261055
transform 1 0 23136 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_2  output370
timestamp 1621261055
transform 1 0 21408 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_215
timestamp 1621261055
transform 1 0 21792 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_223
timestamp 1621261055
transform 1 0 22560 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_225
timestamp 1621261055
transform 1 0 22752 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1033
timestamp 1621261055
transform 1 0 25344 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input7
timestamp 1621261055
transform 1 0 24000 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_234
timestamp 1621261055
transform 1 0 23616 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_242
timestamp 1621261055
transform 1 0 24384 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_250
timestamp 1621261055
transform 1 0 25152 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__buf_2  input8
timestamp 1621261055
transform 1 0 25824 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input9
timestamp 1621261055
transform 1 0 26976 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_253
timestamp 1621261055
transform 1 0 25440 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_262
timestamp 1621261055
transform 1 0 26304 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_266
timestamp 1621261055
transform 1 0 26688 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_268
timestamp 1621261055
transform 1 0 26880 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_273
timestamp 1621261055
transform 1 0 27360 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1034
timestamp 1621261055
transform 1 0 28032 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input10
timestamp 1621261055
transform 1 0 28608 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_277
timestamp 1621261055
transform 1 0 27744 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_279
timestamp 1621261055
transform 1 0 27936 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_281
timestamp 1621261055
transform 1 0 28128 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_285
timestamp 1621261055
transform 1 0 28512 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_291
timestamp 1621261055
transform 1 0 29088 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1035
timestamp 1621261055
transform 1 0 30720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input11
timestamp 1621261055
transform 1 0 29952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_299
timestamp 1621261055
transform 1 0 29856 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_304
timestamp 1621261055
transform 1 0 30336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_309
timestamp 1621261055
transform 1 0 30816 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1036
timestamp 1621261055
transform 1 0 33408 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input13
timestamp 1621261055
transform 1 0 31680 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_2  output377
timestamp 1621261055
transform 1 0 32544 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_317
timestamp 1621261055
transform 1 0 31584 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_323
timestamp 1621261055
transform 1 0 32160 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_331
timestamp 1621261055
transform 1 0 32928 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_335
timestamp 1621261055
transform 1 0 33312 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input14
timestamp 1621261055
transform 1 0 33888 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input15
timestamp 1621261055
transform 1 0 34848 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_337
timestamp 1621261055
transform 1 0 33504 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_346
timestamp 1621261055
transform 1 0 34368 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_350
timestamp 1621261055
transform 1 0 34752 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_356
timestamp 1621261055
transform 1 0 35328 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1037
timestamp 1621261055
transform 1 0 36096 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input16
timestamp 1621261055
transform 1 0 36576 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_365
timestamp 1621261055
transform 1 0 36192 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_373
timestamp 1621261055
transform 1 0 36960 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1038
timestamp 1621261055
transform 1 0 38784 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input17 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 37824 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__fill_1  FILLER_81_381
timestamp 1621261055
transform 1 0 37728 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_388
timestamp 1621261055
transform 1 0 38400 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_393
timestamp 1621261055
transform 1 0 38880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1039
timestamp 1621261055
transform 1 0 41472 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input18
timestamp 1621261055
transform 1 0 39648 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_2  output383
timestamp 1621261055
transform -1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_13
timestamp 1621261055
transform -1 0 40608 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_14
timestamp 1621261055
transform -1 0 41184 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_407
timestamp 1621261055
transform 1 0 40224 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_417
timestamp 1621261055
transform 1 0 41184 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_419
timestamp 1621261055
transform 1 0 41376 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input19
timestamp 1621261055
transform 1 0 41952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_4  input20
timestamp 1621261055
transform 1 0 42816 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_421
timestamp 1621261055
transform 1 0 41568 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_429
timestamp 1621261055
transform 1 0 42336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_433
timestamp 1621261055
transform 1 0 42720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_440
timestamp 1621261055
transform 1 0 43392 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1040
timestamp 1621261055
transform 1 0 44160 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input21
timestamp 1621261055
transform 1 0 44640 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_449
timestamp 1621261055
transform 1 0 44256 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_459
timestamp 1621261055
transform 1 0 45216 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1041
timestamp 1621261055
transform 1 0 46848 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input22
timestamp 1621261055
transform 1 0 45888 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input24
timestamp 1621261055
transform 1 0 47520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_463
timestamp 1621261055
transform 1 0 45600 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_465
timestamp 1621261055
transform 1 0 45792 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_472
timestamp 1621261055
transform 1 0 46464 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_477
timestamp 1621261055
transform 1 0 46944 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_481
timestamp 1621261055
transform 1 0 47328 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1042
timestamp 1621261055
transform 1 0 49536 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input25
timestamp 1621261055
transform 1 0 48576 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_487
timestamp 1621261055
transform 1 0 47904 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_491
timestamp 1621261055
transform 1 0 48288 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_493
timestamp 1621261055
transform 1 0 48480 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_500
timestamp 1621261055
transform 1 0 49152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_4  input26
timestamp 1621261055
transform 1 0 50688 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_8  FILLER_81_505
timestamp 1621261055
transform 1 0 49632 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_513
timestamp 1621261055
transform 1 0 50400 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_515
timestamp 1621261055
transform 1 0 50592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_522
timestamp 1621261055
transform 1 0 51264 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1043
timestamp 1621261055
transform 1 0 52224 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input27
timestamp 1621261055
transform 1 0 52704 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_530
timestamp 1621261055
transform 1 0 52032 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_533
timestamp 1621261055
transform 1 0 52320 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_541
timestamp 1621261055
transform 1 0 53088 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1044
timestamp 1621261055
transform 1 0 54912 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input28
timestamp 1621261055
transform 1 0 53856 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_4  input29
timestamp 1621261055
transform 1 0 55392 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_555
timestamp 1621261055
transform 1 0 54432 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_559
timestamp 1621261055
transform 1 0 54816 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_561
timestamp 1621261055
transform 1 0 55008 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1045
timestamp 1621261055
transform 1 0 57600 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input31
timestamp 1621261055
transform 1 0 56640 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_571
timestamp 1621261055
transform 1 0 55968 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_575
timestamp 1621261055
transform 1 0 56352 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_577
timestamp 1621261055
transform 1 0 56544 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_584
timestamp 1621261055
transform 1 0 57216 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_163
timestamp 1621261055
transform -1 0 58848 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_589
timestamp 1621261055
transform 1 0 57696 0 1 56610
box -38 -49 806 715
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 12980 0 13036 800 6 la_data_in[0]
port 114 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_data_in[100]
port 115 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_data_in[101]
port 116 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[102]
port 117 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[103]
port 118 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[104]
port 119 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_data_in[105]
port 120 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_data_in[106]
port 121 nsew signal input
rlabel metal2 s 52244 0 52300 800 6 la_data_in[107]
port 122 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[108]
port 123 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[109]
port 124 nsew signal input
rlabel metal2 s 16628 0 16684 800 6 la_data_in[10]
port 125 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[110]
port 126 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_data_in[111]
port 127 nsew signal input
rlabel metal2 s 54068 0 54124 800 6 la_data_in[112]
port 128 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[113]
port 129 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[114]
port 130 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[115]
port 131 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[116]
port 132 nsew signal input
rlabel metal2 s 55892 0 55948 800 6 la_data_in[117]
port 133 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[118]
port 134 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[119]
port 135 nsew signal input
rlabel metal2 s 17012 0 17068 800 6 la_data_in[11]
port 136 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[120]
port 137 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[121]
port 138 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[122]
port 139 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[123]
port 140 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[124]
port 141 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[125]
port 142 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[126]
port 143 nsew signal input
rlabel metal2 s 59636 0 59692 800 6 la_data_in[127]
port 144 nsew signal input
rlabel metal2 s 17396 0 17452 800 6 la_data_in[12]
port 145 nsew signal input
rlabel metal2 s 17684 0 17740 800 6 la_data_in[13]
port 146 nsew signal input
rlabel metal2 s 18068 0 18124 800 6 la_data_in[14]
port 147 nsew signal input
rlabel metal2 s 18452 0 18508 800 6 la_data_in[15]
port 148 nsew signal input
rlabel metal2 s 18836 0 18892 800 6 la_data_in[16]
port 149 nsew signal input
rlabel metal2 s 19220 0 19276 800 6 la_data_in[17]
port 150 nsew signal input
rlabel metal2 s 19604 0 19660 800 6 la_data_in[18]
port 151 nsew signal input
rlabel metal2 s 19892 0 19948 800 6 la_data_in[19]
port 152 nsew signal input
rlabel metal2 s 13364 0 13420 800 6 la_data_in[1]
port 153 nsew signal input
rlabel metal2 s 20276 0 20332 800 6 la_data_in[20]
port 154 nsew signal input
rlabel metal2 s 20660 0 20716 800 6 la_data_in[21]
port 155 nsew signal input
rlabel metal2 s 21044 0 21100 800 6 la_data_in[22]
port 156 nsew signal input
rlabel metal2 s 21428 0 21484 800 6 la_data_in[23]
port 157 nsew signal input
rlabel metal2 s 21812 0 21868 800 6 la_data_in[24]
port 158 nsew signal input
rlabel metal2 s 22100 0 22156 800 6 la_data_in[25]
port 159 nsew signal input
rlabel metal2 s 22484 0 22540 800 6 la_data_in[26]
port 160 nsew signal input
rlabel metal2 s 22868 0 22924 800 6 la_data_in[27]
port 161 nsew signal input
rlabel metal2 s 23252 0 23308 800 6 la_data_in[28]
port 162 nsew signal input
rlabel metal2 s 23636 0 23692 800 6 la_data_in[29]
port 163 nsew signal input
rlabel metal2 s 13652 0 13708 800 6 la_data_in[2]
port 164 nsew signal input
rlabel metal2 s 24020 0 24076 800 6 la_data_in[30]
port 165 nsew signal input
rlabel metal2 s 24308 0 24364 800 6 la_data_in[31]
port 166 nsew signal input
rlabel metal2 s 24692 0 24748 800 6 la_data_in[32]
port 167 nsew signal input
rlabel metal2 s 25076 0 25132 800 6 la_data_in[33]
port 168 nsew signal input
rlabel metal2 s 25460 0 25516 800 6 la_data_in[34]
port 169 nsew signal input
rlabel metal2 s 25844 0 25900 800 6 la_data_in[35]
port 170 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_in[36]
port 171 nsew signal input
rlabel metal2 s 26516 0 26572 800 6 la_data_in[37]
port 172 nsew signal input
rlabel metal2 s 26900 0 26956 800 6 la_data_in[38]
port 173 nsew signal input
rlabel metal2 s 27284 0 27340 800 6 la_data_in[39]
port 174 nsew signal input
rlabel metal2 s 14036 0 14092 800 6 la_data_in[3]
port 175 nsew signal input
rlabel metal2 s 27668 0 27724 800 6 la_data_in[40]
port 176 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_data_in[41]
port 177 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 la_data_in[42]
port 178 nsew signal input
rlabel metal2 s 28724 0 28780 800 6 la_data_in[43]
port 179 nsew signal input
rlabel metal2 s 29108 0 29164 800 6 la_data_in[44]
port 180 nsew signal input
rlabel metal2 s 29492 0 29548 800 6 la_data_in[45]
port 181 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_data_in[46]
port 182 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_data_in[47]
port 183 nsew signal input
rlabel metal2 s 30548 0 30604 800 6 la_data_in[48]
port 184 nsew signal input
rlabel metal2 s 30932 0 30988 800 6 la_data_in[49]
port 185 nsew signal input
rlabel metal2 s 14420 0 14476 800 6 la_data_in[4]
port 186 nsew signal input
rlabel metal2 s 31316 0 31372 800 6 la_data_in[50]
port 187 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_data_in[51]
port 188 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_data_in[52]
port 189 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_data_in[53]
port 190 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 la_data_in[54]
port 191 nsew signal input
rlabel metal2 s 33140 0 33196 800 6 la_data_in[55]
port 192 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_data_in[56]
port 193 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_data_in[57]
port 194 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_data_in[58]
port 195 nsew signal input
rlabel metal2 s 34580 0 34636 800 6 la_data_in[59]
port 196 nsew signal input
rlabel metal2 s 14804 0 14860 800 6 la_data_in[5]
port 197 nsew signal input
rlabel metal2 s 34964 0 35020 800 6 la_data_in[60]
port 198 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_data_in[61]
port 199 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_data_in[62]
port 200 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_data_in[63]
port 201 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_data_in[64]
port 202 nsew signal input
rlabel metal2 s 36788 0 36844 800 6 la_data_in[65]
port 203 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_data_in[66]
port 204 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_data_in[67]
port 205 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_data_in[68]
port 206 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_data_in[69]
port 207 nsew signal input
rlabel metal2 s 15188 0 15244 800 6 la_data_in[6]
port 208 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_data_in[70]
port 209 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_data_in[71]
port 210 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_data_in[72]
port 211 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_data_in[73]
port 212 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_data_in[74]
port 213 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_data_in[75]
port 214 nsew signal input
rlabel metal2 s 40916 0 40972 800 6 la_data_in[76]
port 215 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_data_in[77]
port 216 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_data_in[78]
port 217 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_data_in[79]
port 218 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 219 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_data_in[80]
port 220 nsew signal input
rlabel metal2 s 42740 0 42796 800 6 la_data_in[81]
port 221 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_data_in[82]
port 222 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_data_in[83]
port 223 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_data_in[84]
port 224 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_data_in[85]
port 225 nsew signal input
rlabel metal2 s 44564 0 44620 800 6 la_data_in[86]
port 226 nsew signal input
rlabel metal2 s 44948 0 45004 800 6 la_data_in[87]
port 227 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_data_in[88]
port 228 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_data_in[89]
port 229 nsew signal input
rlabel metal2 s 15860 0 15916 800 6 la_data_in[8]
port 230 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_data_in[90]
port 231 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_data_in[91]
port 232 nsew signal input
rlabel metal2 s 46772 0 46828 800 6 la_data_in[92]
port 233 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[93]
port 234 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_data_in[94]
port 235 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_data_in[95]
port 236 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_data_in[96]
port 237 nsew signal input
rlabel metal2 s 48596 0 48652 800 6 la_data_in[97]
port 238 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[98]
port 239 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[99]
port 240 nsew signal input
rlabel metal2 s 16244 0 16300 800 6 la_data_in[9]
port 241 nsew signal input
rlabel metal2 s 13076 0 13132 800 6 la_data_out[0]
port 242 nsew signal tristate
rlabel metal2 s 49844 0 49900 800 6 la_data_out[100]
port 243 nsew signal tristate
rlabel metal2 s 50132 0 50188 800 6 la_data_out[101]
port 244 nsew signal tristate
rlabel metal2 s 50516 0 50572 800 6 la_data_out[102]
port 245 nsew signal tristate
rlabel metal2 s 50900 0 50956 800 6 la_data_out[103]
port 246 nsew signal tristate
rlabel metal2 s 51284 0 51340 800 6 la_data_out[104]
port 247 nsew signal tristate
rlabel metal2 s 51668 0 51724 800 6 la_data_out[105]
port 248 nsew signal tristate
rlabel metal2 s 52052 0 52108 800 6 la_data_out[106]
port 249 nsew signal tristate
rlabel metal2 s 52340 0 52396 800 6 la_data_out[107]
port 250 nsew signal tristate
rlabel metal2 s 52724 0 52780 800 6 la_data_out[108]
port 251 nsew signal tristate
rlabel metal2 s 53108 0 53164 800 6 la_data_out[109]
port 252 nsew signal tristate
rlabel metal2 s 16724 0 16780 800 6 la_data_out[10]
port 253 nsew signal tristate
rlabel metal2 s 53492 0 53548 800 6 la_data_out[110]
port 254 nsew signal tristate
rlabel metal2 s 53876 0 53932 800 6 la_data_out[111]
port 255 nsew signal tristate
rlabel metal2 s 54260 0 54316 800 6 la_data_out[112]
port 256 nsew signal tristate
rlabel metal2 s 54548 0 54604 800 6 la_data_out[113]
port 257 nsew signal tristate
rlabel metal2 s 54932 0 54988 800 6 la_data_out[114]
port 258 nsew signal tristate
rlabel metal2 s 55316 0 55372 800 6 la_data_out[115]
port 259 nsew signal tristate
rlabel metal2 s 55700 0 55756 800 6 la_data_out[116]
port 260 nsew signal tristate
rlabel metal2 s 56084 0 56140 800 6 la_data_out[117]
port 261 nsew signal tristate
rlabel metal2 s 56468 0 56524 800 6 la_data_out[118]
port 262 nsew signal tristate
rlabel metal2 s 56756 0 56812 800 6 la_data_out[119]
port 263 nsew signal tristate
rlabel metal2 s 17108 0 17164 800 6 la_data_out[11]
port 264 nsew signal tristate
rlabel metal2 s 57140 0 57196 800 6 la_data_out[120]
port 265 nsew signal tristate
rlabel metal2 s 57524 0 57580 800 6 la_data_out[121]
port 266 nsew signal tristate
rlabel metal2 s 57908 0 57964 800 6 la_data_out[122]
port 267 nsew signal tristate
rlabel metal2 s 58292 0 58348 800 6 la_data_out[123]
port 268 nsew signal tristate
rlabel metal2 s 58580 0 58636 800 6 la_data_out[124]
port 269 nsew signal tristate
rlabel metal2 s 58964 0 59020 800 6 la_data_out[125]
port 270 nsew signal tristate
rlabel metal2 s 59348 0 59404 800 6 la_data_out[126]
port 271 nsew signal tristate
rlabel metal2 s 59732 0 59788 800 6 la_data_out[127]
port 272 nsew signal tristate
rlabel metal2 s 17492 0 17548 800 6 la_data_out[12]
port 273 nsew signal tristate
rlabel metal2 s 17876 0 17932 800 6 la_data_out[13]
port 274 nsew signal tristate
rlabel metal2 s 18260 0 18316 800 6 la_data_out[14]
port 275 nsew signal tristate
rlabel metal2 s 18548 0 18604 800 6 la_data_out[15]
port 276 nsew signal tristate
rlabel metal2 s 18932 0 18988 800 6 la_data_out[16]
port 277 nsew signal tristate
rlabel metal2 s 19316 0 19372 800 6 la_data_out[17]
port 278 nsew signal tristate
rlabel metal2 s 19700 0 19756 800 6 la_data_out[18]
port 279 nsew signal tristate
rlabel metal2 s 20084 0 20140 800 6 la_data_out[19]
port 280 nsew signal tristate
rlabel metal2 s 13460 0 13516 800 6 la_data_out[1]
port 281 nsew signal tristate
rlabel metal2 s 20468 0 20524 800 6 la_data_out[20]
port 282 nsew signal tristate
rlabel metal2 s 20756 0 20812 800 6 la_data_out[21]
port 283 nsew signal tristate
rlabel metal2 s 21140 0 21196 800 6 la_data_out[22]
port 284 nsew signal tristate
rlabel metal2 s 21524 0 21580 800 6 la_data_out[23]
port 285 nsew signal tristate
rlabel metal2 s 21908 0 21964 800 6 la_data_out[24]
port 286 nsew signal tristate
rlabel metal2 s 22292 0 22348 800 6 la_data_out[25]
port 287 nsew signal tristate
rlabel metal2 s 22580 0 22636 800 6 la_data_out[26]
port 288 nsew signal tristate
rlabel metal2 s 22964 0 23020 800 6 la_data_out[27]
port 289 nsew signal tristate
rlabel metal2 s 23348 0 23404 800 6 la_data_out[28]
port 290 nsew signal tristate
rlabel metal2 s 23732 0 23788 800 6 la_data_out[29]
port 291 nsew signal tristate
rlabel metal2 s 13844 0 13900 800 6 la_data_out[2]
port 292 nsew signal tristate
rlabel metal2 s 24116 0 24172 800 6 la_data_out[30]
port 293 nsew signal tristate
rlabel metal2 s 24500 0 24556 800 6 la_data_out[31]
port 294 nsew signal tristate
rlabel metal2 s 24788 0 24844 800 6 la_data_out[32]
port 295 nsew signal tristate
rlabel metal2 s 25172 0 25228 800 6 la_data_out[33]
port 296 nsew signal tristate
rlabel metal2 s 25556 0 25612 800 6 la_data_out[34]
port 297 nsew signal tristate
rlabel metal2 s 25940 0 25996 800 6 la_data_out[35]
port 298 nsew signal tristate
rlabel metal2 s 26324 0 26380 800 6 la_data_out[36]
port 299 nsew signal tristate
rlabel metal2 s 26708 0 26764 800 6 la_data_out[37]
port 300 nsew signal tristate
rlabel metal2 s 26996 0 27052 800 6 la_data_out[38]
port 301 nsew signal tristate
rlabel metal2 s 27380 0 27436 800 6 la_data_out[39]
port 302 nsew signal tristate
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 303 nsew signal tristate
rlabel metal2 s 27764 0 27820 800 6 la_data_out[40]
port 304 nsew signal tristate
rlabel metal2 s 28148 0 28204 800 6 la_data_out[41]
port 305 nsew signal tristate
rlabel metal2 s 28532 0 28588 800 6 la_data_out[42]
port 306 nsew signal tristate
rlabel metal2 s 28916 0 28972 800 6 la_data_out[43]
port 307 nsew signal tristate
rlabel metal2 s 29204 0 29260 800 6 la_data_out[44]
port 308 nsew signal tristate
rlabel metal2 s 29588 0 29644 800 6 la_data_out[45]
port 309 nsew signal tristate
rlabel metal2 s 29972 0 30028 800 6 la_data_out[46]
port 310 nsew signal tristate
rlabel metal2 s 30356 0 30412 800 6 la_data_out[47]
port 311 nsew signal tristate
rlabel metal2 s 30740 0 30796 800 6 la_data_out[48]
port 312 nsew signal tristate
rlabel metal2 s 31028 0 31084 800 6 la_data_out[49]
port 313 nsew signal tristate
rlabel metal2 s 14516 0 14572 800 6 la_data_out[4]
port 314 nsew signal tristate
rlabel metal2 s 31412 0 31468 800 6 la_data_out[50]
port 315 nsew signal tristate
rlabel metal2 s 31796 0 31852 800 6 la_data_out[51]
port 316 nsew signal tristate
rlabel metal2 s 32180 0 32236 800 6 la_data_out[52]
port 317 nsew signal tristate
rlabel metal2 s 32564 0 32620 800 6 la_data_out[53]
port 318 nsew signal tristate
rlabel metal2 s 32948 0 33004 800 6 la_data_out[54]
port 319 nsew signal tristate
rlabel metal2 s 33236 0 33292 800 6 la_data_out[55]
port 320 nsew signal tristate
rlabel metal2 s 33620 0 33676 800 6 la_data_out[56]
port 321 nsew signal tristate
rlabel metal2 s 34004 0 34060 800 6 la_data_out[57]
port 322 nsew signal tristate
rlabel metal2 s 34388 0 34444 800 6 la_data_out[58]
port 323 nsew signal tristate
rlabel metal2 s 34772 0 34828 800 6 la_data_out[59]
port 324 nsew signal tristate
rlabel metal2 s 14900 0 14956 800 6 la_data_out[5]
port 325 nsew signal tristate
rlabel metal2 s 35156 0 35212 800 6 la_data_out[60]
port 326 nsew signal tristate
rlabel metal2 s 35444 0 35500 800 6 la_data_out[61]
port 327 nsew signal tristate
rlabel metal2 s 35828 0 35884 800 6 la_data_out[62]
port 328 nsew signal tristate
rlabel metal2 s 36212 0 36268 800 6 la_data_out[63]
port 329 nsew signal tristate
rlabel metal2 s 36596 0 36652 800 6 la_data_out[64]
port 330 nsew signal tristate
rlabel metal2 s 36980 0 37036 800 6 la_data_out[65]
port 331 nsew signal tristate
rlabel metal2 s 37364 0 37420 800 6 la_data_out[66]
port 332 nsew signal tristate
rlabel metal2 s 37652 0 37708 800 6 la_data_out[67]
port 333 nsew signal tristate
rlabel metal2 s 38036 0 38092 800 6 la_data_out[68]
port 334 nsew signal tristate
rlabel metal2 s 38420 0 38476 800 6 la_data_out[69]
port 335 nsew signal tristate
rlabel metal2 s 15284 0 15340 800 6 la_data_out[6]
port 336 nsew signal tristate
rlabel metal2 s 38804 0 38860 800 6 la_data_out[70]
port 337 nsew signal tristate
rlabel metal2 s 39188 0 39244 800 6 la_data_out[71]
port 338 nsew signal tristate
rlabel metal2 s 39476 0 39532 800 6 la_data_out[72]
port 339 nsew signal tristate
rlabel metal2 s 39860 0 39916 800 6 la_data_out[73]
port 340 nsew signal tristate
rlabel metal2 s 40244 0 40300 800 6 la_data_out[74]
port 341 nsew signal tristate
rlabel metal2 s 40628 0 40684 800 6 la_data_out[75]
port 342 nsew signal tristate
rlabel metal2 s 41012 0 41068 800 6 la_data_out[76]
port 343 nsew signal tristate
rlabel metal2 s 41396 0 41452 800 6 la_data_out[77]
port 344 nsew signal tristate
rlabel metal2 s 41684 0 41740 800 6 la_data_out[78]
port 345 nsew signal tristate
rlabel metal2 s 42068 0 42124 800 6 la_data_out[79]
port 346 nsew signal tristate
rlabel metal2 s 15668 0 15724 800 6 la_data_out[7]
port 347 nsew signal tristate
rlabel metal2 s 42452 0 42508 800 6 la_data_out[80]
port 348 nsew signal tristate
rlabel metal2 s 42836 0 42892 800 6 la_data_out[81]
port 349 nsew signal tristate
rlabel metal2 s 43220 0 43276 800 6 la_data_out[82]
port 350 nsew signal tristate
rlabel metal2 s 43604 0 43660 800 6 la_data_out[83]
port 351 nsew signal tristate
rlabel metal2 s 43892 0 43948 800 6 la_data_out[84]
port 352 nsew signal tristate
rlabel metal2 s 44276 0 44332 800 6 la_data_out[85]
port 353 nsew signal tristate
rlabel metal2 s 44660 0 44716 800 6 la_data_out[86]
port 354 nsew signal tristate
rlabel metal2 s 45044 0 45100 800 6 la_data_out[87]
port 355 nsew signal tristate
rlabel metal2 s 45428 0 45484 800 6 la_data_out[88]
port 356 nsew signal tristate
rlabel metal2 s 45812 0 45868 800 6 la_data_out[89]
port 357 nsew signal tristate
rlabel metal2 s 16052 0 16108 800 6 la_data_out[8]
port 358 nsew signal tristate
rlabel metal2 s 46100 0 46156 800 6 la_data_out[90]
port 359 nsew signal tristate
rlabel metal2 s 46484 0 46540 800 6 la_data_out[91]
port 360 nsew signal tristate
rlabel metal2 s 46868 0 46924 800 6 la_data_out[92]
port 361 nsew signal tristate
rlabel metal2 s 47252 0 47308 800 6 la_data_out[93]
port 362 nsew signal tristate
rlabel metal2 s 47636 0 47692 800 6 la_data_out[94]
port 363 nsew signal tristate
rlabel metal2 s 48020 0 48076 800 6 la_data_out[95]
port 364 nsew signal tristate
rlabel metal2 s 48308 0 48364 800 6 la_data_out[96]
port 365 nsew signal tristate
rlabel metal2 s 48692 0 48748 800 6 la_data_out[97]
port 366 nsew signal tristate
rlabel metal2 s 49076 0 49132 800 6 la_data_out[98]
port 367 nsew signal tristate
rlabel metal2 s 49460 0 49516 800 6 la_data_out[99]
port 368 nsew signal tristate
rlabel metal2 s 16340 0 16396 800 6 la_data_out[9]
port 369 nsew signal tristate
rlabel metal2 s 13172 0 13228 800 6 la_oen[0]
port 370 nsew signal input
rlabel metal2 s 49940 0 49996 800 6 la_oen[100]
port 371 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oen[101]
port 372 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oen[102]
port 373 nsew signal input
rlabel metal2 s 50996 0 51052 800 6 la_oen[103]
port 374 nsew signal input
rlabel metal2 s 51380 0 51436 800 6 la_oen[104]
port 375 nsew signal input
rlabel metal2 s 51764 0 51820 800 6 la_oen[105]
port 376 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oen[106]
port 377 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oen[107]
port 378 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oen[108]
port 379 nsew signal input
rlabel metal2 s 53204 0 53260 800 6 la_oen[109]
port 380 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_oen[10]
port 381 nsew signal input
rlabel metal2 s 53588 0 53644 800 6 la_oen[110]
port 382 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oen[111]
port 383 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oen[112]
port 384 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oen[113]
port 385 nsew signal input
rlabel metal2 s 55028 0 55084 800 6 la_oen[114]
port 386 nsew signal input
rlabel metal2 s 55412 0 55468 800 6 la_oen[115]
port 387 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oen[116]
port 388 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oen[117]
port 389 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oen[118]
port 390 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oen[119]
port 391 nsew signal input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 392 nsew signal input
rlabel metal2 s 57236 0 57292 800 6 la_oen[120]
port 393 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oen[121]
port 394 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oen[122]
port 395 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oen[123]
port 396 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oen[124]
port 397 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oen[125]
port 398 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oen[126]
port 399 nsew signal input
rlabel metal2 s 59828 0 59884 800 6 la_oen[127]
port 400 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_oen[12]
port 401 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_oen[13]
port 402 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_oen[14]
port 403 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_oen[15]
port 404 nsew signal input
rlabel metal2 s 19028 0 19084 800 6 la_oen[16]
port 405 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 406 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_oen[18]
port 407 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_oen[19]
port 408 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_oen[1]
port 409 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_oen[20]
port 410 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_oen[21]
port 411 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_oen[22]
port 412 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 413 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_oen[24]
port 414 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_oen[25]
port 415 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_oen[26]
port 416 nsew signal input
rlabel metal2 s 23156 0 23212 800 6 la_oen[27]
port 417 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_oen[28]
port 418 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 419 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_oen[2]
port 420 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_oen[30]
port 421 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_oen[31]
port 422 nsew signal input
rlabel metal2 s 24980 0 25036 800 6 la_oen[32]
port 423 nsew signal input
rlabel metal2 s 25364 0 25420 800 6 la_oen[33]
port 424 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_oen[34]
port 425 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 426 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_oen[36]
port 427 nsew signal input
rlabel metal2 s 26804 0 26860 800 6 la_oen[37]
port 428 nsew signal input
rlabel metal2 s 27188 0 27244 800 6 la_oen[38]
port 429 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_oen[39]
port 430 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_oen[3]
port 431 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_oen[40]
port 432 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 433 nsew signal input
rlabel metal2 s 28628 0 28684 800 6 la_oen[42]
port 434 nsew signal input
rlabel metal2 s 29012 0 29068 800 6 la_oen[43]
port 435 nsew signal input
rlabel metal2 s 29396 0 29452 800 6 la_oen[44]
port 436 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_oen[45]
port 437 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_oen[46]
port 438 nsew signal input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 439 nsew signal input
rlabel metal2 s 30836 0 30892 800 6 la_oen[48]
port 440 nsew signal input
rlabel metal2 s 31220 0 31276 800 6 la_oen[49]
port 441 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_oen[4]
port 442 nsew signal input
rlabel metal2 s 31604 0 31660 800 6 la_oen[50]
port 443 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_oen[51]
port 444 nsew signal input
rlabel metal2 s 32276 0 32332 800 6 la_oen[52]
port 445 nsew signal input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 446 nsew signal input
rlabel metal2 s 33044 0 33100 800 6 la_oen[54]
port 447 nsew signal input
rlabel metal2 s 33428 0 33484 800 6 la_oen[55]
port 448 nsew signal input
rlabel metal2 s 33812 0 33868 800 6 la_oen[56]
port 449 nsew signal input
rlabel metal2 s 34100 0 34156 800 6 la_oen[57]
port 450 nsew signal input
rlabel metal2 s 34484 0 34540 800 6 la_oen[58]
port 451 nsew signal input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 452 nsew signal input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 453 nsew signal input
rlabel metal2 s 35252 0 35308 800 6 la_oen[60]
port 454 nsew signal input
rlabel metal2 s 35636 0 35692 800 6 la_oen[61]
port 455 nsew signal input
rlabel metal2 s 36020 0 36076 800 6 la_oen[62]
port 456 nsew signal input
rlabel metal2 s 36308 0 36364 800 6 la_oen[63]
port 457 nsew signal input
rlabel metal2 s 36692 0 36748 800 6 la_oen[64]
port 458 nsew signal input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 459 nsew signal input
rlabel metal2 s 37460 0 37516 800 6 la_oen[66]
port 460 nsew signal input
rlabel metal2 s 37844 0 37900 800 6 la_oen[67]
port 461 nsew signal input
rlabel metal2 s 38132 0 38188 800 6 la_oen[68]
port 462 nsew signal input
rlabel metal2 s 38516 0 38572 800 6 la_oen[69]
port 463 nsew signal input
rlabel metal2 s 15380 0 15436 800 6 la_oen[6]
port 464 nsew signal input
rlabel metal2 s 38900 0 38956 800 6 la_oen[70]
port 465 nsew signal input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 466 nsew signal input
rlabel metal2 s 39668 0 39724 800 6 la_oen[72]
port 467 nsew signal input
rlabel metal2 s 40052 0 40108 800 6 la_oen[73]
port 468 nsew signal input
rlabel metal2 s 40340 0 40396 800 6 la_oen[74]
port 469 nsew signal input
rlabel metal2 s 40724 0 40780 800 6 la_oen[75]
port 470 nsew signal input
rlabel metal2 s 41108 0 41164 800 6 la_oen[76]
port 471 nsew signal input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 472 nsew signal input
rlabel metal2 s 41876 0 41932 800 6 la_oen[78]
port 473 nsew signal input
rlabel metal2 s 42260 0 42316 800 6 la_oen[79]
port 474 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_oen[7]
port 475 nsew signal input
rlabel metal2 s 42548 0 42604 800 6 la_oen[80]
port 476 nsew signal input
rlabel metal2 s 42932 0 42988 800 6 la_oen[81]
port 477 nsew signal input
rlabel metal2 s 43316 0 43372 800 6 la_oen[82]
port 478 nsew signal input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 479 nsew signal input
rlabel metal2 s 44084 0 44140 800 6 la_oen[84]
port 480 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oen[85]
port 481 nsew signal input
rlabel metal2 s 44756 0 44812 800 6 la_oen[86]
port 482 nsew signal input
rlabel metal2 s 45140 0 45196 800 6 la_oen[87]
port 483 nsew signal input
rlabel metal2 s 45524 0 45580 800 6 la_oen[88]
port 484 nsew signal input
rlabel metal2 s 45908 0 45964 800 6 la_oen[89]
port 485 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_oen[8]
port 486 nsew signal input
rlabel metal2 s 46292 0 46348 800 6 la_oen[90]
port 487 nsew signal input
rlabel metal2 s 46580 0 46636 800 6 la_oen[91]
port 488 nsew signal input
rlabel metal2 s 46964 0 47020 800 6 la_oen[92]
port 489 nsew signal input
rlabel metal2 s 47348 0 47404 800 6 la_oen[93]
port 490 nsew signal input
rlabel metal2 s 47732 0 47788 800 6 la_oen[94]
port 491 nsew signal input
rlabel metal2 s 48116 0 48172 800 6 la_oen[95]
port 492 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oen[96]
port 493 nsew signal input
rlabel metal2 s 48788 0 48844 800 6 la_oen[97]
port 494 nsew signal input
rlabel metal2 s 49172 0 49228 800 6 la_oen[98]
port 495 nsew signal input
rlabel metal2 s 49556 0 49612 800 6 la_oen[99]
port 496 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_oen[9]
port 497 nsew signal input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 498 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 499 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 500 nsew signal tristate
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 501 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_adr_i[10]
port 502 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 503 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 504 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 505 nsew signal input
rlabel metal2 s 6356 0 6412 800 6 wbs_adr_i[14]
port 506 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_adr_i[15]
port 507 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 508 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 509 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 510 nsew signal input
rlabel metal2 s 8180 0 8236 800 6 wbs_adr_i[19]
port 511 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 512 nsew signal input
rlabel metal2 s 8564 0 8620 800 6 wbs_adr_i[20]
port 513 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_adr_i[21]
port 514 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 515 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 516 nsew signal input
rlabel metal2 s 10004 0 10060 800 6 wbs_adr_i[24]
port 517 nsew signal input
rlabel metal2 s 10388 0 10444 800 6 wbs_adr_i[25]
port 518 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_adr_i[26]
port 519 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_adr_i[27]
port 520 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 521 nsew signal input
rlabel metal2 s 11828 0 11884 800 6 wbs_adr_i[29]
port 522 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 523 nsew signal input
rlabel metal2 s 12212 0 12268 800 6 wbs_adr_i[30]
port 524 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_adr_i[31]
port 525 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 526 nsew signal input
rlabel metal2 s 2708 0 2764 800 6 wbs_adr_i[4]
port 527 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 528 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 529 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 530 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 531 nsew signal input
rlabel metal2 s 4532 0 4588 800 6 wbs_adr_i[9]
port 532 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 533 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 534 nsew signal input
rlabel metal2 s 5012 0 5068 800 6 wbs_dat_i[10]
port 535 nsew signal input
rlabel metal2 s 5396 0 5452 800 6 wbs_dat_i[11]
port 536 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 537 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 538 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 539 nsew signal input
rlabel metal2 s 6836 0 6892 800 6 wbs_dat_i[15]
port 540 nsew signal input
rlabel metal2 s 7220 0 7276 800 6 wbs_dat_i[16]
port 541 nsew signal input
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_i[17]
port 542 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 543 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 544 nsew signal input
rlabel metal2 s 1364 0 1420 800 6 wbs_dat_i[1]
port 545 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 546 nsew signal input
rlabel metal2 s 9044 0 9100 800 6 wbs_dat_i[21]
port 547 nsew signal input
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_i[22]
port 548 nsew signal input
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_i[23]
port 549 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 550 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 551 nsew signal input
rlabel metal2 s 10868 0 10924 800 6 wbs_dat_i[26]
port 552 nsew signal input
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_i[27]
port 553 nsew signal input
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_i[28]
port 554 nsew signal input
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_i[29]
port 555 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 556 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 557 nsew signal input
rlabel metal2 s 12692 0 12748 800 6 wbs_dat_i[31]
port 558 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 559 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 560 nsew signal input
rlabel metal2 s 3188 0 3244 800 6 wbs_dat_i[5]
port 561 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 562 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 563 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 564 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 565 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 566 nsew signal tristate
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 567 nsew signal tristate
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 568 nsew signal tristate
rlabel metal2 s 5876 0 5932 800 6 wbs_dat_o[12]
port 569 nsew signal tristate
rlabel metal2 s 6260 0 6316 800 6 wbs_dat_o[13]
port 570 nsew signal tristate
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 571 nsew signal tristate
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 572 nsew signal tristate
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 573 nsew signal tristate
rlabel metal2 s 7700 0 7756 800 6 wbs_dat_o[17]
port 574 nsew signal tristate
rlabel metal2 s 8084 0 8140 800 6 wbs_dat_o[18]
port 575 nsew signal tristate
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_o[19]
port 576 nsew signal tristate
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 577 nsew signal tristate
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 578 nsew signal tristate
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 579 nsew signal tristate
rlabel metal2 s 9524 0 9580 800 6 wbs_dat_o[22]
port 580 nsew signal tristate
rlabel metal2 s 9908 0 9964 800 6 wbs_dat_o[23]
port 581 nsew signal tristate
rlabel metal2 s 10292 0 10348 800 6 wbs_dat_o[24]
port 582 nsew signal tristate
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 583 nsew signal tristate
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 584 nsew signal tristate
rlabel metal2 s 11348 0 11404 800 6 wbs_dat_o[27]
port 585 nsew signal tristate
rlabel metal2 s 11732 0 11788 800 6 wbs_dat_o[28]
port 586 nsew signal tristate
rlabel metal2 s 12116 0 12172 800 6 wbs_dat_o[29]
port 587 nsew signal tristate
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 588 nsew signal tristate
rlabel metal2 s 12500 0 12556 800 6 wbs_dat_o[30]
port 589 nsew signal tristate
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 590 nsew signal tristate
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 591 nsew signal tristate
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 592 nsew signal tristate
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 593 nsew signal tristate
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 594 nsew signal tristate
rlabel metal2 s 4052 0 4108 800 6 wbs_dat_o[7]
port 595 nsew signal tristate
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 596 nsew signal tristate
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 597 nsew signal tristate
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 598 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 599 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 600 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 601 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 602 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 603 nsew signal input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 604 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 606 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 607 nsew ground bidirectional
rlabel metal4 s 35636 2664 35956 57276 6 vccd2
port 608 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 57276 6 vccd2
port 609 nsew power bidirectional
rlabel metal4 s 50996 2664 51316 57276 6 vssd2
port 610 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 57276 6 vssd2
port 611 nsew ground bidirectional
rlabel metal4 s 36296 2664 36616 57276 6 vdda1
port 612 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 57276 6 vdda1
port 613 nsew power bidirectional
rlabel metal4 s 51656 2664 51976 57276 6 vssa1
port 614 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 57276 6 vssa1
port 615 nsew ground bidirectional
rlabel metal4 s 36956 2664 37276 57276 6 vdda2
port 616 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 57276 6 vdda2
port 617 nsew power bidirectional
rlabel metal4 s 52316 2664 52636 57276 6 vssa2
port 618 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 57276 6 vssa2
port 619 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
