magic
tech sky130A
timestamp 1621278052
<< end >>
