magic
tech sky130A
magscale 1 2
timestamp 1636962390
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 2304 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1425 48 1455 132
rect 1713 48 1743 132
rect 2001 48 2031 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1425 450 1455 618
rect 1713 450 1743 618
rect 2001 450 2031 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 355 134 413 146
rect 355 132 367 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 739 134 797 146
rect 739 132 751 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 100 751 132
rect 785 132 797 134
rect 931 134 989 146
rect 931 132 943 134
rect 785 100 849 132
rect 591 48 849 100
rect 879 100 943 132
rect 977 132 989 134
rect 1267 134 1325 146
rect 977 100 1037 132
rect 879 48 1037 100
rect 1267 100 1279 134
rect 1313 132 1325 134
rect 1603 134 1661 146
rect 1603 132 1615 134
rect 1313 100 1425 132
rect 1267 48 1425 100
rect 1455 100 1615 132
rect 1649 132 1661 134
rect 1795 134 1853 146
rect 1795 132 1807 134
rect 1649 100 1713 132
rect 1455 48 1713 100
rect 1743 100 1807 132
rect 1841 132 1853 134
rect 2083 134 2141 146
rect 2083 132 2095 134
rect 1841 100 2001 132
rect 1743 48 2001 100
rect 2031 100 2095 132
rect 2129 132 2141 134
rect 2129 100 2189 132
rect 2031 48 2189 100
<< pdiff >>
rect 115 566 273 618
rect 115 532 175 566
rect 209 532 273 566
rect 115 450 273 532
rect 303 485 561 618
rect 303 451 367 485
rect 401 451 561 485
rect 303 450 561 451
rect 591 485 849 618
rect 591 451 751 485
rect 785 451 849 485
rect 591 450 849 451
rect 879 593 1037 618
rect 879 559 943 593
rect 977 559 1037 593
rect 879 450 1037 559
rect 1267 485 1425 618
rect 1267 451 1279 485
rect 1313 451 1425 485
rect 1267 450 1425 451
rect 1455 566 1713 618
rect 1455 532 1519 566
rect 1553 532 1713 566
rect 1455 450 1713 532
rect 1743 593 2001 618
rect 1743 559 1807 593
rect 1841 559 2001 593
rect 1743 450 2001 559
rect 2031 485 2189 618
rect 2031 451 2095 485
rect 2129 451 2189 485
rect 2031 450 2189 451
rect 355 439 413 450
rect 739 439 797 450
rect 1267 439 1325 450
rect 2083 439 2141 450
<< ndiffc >>
rect 127 100 161 134
rect 367 100 401 134
rect 751 100 785 134
rect 943 100 977 134
rect 1279 100 1313 134
rect 1615 100 1649 134
rect 1807 100 1841 134
rect 2095 100 2129 134
<< pdiffc >>
rect 175 532 209 566
rect 367 451 401 485
rect 751 451 785 485
rect 943 559 977 593
rect 1279 451 1313 485
rect 1519 532 1553 566
rect 1807 559 1841 593
rect 2095 451 2129 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1425 618 1455 644
rect 1713 618 1743 644
rect 2001 618 2031 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1425 418 1455 450
rect 1713 418 1743 450
rect 2001 418 2031 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1425 132 1455 165
rect 1713 132 1743 165
rect 2001 132 2031 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1425 22 1455 48
rect 1713 22 1743 48
rect 2001 22 2031 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 1999 181 2033 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2304 683
rect 31 618 2273 649
rect 927 593 993 618
rect 159 566 225 582
rect 159 532 175 566
rect 209 532 225 566
rect 927 559 943 593
rect 977 559 993 593
rect 1791 593 1857 618
rect 927 543 993 559
rect 1503 566 1569 582
rect 159 516 225 532
rect 1503 532 1519 566
rect 1553 532 1569 566
rect 1791 559 1807 593
rect 1841 559 1857 593
rect 1791 543 1857 559
rect 1503 516 1569 532
rect 351 485 417 501
rect 351 452 367 485
rect 355 451 367 452
rect 401 451 417 485
rect 735 485 801 501
rect 355 435 417 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 367 377 401 435
rect 255 215 321 231
rect 255 181 271 215
rect 305 184 321 215
rect 305 181 317 184
rect 255 165 317 181
rect 367 150 401 343
rect 735 451 751 485
rect 785 452 801 485
rect 1263 485 1329 501
rect 2079 485 2145 501
rect 785 451 797 452
rect 735 435 797 451
rect 1263 451 1279 485
rect 1313 451 1329 485
rect 1263 435 1329 451
rect 2079 452 2095 485
rect 463 296 497 424
rect 1423 418 1457 451
rect 2083 451 2095 452
rect 2129 451 2145 485
rect 2083 435 2145 451
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 559 231 593 352
rect 847 242 881 352
rect 655 231 881 242
rect 1423 231 1457 352
rect 1711 231 1745 352
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 655 215 897 231
rect 655 208 847 215
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 351 134 417 150
rect 351 100 367 134
rect 401 100 417 134
rect 655 134 689 208
rect 831 181 847 208
rect 881 184 897 215
rect 1407 215 1473 231
rect 881 181 893 184
rect 831 165 893 181
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1695 215 1761 231
rect 1695 184 1711 215
rect 1407 165 1473 181
rect 1699 181 1711 184
rect 1745 184 1761 215
rect 1983 215 2049 231
rect 1745 181 1757 184
rect 1699 165 1757 181
rect 1983 181 1999 215
rect 2033 184 2049 215
rect 2033 181 2045 184
rect 1983 165 2045 181
rect 735 134 797 150
rect 735 100 751 134
rect 785 131 797 134
rect 927 134 993 150
rect 785 100 801 131
rect 351 84 417 100
rect 735 84 801 100
rect 927 100 943 134
rect 977 100 993 134
rect 927 84 993 100
rect 1263 134 1329 150
rect 1263 100 1279 134
rect 1313 100 1329 134
rect 1263 84 1329 100
rect 1599 134 1665 150
rect 1599 100 1615 134
rect 1649 100 1665 134
rect 1599 84 1665 100
rect 1791 134 1857 150
rect 1791 100 1807 134
rect 1841 100 1857 134
rect 1791 84 1857 100
rect 2079 134 2145 150
rect 2079 100 2095 134
rect 2129 100 2145 134
rect 2079 84 2145 100
rect 943 48 977 84
rect 1807 48 1841 84
rect 31 17 2273 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2304 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 175 532 209 566
rect 1519 532 1553 566
rect 1807 559 1841 593
rect 271 368 305 402
rect 367 343 401 377
rect 271 181 305 215
rect 463 424 497 458
rect 751 451 785 485
rect 1279 451 1313 485
rect 1423 451 1457 485
rect 2095 451 2129 485
rect 1999 368 2033 402
rect 463 262 497 296
rect 559 181 593 215
rect 127 100 161 134
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 655 100 689 134
rect 751 100 785 134
rect 1279 100 1313 134
rect 1615 100 1649 134
rect 2095 100 2129 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2304 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2304 683
rect 0 618 2304 649
rect 1795 593 1853 618
rect 163 566 221 578
rect 163 532 175 566
rect 209 563 221 566
rect 1507 566 1565 578
rect 1507 563 1519 566
rect 209 535 1519 563
rect 209 532 221 535
rect 163 520 221 532
rect 1507 532 1519 535
rect 1553 532 1565 566
rect 1795 559 1807 593
rect 1841 559 1853 593
rect 1795 547 1853 559
rect 1507 520 1565 532
rect 739 485 797 497
rect 130 470 494 482
rect 130 458 509 470
rect 130 454 463 458
rect 130 146 158 454
rect 451 424 463 454
rect 497 424 509 458
rect 739 451 751 485
rect 785 482 797 485
rect 1267 485 1325 497
rect 1267 482 1279 485
rect 785 454 1279 482
rect 785 451 797 454
rect 739 439 797 451
rect 1267 451 1279 454
rect 1313 451 1325 485
rect 1267 439 1325 451
rect 1411 485 1469 497
rect 1411 451 1423 485
rect 1457 482 1469 485
rect 2083 485 2141 497
rect 2083 482 2095 485
rect 1457 454 2095 482
rect 1457 451 1469 454
rect 1411 439 1469 451
rect 2083 451 2095 454
rect 2129 451 2141 485
rect 2083 439 2141 451
rect 259 402 317 414
rect 451 412 509 424
rect 259 368 271 402
rect 305 368 317 402
rect 1987 402 2045 414
rect 259 356 317 368
rect 355 377 413 389
rect 274 227 302 356
rect 355 343 367 377
rect 401 374 413 377
rect 1987 374 1999 402
rect 401 368 1999 374
rect 2033 368 2045 402
rect 401 356 2045 368
rect 401 346 2030 356
rect 401 343 413 346
rect 355 331 413 343
rect 451 296 509 308
rect 451 262 463 296
rect 497 293 509 296
rect 497 265 1838 293
rect 497 262 509 265
rect 451 250 509 262
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 212 605 215
rect 1699 215 1757 227
rect 1699 212 1711 215
rect 593 184 1711 212
rect 593 181 605 184
rect 547 169 605 181
rect 1699 181 1711 184
rect 1745 181 1757 215
rect 1699 169 1757 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 274 131 302 169
rect 643 134 701 146
rect 643 131 655 134
rect 274 103 655 131
rect 115 88 173 100
rect 643 100 655 103
rect 689 100 701 134
rect 643 88 701 100
rect 739 134 797 146
rect 739 100 751 134
rect 785 131 797 134
rect 1267 134 1325 146
rect 1267 131 1279 134
rect 785 103 1279 131
rect 785 100 797 103
rect 739 88 797 100
rect 1267 100 1279 103
rect 1313 100 1325 134
rect 1267 88 1325 100
rect 1603 134 1661 146
rect 1603 100 1615 134
rect 1649 131 1661 134
rect 1810 131 1838 265
rect 2002 227 2030 346
rect 1987 215 2045 227
rect 1987 181 1999 215
rect 2033 181 2045 215
rect 1987 169 2045 181
rect 2098 146 2126 439
rect 1649 103 1838 131
rect 2083 134 2141 146
rect 1649 100 1661 103
rect 1603 88 1661 100
rect 2083 100 2095 134
rect 2129 100 2141 134
rect 2083 88 2141 100
rect 0 17 2304 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2304 17
rect 0 -48 2304 -17
<< labels >>
rlabel metal1 0 618 2304 714 0 VPWR
port 4 se
rlabel metal1 0 618 2304 714 0 VPWR
port 4 se
rlabel metal1 0 -48 2304 48 0 VGND
port 3 se
rlabel metal1 0 -48 2304 48 0 VGND
port 3 se
rlabel metal1 2083 88 2141 146 0 C
port 2 se
rlabel metal1 2098 146 2126 439 0 C
port 2 se
rlabel metal1 1411 439 1469 454 0 C
port 2 se
rlabel metal1 2083 439 2141 454 0 C
port 2 se
rlabel metal1 1411 454 2141 482 0 C
port 2 se
rlabel metal1 1411 482 1469 497 0 C
port 2 se
rlabel metal1 2083 482 2141 497 0 C
port 2 se
rlabel metal1 547 169 605 184 0 B
port 1 se
rlabel metal1 1699 169 1757 184 0 B
port 1 se
rlabel metal1 547 184 1757 212 0 B
port 1 se
rlabel metal1 547 212 605 227 0 B
port 1 se
rlabel metal1 1699 212 1757 227 0 B
port 1 se
rlabel metal1 643 88 701 103 0 A
port 0 se
rlabel metal1 274 103 701 131 0 A
port 0 se
rlabel metal1 643 131 701 146 0 A
port 0 se
rlabel metal1 274 131 302 169 0 A
port 0 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel locali 0 -17 2304 17 4 VGND
port 3 se ground default abutment
rlabel locali 31 17 2273 48 4 VGND
port 3 se ground default abutment
rlabel locali 0 649 2304 683 4 VPWR
port 4 se power default abutment
rlabel locali 31 618 2273 649 4 VGND
port 3 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 2304 666
<< end >>
