MACRO INVX8
 CLASS CORE ;
 FOREIGN INVX8 0 0 ;
 SIZE 7.2 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 7.20000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 7.20000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 3.69500000 0.44000000 3.98500000 0.51500000 ;
        RECT 6.09500000 0.44000000 6.38500000 0.51500000 ;
        RECT 3.69500000 0.51500000 6.38500000 0.65500000 ;
        RECT 0.81500000 0.44000000 1.10500000 0.73000000 ;
        RECT 3.69500000 0.65500000 3.98500000 0.73000000 ;
        RECT 6.09500000 0.65500000 6.38500000 0.73000000 ;
        RECT 0.89000000 0.73000000 1.03000000 2.19500000 ;
        RECT 6.17000000 0.73000000 6.31000000 2.19500000 ;
        RECT 0.81500000 2.19500000 1.10500000 2.27000000 ;
        RECT 3.69500000 2.19500000 3.98500000 2.27000000 ;
        RECT 6.09500000 2.19500000 6.38500000 2.27000000 ;
        RECT 0.81500000 2.27000000 6.38500000 2.41000000 ;
        RECT 0.81500000 2.41000000 1.10500000 2.48500000 ;
        RECT 3.69500000 2.41000000 3.98500000 2.48500000 ;
        RECT 6.09500000 2.41000000 6.38500000 2.48500000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 2.73500000 0.84500000 3.02500000 1.13500000 ;
        RECT 4.17500000 0.84500000 4.46500000 1.13500000 ;
        RECT 5.61500000 0.84500000 5.90500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 2.81000000 1.13500000 2.95000000 1.78000000 ;
        RECT 4.25000000 1.13500000 4.39000000 1.78000000 ;
        RECT 5.69000000 1.13500000 5.83000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 1.85500000 ;
        RECT 2.73500000 1.78000000 3.02500000 1.85500000 ;
        RECT 4.17500000 1.78000000 4.46500000 1.85500000 ;
        RECT 5.61500000 1.78000000 5.90500000 1.85500000 ;
        RECT 1.29500000 1.85500000 5.90500000 1.99500000 ;
        RECT 1.29500000 1.99500000 1.58500000 2.07000000 ;
        RECT 2.73500000 1.99500000 3.02500000 2.07000000 ;
        RECT 4.17500000 1.99500000 4.46500000 2.07000000 ;
        RECT 5.61500000 1.99500000 5.90500000 2.07000000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 5.67500000 0.90500000 5.84500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 0.87500000 2.25500000 1.04500000 2.42500000 ;
     RECT 3.75500000 2.25500000 3.92500000 2.42500000 ;
     RECT 6.15500000 2.25500000 6.32500000 2.42500000 ;
     RECT 1.83500000 2.84000000 2.00500000 3.01000000 ;
     RECT 4.71500000 2.84000000 4.88500000 3.01000000 ;

    LAYER ndiffc ;
     RECT 1.83500000 0.32000000 2.00500000 0.49000000 ;
     RECT 4.71500000 0.32000000 4.88500000 0.49000000 ;
     RECT 0.87500000 0.50000000 1.04500000 0.67000000 ;
     RECT 3.75500000 0.50000000 3.92500000 0.67000000 ;
     RECT 6.15500000 0.50000000 6.32500000 0.67000000 ;

    LAYER li1 ;
     RECT 1.83500000 0.09500000 2.00500000 0.24000000 ;
     RECT 1.75500000 0.24000000 2.08500000 0.57000000 ;
     RECT 4.71500000 0.09500000 4.88500000 0.24000000 ;
     RECT 4.63500000 0.24000000 4.96500000 0.57000000 ;
     RECT 0.79500000 0.42000000 1.12500000 0.75000000 ;
     RECT 3.67500000 0.42000000 4.00500000 0.75000000 ;
     RECT 6.07500000 0.42000000 6.40500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 2.71500000 0.82500000 3.04500000 1.15500000 ;
     RECT 4.15500000 0.82500000 4.48500000 1.15500000 ;
     RECT 5.59500000 0.82500000 5.92500000 1.15500000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 2.71500000 1.76000000 3.04500000 2.09000000 ;
     RECT 4.15500000 1.76000000 4.48500000 2.09000000 ;
     RECT 5.59500000 1.76000000 5.92500000 2.09000000 ;
     RECT 0.79500000 2.17500000 1.12500000 2.50500000 ;
     RECT 3.67500000 2.17500000 4.00500000 2.50500000 ;
     RECT 6.07500000 2.17500000 6.40500000 2.50500000 ;
     RECT 1.75500000 2.76000000 2.08500000 3.09000000 ;
     RECT 4.63500000 2.76000000 4.96500000 3.09000000 ;

    LAYER viali ;
     RECT 1.83500000 0.09500000 2.00500000 0.26500000 ;
     RECT 4.71500000 0.09500000 4.88500000 0.26500000 ;
     RECT 0.87500000 0.50000000 1.04500000 0.67000000 ;
     RECT 3.75500000 0.50000000 3.92500000 0.67000000 ;
     RECT 6.15500000 0.50000000 6.32500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 5.67500000 0.90500000 5.84500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;
     RECT 0.87500000 2.25500000 1.04500000 2.42500000 ;
     RECT 3.75500000 2.25500000 3.92500000 2.42500000 ;
     RECT 6.15500000 2.25500000 6.32500000 2.42500000 ;
     RECT 1.83500000 2.84000000 2.00500000 3.01000000 ;
     RECT 4.71500000 2.84000000 4.88500000 3.01000000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 7.20000000 0.24000000 ;
     RECT 1.77500000 0.24000000 2.06500000 0.32500000 ;
     RECT 4.65500000 0.24000000 4.94500000 0.32500000 ;
     RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
     RECT 2.73500000 0.84500000 3.02500000 1.13500000 ;
     RECT 4.17500000 0.84500000 4.46500000 1.13500000 ;
     RECT 5.61500000 0.84500000 5.90500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
     RECT 2.81000000 1.13500000 2.95000000 1.78000000 ;
     RECT 4.25000000 1.13500000 4.39000000 1.78000000 ;
     RECT 5.69000000 1.13500000 5.83000000 1.78000000 ;
     RECT 1.29500000 1.78000000 1.58500000 1.85500000 ;
     RECT 2.73500000 1.78000000 3.02500000 1.85500000 ;
     RECT 4.17500000 1.78000000 4.46500000 1.85500000 ;
     RECT 5.61500000 1.78000000 5.90500000 1.85500000 ;
     RECT 1.29500000 1.85500000 5.90500000 1.99500000 ;
     RECT 1.29500000 1.99500000 1.58500000 2.07000000 ;
     RECT 2.73500000 1.99500000 3.02500000 2.07000000 ;
     RECT 4.17500000 1.99500000 4.46500000 2.07000000 ;
     RECT 5.61500000 1.99500000 5.90500000 2.07000000 ;
     RECT 3.69500000 0.44000000 3.98500000 0.51500000 ;
     RECT 6.09500000 0.44000000 6.38500000 0.51500000 ;
     RECT 3.69500000 0.51500000 6.38500000 0.65500000 ;
     RECT 0.81500000 0.44000000 1.10500000 0.73000000 ;
     RECT 3.69500000 0.65500000 3.98500000 0.73000000 ;
     RECT 6.09500000 0.65500000 6.38500000 0.73000000 ;
     RECT 0.89000000 0.73000000 1.03000000 2.19500000 ;
     RECT 6.17000000 0.73000000 6.31000000 2.19500000 ;
     RECT 0.81500000 2.19500000 1.10500000 2.27000000 ;
     RECT 3.69500000 2.19500000 3.98500000 2.27000000 ;
     RECT 6.09500000 2.19500000 6.38500000 2.27000000 ;
     RECT 0.81500000 2.27000000 6.38500000 2.41000000 ;
     RECT 0.81500000 2.41000000 1.10500000 2.48500000 ;
     RECT 3.69500000 2.41000000 3.98500000 2.48500000 ;
     RECT 6.09500000 2.41000000 6.38500000 2.48500000 ;
     RECT 1.77500000 2.78000000 2.06500000 3.09000000 ;
     RECT 4.65500000 2.78000000 4.94500000 3.09000000 ;
     RECT 0.00000000 3.09000000 7.20000000 3.57000000 ;

 END
END INVX8
