magic
tech sky130A
timestamp 1621276911
<< end >>
