VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OR2X1
  CLASS CORE ;
  FOREIGN OR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.780 1.585 2.070 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 1.780 3.025 2.070 ;
        RECT 2.810 1.540 2.950 1.780 ;
        RECT 2.735 1.250 3.025 1.540 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA 0.914200 ;
    PORT
      LAYER met1 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 3.215 0.440 3.505 0.730 ;
        RECT 0.650 0.240 0.790 0.440 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 3.215 2.735 3.505 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.155 3.090 5.605 3.245 ;
        RECT 3.195 2.715 3.525 3.090 ;
      LAYER mcon ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 3.275 2.795 3.445 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 4.655 2.195 4.945 2.485 ;
        RECT 4.730 0.730 4.870 2.195 ;
        RECT 4.655 0.440 4.945 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 5.760 3.330 ;
      LAYER li1 ;
        RECT 0.795 2.260 1.125 2.505 ;
        RECT 0.795 2.175 1.105 2.260 ;
        RECT 4.635 2.175 4.965 2.505 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 2.005 4.465 2.090 ;
        RECT 4.155 1.760 4.485 2.005 ;
        RECT 1.355 1.155 1.525 1.760 ;
        RECT 2.795 1.155 2.965 1.480 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 2.715 0.920 3.045 1.155 ;
        RECT 2.735 0.825 3.045 0.920 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 4.155 0.825 4.465 0.920 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 2.235 0.420 2.565 0.750 ;
        RECT 3.215 0.655 3.525 0.750 ;
        RECT 3.195 0.420 3.525 0.655 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 0.155 0.085 5.605 0.240 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.875 2.255 1.045 2.425 ;
        RECT 4.715 2.255 4.885 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 2.795 1.310 2.965 1.480 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 2.315 0.500 2.485 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
      LAYER met1 ;
        RECT 0.815 2.195 1.105 2.485 ;
        RECT 0.890 1.060 1.030 2.195 ;
        RECT 4.175 1.780 4.465 2.070 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 4.175 1.060 4.465 1.135 ;
        RECT 0.890 0.920 4.465 1.060 ;
        RECT 2.330 0.730 2.470 0.920 ;
        RECT 4.175 0.845 4.465 0.920 ;
        RECT 2.255 0.440 2.545 0.730 ;
  END
END OR2X1
END LIBRARY

