VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 7.200 3.570 ;
        RECT 1.780 3.010 2.070 3.090 ;
        RECT 1.780 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.070 3.010 ;
        RECT 1.780 2.780 2.070 2.840 ;
        RECT 4.660 3.010 4.950 3.090 ;
        RECT 4.660 2.840 4.720 3.010 ;
        RECT 4.890 2.840 4.950 3.010 ;
        RECT 4.660 2.780 4.950 2.840 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.270 2.070 0.330 ;
        RECT 1.780 0.240 1.840 0.270 ;
        RECT 2.010 0.240 2.070 0.270 ;
        RECT 4.660 0.270 4.950 0.330 ;
        RECT 4.660 0.240 4.720 0.270 ;
        RECT 4.890 0.240 4.950 0.270 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.820 2.410 1.110 2.490 ;
        RECT 3.700 2.410 3.990 2.490 ;
        RECT 6.100 2.410 6.390 2.490 ;
        RECT 0.820 2.270 6.390 2.410 ;
        RECT 0.820 2.200 1.110 2.270 ;
        RECT 3.700 2.200 3.990 2.270 ;
        RECT 6.100 2.200 6.390 2.270 ;
        RECT 0.890 0.730 1.030 2.200 ;
        RECT 6.170 0.730 6.310 2.200 ;
        RECT 0.820 0.440 1.110 0.730 ;
        RECT 3.700 0.660 3.990 0.730 ;
        RECT 6.100 0.660 6.390 0.730 ;
        RECT 3.700 0.520 6.390 0.660 ;
        RECT 3.700 0.440 3.990 0.520 ;
        RECT 6.100 0.440 6.390 0.520 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 2.000 1.590 2.070 ;
        RECT 2.740 2.000 3.030 2.070 ;
        RECT 4.180 2.000 4.470 2.070 ;
        RECT 5.620 2.000 5.910 2.070 ;
        RECT 1.300 1.860 5.910 2.000 ;
        RECT 1.300 1.780 1.590 1.860 ;
        RECT 2.740 1.780 3.030 1.860 ;
        RECT 4.180 1.780 4.470 1.860 ;
        RECT 5.620 1.780 5.910 1.860 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 5.690 1.140 5.830 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
        RECT 2.740 0.850 3.030 1.140 ;
        RECT 4.180 0.850 4.470 1.140 ;
        RECT 5.620 0.850 5.910 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 3.010 2.090 3.090 ;
        RECT 1.760 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.090 3.010 ;
        RECT 1.760 2.760 2.090 2.840 ;
        RECT 4.640 3.010 4.970 3.090 ;
        RECT 4.640 2.840 4.720 3.010 ;
        RECT 4.890 2.840 4.970 3.010 ;
        RECT 4.640 2.760 4.970 2.840 ;
        RECT 0.800 2.430 1.130 2.510 ;
        RECT 0.800 2.260 0.880 2.430 ;
        RECT 1.050 2.260 1.130 2.430 ;
        RECT 0.800 2.180 1.130 2.260 ;
        RECT 3.680 2.430 4.010 2.510 ;
        RECT 3.680 2.260 3.760 2.430 ;
        RECT 3.930 2.260 4.010 2.430 ;
        RECT 6.080 2.430 6.410 2.510 ;
        RECT 6.080 2.260 6.160 2.430 ;
        RECT 6.330 2.260 6.410 2.430 ;
        RECT 3.680 2.180 3.990 2.260 ;
        RECT 6.100 2.180 6.410 2.260 ;
        RECT 1.300 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 2.010 5.930 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.920 4.240 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.180 0.910 4.240 0.920 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.180 0.830 4.490 0.910 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.600 0.830 5.930 0.910 ;
        RECT 0.800 0.670 1.110 0.750 ;
        RECT 0.800 0.500 0.880 0.670 ;
        RECT 1.050 0.660 1.110 0.670 ;
        RECT 3.680 0.670 4.010 0.750 ;
        RECT 1.050 0.500 1.130 0.660 ;
        RECT 0.800 0.420 1.130 0.500 ;
        RECT 1.760 0.490 2.090 0.570 ;
        RECT 1.760 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.090 0.490 ;
        RECT 3.680 0.500 3.760 0.670 ;
        RECT 3.930 0.500 4.010 0.670 ;
        RECT 6.100 0.670 6.410 0.750 ;
        RECT 6.100 0.660 6.160 0.670 ;
        RECT 3.680 0.420 4.010 0.500 ;
        RECT 4.640 0.490 4.970 0.570 ;
        RECT 1.760 0.270 2.090 0.320 ;
        RECT 1.760 0.240 1.840 0.270 ;
        RECT 2.010 0.240 2.090 0.270 ;
        RECT 4.640 0.320 4.720 0.490 ;
        RECT 4.890 0.320 4.970 0.490 ;
        RECT 6.080 0.500 6.160 0.660 ;
        RECT 6.330 0.500 6.410 0.670 ;
        RECT 6.080 0.420 6.410 0.500 ;
        RECT 4.640 0.270 4.970 0.320 ;
        RECT 4.640 0.240 4.720 0.270 ;
        RECT 4.890 0.240 4.970 0.270 ;
  END
END INVX8
END LIBRARY

