VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX1
  CLASS CORE ;
  FOREIGN INVX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 2.880 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.880 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 2.150 2.070 2.440 ;
        RECT 1.850 0.690 1.990 2.150 ;
        RECT 1.780 0.400 2.070 0.690 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END A
END INVX1
END LIBRARY

