magic
tech sky130A
magscale 1 2
timestamp 1624917773
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 2016 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
rect 1713 48 1743 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
rect 1713 450 1743 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 931 134 989 146
rect 931 132 943 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 102 561 132
rect 303 68 367 102
rect 401 68 561 102
rect 303 48 561 68
rect 591 48 849 132
rect 879 100 943 132
rect 977 132 989 134
rect 1795 134 1853 146
rect 1795 132 1807 134
rect 977 100 1137 132
rect 879 48 1137 100
rect 1167 48 1425 132
rect 1455 102 1713 132
rect 1455 68 1519 102
rect 1553 68 1713 102
rect 1455 48 1713 68
rect 1743 100 1807 132
rect 1841 132 1853 134
rect 1841 100 1901 132
rect 1743 48 1901 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 598 561 618
rect 303 564 367 598
rect 401 564 561 598
rect 303 450 561 564
rect 591 450 849 618
rect 879 485 1137 618
rect 879 451 943 485
rect 977 451 1137 485
rect 879 450 1137 451
rect 1167 450 1425 618
rect 1455 598 1713 618
rect 1455 564 1519 598
rect 1553 564 1713 598
rect 1455 450 1713 564
rect 1743 485 1901 618
rect 1743 451 1807 485
rect 1841 451 1901 485
rect 1743 450 1901 451
rect 115 439 173 450
rect 931 439 989 450
rect 1795 439 1853 450
<< ndiffc >>
rect 127 100 161 134
rect 367 68 401 102
rect 943 100 977 134
rect 1519 68 1553 102
rect 1807 100 1841 134
<< pdiffc >>
rect 127 451 161 485
rect 367 564 401 598
rect 943 451 977 485
rect 1519 564 1553 598
rect 1807 451 1841 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 1713 618 1743 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 1713 418 1743 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 1713 132 1743 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
rect 1713 22 1743 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 31 618 1985 649
rect 351 598 417 618
rect 351 564 367 598
rect 401 564 417 598
rect 1503 598 1569 618
rect 351 548 417 564
rect 1503 564 1519 598
rect 1553 564 1569 598
rect 1503 548 1569 564
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 559 418 593 532
rect 927 485 993 501
rect 927 452 943 485
rect 847 418 881 451
rect 931 451 943 452
rect 977 451 993 485
rect 1791 485 1857 501
rect 1791 452 1807 485
rect 931 435 993 451
rect 1795 451 1807 452
rect 1841 451 1857 485
rect 1795 435 1857 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 559 323 593 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 184 897 215
rect 881 181 893 184
rect 831 165 893 181
rect 943 150 977 435
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1711 231 1745 352
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 927 134 993 150
rect 111 84 177 100
rect 351 102 417 118
rect 351 68 367 102
rect 401 68 417 102
rect 927 100 943 134
rect 977 100 993 134
rect 1795 134 1857 150
rect 1795 131 1807 134
rect 927 84 993 100
rect 1503 102 1569 118
rect 351 48 417 68
rect 1503 68 1519 102
rect 1553 68 1569 102
rect 1791 100 1807 131
rect 1841 100 1857 134
rect 1791 84 1857 100
rect 1503 48 1569 68
rect 31 17 1985 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 367 564 401 598
rect 559 532 593 566
rect 127 451 161 485
rect 847 451 881 485
rect 1807 451 1841 485
rect 271 368 305 402
rect 559 289 593 323
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 127 100 161 134
rect 367 68 401 102
rect 943 100 977 134
rect 1519 68 1553 102
rect 1807 100 1841 134
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 714
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 618 2016 649
rect 355 598 413 618
rect 355 564 367 598
rect 401 564 413 598
rect 355 552 413 564
rect 547 566 605 578
rect 547 532 559 566
rect 593 563 605 566
rect 593 535 1742 563
rect 593 532 605 535
rect 547 520 605 532
rect 115 485 173 497
rect 115 451 127 485
rect 161 482 173 485
rect 835 485 893 497
rect 835 482 847 485
rect 161 454 847 482
rect 161 451 173 454
rect 115 439 173 451
rect 835 451 847 454
rect 881 482 893 485
rect 881 454 1262 482
rect 881 451 893 454
rect 835 439 893 451
rect 130 146 158 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 399 317 402
rect 1123 402 1181 414
rect 1123 399 1135 402
rect 305 371 1135 399
rect 305 368 317 371
rect 259 356 317 368
rect 274 227 302 356
rect 547 323 605 335
rect 547 289 559 323
rect 593 289 605 323
rect 547 277 605 289
rect 562 227 590 277
rect 850 227 878 371
rect 1123 368 1135 371
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 181 605 215
rect 547 169 605 181
rect 835 215 893 227
rect 835 181 847 215
rect 881 181 893 215
rect 835 169 893 181
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 212 1181 215
rect 1234 212 1262 454
rect 1714 414 1742 535
rect 1795 485 1853 497
rect 1795 451 1807 485
rect 1841 451 1853 485
rect 1795 439 1853 451
rect 1411 402 1469 414
rect 1411 368 1423 402
rect 1457 368 1469 402
rect 1411 356 1469 368
rect 1699 402 1757 414
rect 1699 368 1711 402
rect 1745 368 1757 402
rect 1699 356 1757 368
rect 1426 227 1454 356
rect 1169 184 1262 212
rect 1411 215 1469 227
rect 1169 181 1181 184
rect 1123 169 1181 181
rect 1411 181 1423 215
rect 1457 212 1469 215
rect 1810 212 1838 439
rect 1457 184 1838 212
rect 1457 181 1469 184
rect 1411 169 1469 181
rect 1810 146 1838 184
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 931 134 989 146
rect 115 88 173 100
rect 355 102 413 114
rect 355 68 367 102
rect 401 68 413 102
rect 931 100 943 134
rect 977 100 989 134
rect 1795 134 1853 146
rect 931 88 989 100
rect 1507 102 1565 114
rect 355 48 413 68
rect 1507 68 1519 102
rect 1553 68 1565 102
rect 1795 100 1807 134
rect 1841 100 1853 134
rect 1795 88 1853 100
rect 1507 48 1565 68
rect 0 17 2016 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -48 2016 -17
<< labels >>
rlabel metal1 0 618 2016 714 0 VPWR
port 3 se
rlabel metal1 0 618 2016 714 0 VPWR
port 3 se
rlabel metal1 0 -48 2016 48 0 VGND
port 2 se
rlabel metal1 931 88 989 146 0 Y
port 4 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 835 169 893 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 259 356 317 371 0 A
port 0 se
rlabel metal1 850 227 878 371 0 A
port 0 se
rlabel metal1 1123 356 1181 371 0 A
port 0 se
rlabel metal1 259 371 1181 399 0 A
port 0 se
rlabel metal1 259 399 317 414 0 A
port 0 se
rlabel metal1 1123 399 1181 414 0 A
port 0 se
rlabel metal1 547 169 605 227 0 B
port 1 se
rlabel metal1 562 227 590 277 0 B
port 1 se
rlabel metal1 547 277 605 335 0 B
port 1 se
rlabel locali 0 -17 2016 17 4 VGND
port 2 se ground default abutment
rlabel locali 31 17 1985 48 4 VGND
port 2 se ground default abutment
rlabel locali 0 649 2016 683 4 VPWR
port 3 se power default abutment
rlabel locali 31 618 1985 649 4 VGND
port 2 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 2016 666
<< end >>
