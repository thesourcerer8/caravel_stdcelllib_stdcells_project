VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 0.580 2.970 0.870 3.090 ;
        RECT 0.580 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.870 2.970 ;
        RECT 0.580 2.740 0.870 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 0.560 2.970 0.890 3.090 ;
        RECT 0.560 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.890 2.970 ;
        RECT 0.560 2.720 0.890 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.760 0.670 2.090 0.750 ;
        RECT 1.760 0.500 1.840 0.670 ;
        RECT 2.010 0.500 2.090 0.670 ;
        RECT 1.760 0.420 2.090 0.500 ;
        RECT 1.840 0.240 2.010 0.420 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.220 2.200 3.510 2.490 ;
        RECT 3.290 0.730 3.430 2.200 ;
        RECT 0.820 0.660 1.110 0.730 ;
        RECT 3.220 0.660 3.510 0.730 ;
        RECT 0.820 0.520 3.510 0.660 ;
        RECT 0.820 0.440 1.110 0.520 ;
        RECT 3.220 0.440 3.510 0.520 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 2.740 0.850 3.030 1.140 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 3.200 2.430 3.530 2.510 ;
        RECT 3.200 2.260 3.280 2.430 ;
        RECT 3.450 2.260 3.530 2.430 ;
        RECT 3.220 2.180 3.530 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.920 1.610 1.080 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 1.530 0.910 1.590 0.920 ;
        RECT 1.280 0.830 1.590 0.910 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.920 3.050 1.080 ;
        RECT 2.970 0.910 3.030 0.920 ;
        RECT 2.720 0.830 3.030 0.910 ;
        RECT 0.800 0.670 1.110 0.750 ;
        RECT 0.800 0.500 0.880 0.670 ;
        RECT 1.050 0.660 1.110 0.670 ;
        RECT 3.200 0.670 3.530 0.750 ;
        RECT 1.050 0.500 1.130 0.660 ;
        RECT 0.800 0.420 1.130 0.500 ;
        RECT 3.200 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.530 0.670 ;
        RECT 3.200 0.420 3.530 0.500 ;
  END
END NOR2X1
END LIBRARY

