VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 1.385 3.025 1.675 ;
        RECT 2.810 1.135 2.950 1.385 ;
        RECT 2.735 0.845 3.025 1.135 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA 0.562100 ;
    PORT
      LAYER met1 ;
        RECT 3.215 0.440 3.505 0.730 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 0.575 2.735 0.865 3.090 ;
        RECT 3.215 2.735 3.505 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 0.663600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.155 3.215 5.605 3.245 ;
        RECT 0.155 3.090 3.025 3.215 ;
        RECT 3.695 3.090 5.605 3.215 ;
        RECT 0.555 2.715 0.885 3.090 ;
      LAYER mcon ;
        RECT 3.275 3.245 3.445 3.415 ;
        RECT 0.635 2.795 0.805 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 4.655 2.195 4.945 2.485 ;
        RECT 4.730 0.730 4.870 2.195 ;
        RECT 4.655 0.440 4.945 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 5.760 3.330 ;
      LAYER li1 ;
        RECT 3.195 2.715 3.525 3.045 ;
        RECT 1.755 2.260 2.085 2.505 ;
        RECT 4.635 2.260 4.965 2.505 ;
        RECT 1.775 2.175 2.085 2.260 ;
        RECT 4.655 2.175 4.965 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 2.795 1.445 2.965 1.760 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.295 0.825 1.605 0.920 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 4.155 0.825 4.465 0.920 ;
        RECT 0.795 0.420 1.125 0.750 ;
        RECT 3.215 0.655 3.525 0.750 ;
        RECT 3.195 0.420 3.525 0.655 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 0.155 0.085 5.605 0.240 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 3.275 2.795 3.445 2.965 ;
        RECT 1.835 2.255 2.005 2.425 ;
        RECT 4.715 2.255 4.885 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 0.875 0.500 1.045 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 3.275 -0.085 3.445 0.085 ;
      LAYER met1 ;
        RECT 1.775 2.195 2.065 2.485 ;
        RECT 1.850 1.995 1.990 2.195 ;
        RECT 4.175 1.995 4.465 2.070 ;
        RECT 1.850 1.855 4.465 1.995 ;
        RECT 0.815 0.655 1.105 0.730 ;
        RECT 1.850 0.655 1.990 1.855 ;
        RECT 4.175 1.780 4.465 1.855 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 4.175 0.845 4.465 1.135 ;
        RECT 0.815 0.515 1.990 0.655 ;
        RECT 0.815 0.440 1.105 0.515 ;
  END
END AND2X1
END LIBRARY

