VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 12.960 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.960 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 10.660 2.370 11.190 2.440 ;
        RECT 10.660 2.230 12.070 2.370 ;
        RECT 10.660 2.150 11.190 2.230 ;
        RECT 11.930 0.750 12.070 2.230 ;
        RECT 10.900 0.610 11.190 0.690 ;
        RECT 11.690 0.610 12.070 0.750 ;
        RECT 10.900 0.470 11.830 0.610 ;
        RECT 10.900 0.400 11.190 0.470 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.370 2.630 2.950 2.770 ;
        RECT 1.370 2.040 1.510 2.630 ;
        RECT 2.810 2.040 2.950 2.630 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 2.740 1.750 3.030 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END A
END CLKBUF1
END LIBRARY

