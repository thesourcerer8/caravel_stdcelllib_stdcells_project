magic
tech sky130A
timestamp 1621276817
<< end >>
