VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 10.080 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.140 0.660 5.430 0.730 ;
        RECT 6.100 0.660 6.390 0.730 ;
        RECT 5.140 0.520 6.390 0.660 ;
        RECT 5.140 0.440 5.430 0.520 ;
        RECT 6.100 0.440 6.390 0.520 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 8.500 1.780 8.790 2.070 ;
        RECT 2.740 1.470 3.030 1.540 ;
        RECT 8.570 1.470 8.710 1.780 ;
        RECT 2.740 1.330 8.710 1.470 ;
        RECT 2.740 1.250 3.030 1.330 ;
        RECT 8.570 1.140 8.710 1.330 ;
        RECT 8.500 0.850 8.790 1.140 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.390 1.590 1.680 ;
        RECT 1.370 1.140 1.510 1.390 ;
        RECT 1.300 0.930 1.590 1.140 ;
        RECT 1.300 0.850 2.230 0.930 ;
        RECT 1.370 0.790 2.230 0.850 ;
        RECT 2.090 0.660 2.230 0.790 ;
        RECT 4.180 0.660 4.470 0.730 ;
        RECT 2.090 0.520 4.470 0.660 ;
        RECT 4.180 0.440 4.470 0.520 ;
    END
  END A
END XOR2X1
END LIBRARY

