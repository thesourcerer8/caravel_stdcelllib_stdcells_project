MACRO CLKBUF1
 CLASS CORE ;
 FOREIGN CLKBUF1 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 12.96000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 12.96000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 10.89500000 0.39500000 11.18500000 0.47000000 ;
        RECT 10.89500000 0.47000000 11.83000000 0.60500000 ;
        RECT 10.89500000 0.60500000 12.07000000 0.61000000 ;
        RECT 10.89500000 0.61000000 11.18500000 0.68500000 ;
        RECT 11.69000000 0.61000000 12.07000000 0.74500000 ;
        RECT 10.65500000 2.15000000 11.18500000 2.22500000 ;
        RECT 11.93000000 0.74500000 12.07000000 2.22500000 ;
        RECT 10.65500000 2.22500000 12.07000000 2.36500000 ;
        RECT 10.65500000 2.36500000 11.18500000 2.44000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.29500000 0.80000000 1.58500000 1.09000000 ;
        RECT 1.37000000 1.09000000 1.51000000 1.74500000 ;
        RECT 1.29500000 1.74500000 1.58500000 2.03500000 ;
        RECT 2.73500000 1.74500000 3.02500000 2.03500000 ;
        RECT 1.37000000 2.03500000 1.51000000 2.63000000 ;
        RECT 2.81000000 2.03500000 2.95000000 2.63000000 ;
        RECT 1.37000000 2.63000000 2.95000000 2.77000000 ;
    END
  END A


END CLKBUF1
