magic
tech sky130A
timestamp 1624702590
<< nwell >>
rect 0 179 720 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
<< ndiff >>
rect 82 67 111 73
rect 82 66 88 67
rect 58 50 88 66
rect 105 66 111 67
rect 610 67 639 73
rect 610 66 616 67
rect 105 50 137 66
rect 58 24 137 50
rect 152 24 281 66
rect 296 51 425 66
rect 296 34 328 51
rect 345 34 425 51
rect 296 24 425 34
rect 440 24 569 66
rect 584 50 616 66
rect 633 66 639 67
rect 633 50 663 66
rect 584 24 663 50
<< pdiff >>
rect 58 256 137 309
rect 58 239 88 256
rect 105 239 137 256
rect 58 225 137 239
rect 152 299 281 309
rect 152 282 184 299
rect 201 282 281 299
rect 152 225 281 282
rect 296 283 425 309
rect 296 266 376 283
rect 393 266 425 283
rect 296 225 425 266
rect 440 243 569 309
rect 440 226 520 243
rect 537 226 569 243
rect 440 225 569 226
rect 584 283 663 309
rect 584 266 616 283
rect 633 266 663 283
rect 584 225 663 266
rect 514 220 543 225
<< ndiffc >>
rect 88 50 105 67
rect 328 34 345 51
rect 616 50 633 67
<< pdiffc >>
rect 88 239 105 256
rect 184 282 201 299
rect 376 266 393 283
rect 520 226 537 243
rect 616 266 633 283
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
<< locali >>
rect 0 342 720 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 720 342
rect 0 309 720 325
rect 176 299 209 309
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 368 283 401 291
rect 368 266 376 283
rect 393 266 401 283
rect 80 256 113 264
rect 368 258 401 266
rect 608 283 641 291
rect 608 266 616 283
rect 633 266 641 283
rect 608 258 641 266
rect 80 239 88 256
rect 105 239 113 256
rect 80 231 113 239
rect 512 243 545 251
rect 512 226 520 243
rect 537 226 545 243
rect 512 218 545 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 562 201 593 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 92 593 108
rect 585 91 591 92
rect 560 83 591 91
rect 80 67 111 75
rect 80 50 88 67
rect 105 66 111 67
rect 608 67 641 75
rect 105 50 113 66
rect 80 42 113 50
rect 320 51 353 59
rect 320 34 328 51
rect 345 34 353 51
rect 608 50 616 67
rect 633 50 641 67
rect 608 42 641 50
rect 320 24 353 34
rect 0 9 720 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 720 9
rect 0 -24 720 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 304 325 321 342
rect 352 325 369 342
rect 400 325 417 342
rect 448 325 465 342
rect 496 325 513 342
rect 544 325 561 342
rect 592 325 609 342
rect 640 325 657 342
rect 688 325 705 342
rect 184 282 201 299
rect 376 266 393 283
rect 616 266 633 283
rect 88 239 105 256
rect 520 226 537 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
rect 88 50 105 67
rect 616 50 633 67
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
rect 304 -9 321 9
rect 352 -9 369 9
rect 400 -9 417 9
rect 448 -9 465 9
rect 496 -9 513 9
rect 544 -9 561 9
rect 592 -9 609 9
rect 640 -9 657 9
rect 688 -9 705 9
<< metal1 >>
rect 0 342 720 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 720 342
rect 0 309 720 325
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 370 283 399 289
rect 370 266 376 283
rect 393 282 399 283
rect 610 283 639 289
rect 610 282 616 283
rect 393 268 616 282
rect 393 266 399 268
rect 82 256 111 262
rect 82 239 88 256
rect 105 255 111 256
rect 370 260 399 266
rect 610 266 616 268
rect 633 266 639 283
rect 610 260 639 266
rect 370 255 391 260
rect 105 241 391 255
rect 514 243 543 249
rect 105 239 111 241
rect 82 233 111 239
rect 514 226 520 243
rect 537 241 543 243
rect 537 227 631 241
rect 537 226 543 227
rect 514 220 543 226
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 418 201 447 207
rect 418 184 424 201
rect 441 184 447 201
rect 418 178 447 184
rect 562 201 591 207
rect 562 184 568 201
rect 585 184 591 201
rect 562 178 591 184
rect 137 114 151 178
rect 281 114 295 178
rect 425 114 439 178
rect 569 114 583 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 274 108 303 114
rect 274 91 280 108
rect 297 91 303 108
rect 274 85 303 91
rect 418 108 447 114
rect 418 91 424 108
rect 441 91 447 108
rect 418 85 447 91
rect 562 108 591 114
rect 562 91 568 108
rect 585 91 591 108
rect 562 85 591 91
rect 617 73 631 227
rect 82 67 111 73
rect 82 50 88 67
rect 105 66 111 67
rect 610 67 639 73
rect 610 66 616 67
rect 105 52 616 66
rect 105 50 111 52
rect 82 44 111 50
rect 610 50 616 52
rect 633 50 639 67
rect 610 44 639 50
rect 0 9 720 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 720 9
rect 0 -24 720 -9
<< labels >>
rlabel locali 0 309 720 357 0 VDD
port 1 se
rlabel metal1 0 309 720 357 0 VDD
port 2 se
rlabel locali 0 -24 720 24 0 GND
port 3 se
rlabel metal1 0 -24 720 24 0 GND
port 4 se
rlabel metal1 82 44 111 52 0 Y
port 5 se
rlabel metal1 610 44 639 52 0 Y
port 6 se
rlabel metal1 82 52 639 66 0 Y
port 7 se
rlabel metal1 82 66 111 73 0 Y
port 8 se
rlabel metal1 610 66 639 73 0 Y
port 9 se
rlabel metal1 514 220 543 227 0 Y
port 10 se
rlabel metal1 617 73 631 227 0 Y
port 11 se
rlabel metal1 514 227 631 241 0 Y
port 12 se
rlabel metal1 514 241 543 249 0 Y
port 13 se
rlabel metal1 418 85 447 114 0 C
port 14 se
rlabel metal1 425 114 439 178 0 C
port 15 se
rlabel metal1 418 178 447 207 0 C
port 16 se
rlabel metal1 562 85 591 114 0 D
port 17 se
rlabel metal1 569 114 583 178 0 D
port 18 se
rlabel metal1 562 178 591 207 0 D
port 19 se
rlabel metal1 274 85 303 114 0 A
port 20 se
rlabel metal1 281 114 295 178 0 A
port 21 se
rlabel metal1 274 178 303 207 0 A
port 22 se
rlabel metal1 130 85 159 114 0 B
port 23 se
rlabel metal1 137 114 151 178 0 B
port 24 se
rlabel metal1 130 178 159 207 0 B
port 25 se
<< properties >>
string FIXED_BBOX 0 0 720 333
<< end >>
