VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BUFX4
  CLASS CORE ;
  FOREIGN BUFX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 1.780 2.990 2.070 3.090 ;
        RECT 1.780 2.820 1.840 2.990 ;
        RECT 2.010 2.820 2.070 2.990 ;
        RECT 1.780 2.760 2.070 2.820 ;
        RECT 4.660 2.990 4.950 3.090 ;
        RECT 4.660 2.820 4.720 2.990 ;
        RECT 4.890 2.820 4.950 2.990 ;
        RECT 4.660 2.760 4.950 2.820 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 1.760 2.990 2.090 3.090 ;
        RECT 1.760 2.820 1.840 2.990 ;
        RECT 2.010 2.820 2.090 2.990 ;
        RECT 1.760 2.740 2.090 2.820 ;
        RECT 4.640 2.990 4.970 3.090 ;
        RECT 4.640 2.820 4.720 2.990 ;
        RECT 4.890 2.820 4.970 2.990 ;
        RECT 4.640 2.740 4.970 2.820 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.510 2.070 0.570 ;
        RECT 1.780 0.340 1.840 0.510 ;
        RECT 2.010 0.340 2.070 0.510 ;
        RECT 1.780 0.240 2.070 0.340 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.760 0.510 2.090 0.590 ;
        RECT 1.760 0.340 1.840 0.510 ;
        RECT 2.010 0.340 2.090 0.510 ;
        RECT 1.760 0.240 2.090 0.340 ;
        RECT 4.640 0.510 4.970 0.590 ;
        RECT 4.640 0.340 4.720 0.510 ;
        RECT 4.890 0.340 4.970 0.510 ;
        RECT 4.640 0.240 4.970 0.340 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.700 2.410 3.990 2.490 ;
        RECT 3.700 2.270 4.870 2.410 ;
        RECT 3.700 2.200 3.990 2.270 ;
        RECT 3.700 0.660 3.990 0.730 ;
        RECT 4.730 0.660 4.870 2.270 ;
        RECT 3.700 0.520 4.870 0.660 ;
        RECT 3.700 0.440 3.990 0.520 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.540 1.510 1.780 ;
        RECT 1.300 1.250 1.590 1.540 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 3.680 2.430 4.010 2.510 ;
        RECT 3.680 2.260 3.760 2.430 ;
        RECT 3.930 2.260 4.010 2.430 ;
        RECT 3.680 2.180 4.010 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 4.180 2.010 4.490 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 1.360 1.160 1.530 1.310 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.920 4.240 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.180 0.910 4.240 0.920 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.180 0.830 4.490 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 3.680 0.670 4.010 0.750 ;
        RECT 3.680 0.500 3.760 0.670 ;
        RECT 3.930 0.500 4.010 0.670 ;
        RECT 3.680 0.420 4.010 0.500 ;
      LAYER met1 ;
        RECT 0.580 2.430 0.870 2.490 ;
        RECT 0.580 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.870 2.430 ;
        RECT 0.580 2.200 0.870 2.260 ;
        RECT 0.650 1.060 0.790 2.200 ;
        RECT 2.740 2.010 3.030 2.070 ;
        RECT 2.740 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.030 2.010 ;
        RECT 2.740 1.780 3.030 1.840 ;
        RECT 4.180 2.010 4.470 2.070 ;
        RECT 4.180 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.470 2.010 ;
        RECT 4.180 1.780 4.470 1.840 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 2.740 1.080 3.030 1.140 ;
        RECT 2.740 1.060 2.800 1.080 ;
        RECT 0.650 0.920 2.800 1.060 ;
        RECT 0.650 0.730 0.790 0.920 ;
        RECT 2.740 0.910 2.800 0.920 ;
        RECT 2.970 1.060 3.030 1.080 ;
        RECT 4.180 1.080 4.470 1.140 ;
        RECT 4.180 1.060 4.240 1.080 ;
        RECT 2.970 0.920 4.240 1.060 ;
        RECT 2.970 0.910 3.030 0.920 ;
        RECT 2.740 0.850 3.030 0.910 ;
        RECT 4.180 0.910 4.240 0.920 ;
        RECT 4.410 0.910 4.470 1.080 ;
        RECT 4.180 0.850 4.470 0.910 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.870 0.670 ;
        RECT 0.580 0.440 0.870 0.500 ;
  END
END BUFX4
END LIBRARY

