VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 7.540 2.990 7.830 3.090 ;
        RECT 7.540 2.820 7.600 2.990 ;
        RECT 7.770 2.820 7.830 2.990 ;
        RECT 7.540 2.760 7.830 2.820 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 1.760 2.990 2.090 3.090 ;
        RECT 1.760 2.820 1.840 2.990 ;
        RECT 2.010 2.820 2.090 2.990 ;
        RECT 1.760 2.740 2.090 2.820 ;
        RECT 7.520 2.990 7.850 3.090 ;
        RECT 7.520 2.820 7.600 2.990 ;
        RECT 7.770 2.820 7.850 2.990 ;
        RECT 7.520 2.740 7.850 2.820 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.510 2.070 0.570 ;
        RECT 1.780 0.340 1.840 0.510 ;
        RECT 2.010 0.340 2.070 0.510 ;
        RECT 1.780 0.240 2.070 0.340 ;
        RECT 7.540 0.510 7.830 0.570 ;
        RECT 7.540 0.340 7.600 0.510 ;
        RECT 7.770 0.340 7.830 0.510 ;
        RECT 7.540 0.240 7.830 0.340 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.760 0.510 2.090 0.590 ;
        RECT 1.760 0.340 1.840 0.510 ;
        RECT 2.010 0.340 2.090 0.510 ;
        RECT 1.760 0.240 2.090 0.340 ;
        RECT 7.520 0.510 7.850 0.590 ;
        RECT 7.520 0.340 7.600 0.510 ;
        RECT 7.770 0.340 7.850 0.510 ;
        RECT 7.520 0.240 7.850 0.340 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 0.440 4.950 0.730 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 2.000 1.590 2.070 ;
        RECT 2.740 2.000 3.030 2.070 ;
        RECT 1.300 1.860 3.030 2.000 ;
        RECT 1.300 1.780 1.590 1.860 ;
        RECT 2.740 1.780 3.030 1.860 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
        RECT 2.740 0.850 3.030 1.140 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 2.000 4.470 2.070 ;
        RECT 8.500 2.000 8.790 2.070 ;
        RECT 4.180 1.860 8.790 2.000 ;
        RECT 4.180 1.780 4.470 1.860 ;
        RECT 5.690 1.140 5.830 1.860 ;
        RECT 8.500 1.780 8.790 1.860 ;
        RECT 8.570 1.140 8.710 1.780 ;
        RECT 5.620 0.850 5.910 1.140 ;
        RECT 8.500 0.850 8.790 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 4.640 2.430 4.970 2.510 ;
        RECT 4.640 2.260 4.720 2.430 ;
        RECT 4.890 2.260 4.970 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 4.660 2.180 4.970 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.920 4.490 1.080 ;
        RECT 4.410 0.910 4.470 0.920 ;
        RECT 4.160 0.830 4.470 0.910 ;
        RECT 4.720 0.750 4.890 2.180 ;
        RECT 5.680 2.090 5.850 2.260 ;
        RECT 7.120 2.090 7.290 2.660 ;
        RECT 8.960 2.430 9.290 2.510 ;
        RECT 8.960 2.260 9.040 2.430 ;
        RECT 9.210 2.260 9.290 2.430 ;
        RECT 8.980 2.180 9.290 2.260 ;
        RECT 5.600 2.010 5.930 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 7.040 2.010 7.370 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 8.480 2.010 8.810 2.090 ;
        RECT 8.480 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.810 2.010 ;
        RECT 8.480 1.760 8.810 1.840 ;
        RECT 7.120 1.160 7.290 1.760 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.600 0.830 5.930 0.910 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.370 1.080 ;
        RECT 7.040 0.830 7.370 0.910 ;
        RECT 8.480 1.080 8.810 1.160 ;
        RECT 8.480 0.910 8.560 1.080 ;
        RECT 8.730 0.910 8.810 1.080 ;
        RECT 8.480 0.830 8.810 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 4.640 0.670 4.970 0.750 ;
        RECT 4.640 0.500 4.720 0.670 ;
        RECT 4.890 0.500 4.970 0.670 ;
        RECT 8.980 0.670 9.290 0.750 ;
        RECT 8.980 0.660 9.040 0.670 ;
        RECT 4.640 0.420 4.970 0.500 ;
        RECT 8.960 0.500 9.040 0.660 ;
        RECT 9.210 0.500 9.290 0.670 ;
        RECT 8.960 0.420 9.290 0.500 ;
      LAYER met1 ;
        RECT 7.060 2.830 7.350 2.890 ;
        RECT 7.060 2.820 7.120 2.830 ;
        RECT 0.650 2.680 7.120 2.820 ;
        RECT 0.650 2.490 0.790 2.680 ;
        RECT 7.060 2.660 7.120 2.680 ;
        RECT 7.290 2.660 7.350 2.830 ;
        RECT 7.060 2.600 7.350 2.660 ;
        RECT 0.580 2.430 0.870 2.490 ;
        RECT 0.580 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.870 2.430 ;
        RECT 5.620 2.430 5.910 2.490 ;
        RECT 5.620 2.410 5.680 2.430 ;
        RECT 0.580 2.200 0.870 2.260 ;
        RECT 3.770 2.270 5.680 2.410 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 3.770 1.060 3.910 2.270 ;
        RECT 5.620 2.260 5.680 2.270 ;
        RECT 5.850 2.410 5.910 2.430 ;
        RECT 8.980 2.430 9.270 2.490 ;
        RECT 8.980 2.410 9.040 2.430 ;
        RECT 5.850 2.270 9.040 2.410 ;
        RECT 5.850 2.260 5.910 2.270 ;
        RECT 5.620 2.200 5.910 2.260 ;
        RECT 8.980 2.260 9.040 2.270 ;
        RECT 9.210 2.260 9.270 2.430 ;
        RECT 8.980 2.200 9.270 2.260 ;
        RECT 4.180 1.080 4.470 1.140 ;
        RECT 4.180 1.060 4.240 1.080 ;
        RECT 3.770 0.920 4.240 1.060 ;
        RECT 4.180 0.910 4.240 0.920 ;
        RECT 4.410 0.910 4.470 1.080 ;
        RECT 4.180 0.850 4.470 0.910 ;
        RECT 9.050 0.730 9.190 2.200 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.870 0.670 ;
        RECT 0.580 0.440 0.870 0.500 ;
        RECT 8.980 0.670 9.270 0.730 ;
        RECT 8.980 0.500 9.040 0.670 ;
        RECT 9.210 0.500 9.270 0.670 ;
        RECT 8.980 0.440 9.270 0.500 ;
  END
END XNOR2X1
END LIBRARY

