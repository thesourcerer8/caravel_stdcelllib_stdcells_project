VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.840 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 15.840 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.840 0.240 ;
    END
  END gnd
  PIN YS
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 14.740 2.150 15.030 2.440 ;
        RECT 14.810 0.690 14.950 2.150 ;
        RECT 14.740 0.400 15.030 0.690 ;
    END
  END YS
  PIN YC
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 2.370 2.070 2.440 ;
        RECT 0.890 2.230 2.070 2.370 ;
        RECT 0.890 0.610 1.030 2.230 ;
        RECT 1.780 2.150 2.070 2.230 ;
        RECT 1.780 0.610 2.070 0.690 ;
        RECT 0.890 0.470 2.070 0.610 ;
        RECT 1.780 0.400 2.070 0.470 ;
    END
  END YC
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.750 4.470 2.040 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 4.180 0.800 4.470 1.090 ;
        RECT 4.250 0.610 4.390 0.800 ;
        RECT 8.980 0.610 9.270 0.820 ;
        RECT 4.250 0.530 9.270 0.610 ;
        RECT 4.250 0.470 9.190 0.530 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.750 5.910 2.040 ;
        RECT 11.380 1.750 11.670 2.040 ;
        RECT 5.690 1.150 5.830 1.750 ;
        RECT 11.450 1.150 11.590 1.750 ;
        RECT 5.690 1.090 11.590 1.150 ;
        RECT 5.620 1.010 11.670 1.090 ;
        RECT 5.620 0.800 5.910 1.010 ;
        RECT 11.380 0.800 11.670 1.010 ;
    END
  END A
END HAX1
END LIBRARY

